magic
tech sky130A
timestamp 1614974079
<< error_p >>
rect -107 31 -99 39
rect -97 31 -89 39
rect -115 23 -81 31
rect -107 15 -89 23
rect -115 7 -81 15
rect -107 -1 -99 7
rect -97 -1 -89 7
<< nwell >>
rect -142 45 180 131
<< nmos >>
rect -85 -95 -70 -60
rect -24 -95 -9 -60
rect 35 -95 50 -60
rect 100 -95 115 -60
<< pmos >>
rect -85 68 -70 104
rect -24 68 -9 104
rect 35 68 50 104
rect 100 68 115 104
<< ndiff >>
rect -123 -71 -85 -60
rect -123 -88 -116 -71
rect -99 -88 -85 -71
rect -123 -95 -85 -88
rect -70 -95 -24 -60
rect -9 -95 35 -60
rect 50 -71 100 -60
rect 50 -88 67 -71
rect 84 -88 100 -71
rect 50 -95 100 -88
rect 115 -67 163 -60
rect 115 -85 141 -67
rect 158 -85 163 -67
rect 115 -95 163 -85
<< pdiff >>
rect -120 104 -93 105
rect -120 96 -85 104
rect -120 75 -115 96
rect -98 75 -85 96
rect -120 68 -85 75
rect -70 96 -24 104
rect -70 75 -55 96
rect -37 75 -24 96
rect -70 68 -24 75
rect -9 68 35 104
rect 50 98 100 104
rect 50 77 69 98
rect 86 77 100 98
rect 50 68 100 77
rect 115 95 161 104
rect 115 74 140 95
rect 157 74 161 95
rect 115 68 161 74
rect -120 67 -93 68
<< ndiffc >>
rect -116 -88 -99 -71
rect 67 -88 84 -71
rect 141 -85 158 -67
<< pdiffc >>
rect -115 75 -98 96
rect -55 75 -37 96
rect 69 77 86 98
rect 140 74 157 95
<< poly >>
rect -85 104 -70 122
rect -24 104 -9 120
rect 35 104 50 119
rect 100 104 115 120
rect -85 40 -70 68
rect -115 39 -70 40
rect -116 31 -70 39
rect -24 38 -9 68
rect -116 7 -107 31
rect -89 7 -70 31
rect -116 -2 -70 7
rect -49 1 -9 38
rect -85 -60 -70 -2
rect -24 -60 -9 1
rect 35 44 50 68
rect 35 7 72 44
rect 35 -60 50 7
rect 100 -14 115 68
rect 85 -46 115 -14
rect 100 -60 115 -46
rect -85 -114 -70 -95
rect -24 -112 -9 -95
rect 35 -115 50 -95
rect 100 -115 115 -95
<< polycont >>
rect -107 7 -89 31
<< locali >>
rect -120 148 159 179
rect -160 96 -92 105
rect -60 104 -33 148
rect -160 75 -115 96
rect -98 75 -92 96
rect -160 67 -92 75
rect -63 96 -29 104
rect -63 75 -55 96
rect -37 75 -29 96
rect -63 67 -29 75
rect -160 -17 -134 67
rect -1 -17 27 104
rect 65 98 90 148
rect 65 77 69 98
rect 86 77 90 98
rect 65 69 90 77
rect 135 95 161 104
rect 135 74 140 95
rect 157 74 161 95
rect -160 -42 105 -17
rect -160 -60 -134 -42
rect 135 -60 161 74
rect -160 -71 -91 -60
rect -160 -88 -116 -71
rect -99 -88 -91 -71
rect -160 -97 -91 -88
rect 60 -71 90 -60
rect 60 -88 67 -71
rect 84 -88 90 -71
rect 60 -144 90 -88
rect 135 -67 163 -60
rect 135 -85 141 -67
rect 158 -85 163 -67
rect 135 -95 163 -85
rect -116 -175 169 -144
<< metal1 >>
rect -129 139 168 188
rect -115 39 -79 40
rect -116 -2 -79 39
rect -49 1 -24 38
rect 47 7 72 44
rect -123 -136 -79 -135
rect -123 -179 176 -136
rect -123 -181 -80 -179
<< end >>
