* SPICE3 file created from O21ai.ext - technology: sky130A

.option scale=10000u

.subckt O21ai A2 B1 A1 Y VPWR VGND
X0 VGND A1 a_6_20# SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X1 Y B1 a_6_20# SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X2 VPWR B1 Y w_n13_169# sky130_fd_pr__pfet_01v8 w=51 l=15
X3 a_55_199# A1 VPWR w_n13_169# sky130_fd_pr__pfet_01v8 w=51 l=15
X4 a_6_20# A2 VGND SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X5 Y A2 a_55_199# w_n13_169# sky130_fd_pr__pfet_01v8 w=51 l=15
.ends
