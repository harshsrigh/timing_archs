* SPICE3 file created from vsdcell_nand2_1x.ext - technology: sky130A

.option scale=0.01u

.subckt vsdcell_nand2_1x A B VGND Y VPWR
X0 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 w=97 l=15
X1 a_64_41# A VGND VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X2 VPWR B Y VPWR sky130_fd_pr__pfet_01v8 w=97 l=15
X3 Y B a_64_41# VGND sky130_fd_pr__nfet_01v8 w=42 l=15
C0 Y VPWR 0.13fF
C1 A B 0.03fF
C2 a_64_41# Y 0.06fF
C3 Y A 0.02fF
C4 Y B 0.10fF
C5 VPWR A 0.03fF
C6 VPWR B 0.03fF
C7 Y VGND 0.15fF
C8 VPWR VGND 0.86fF
.ends
