magic
tech sky130A
timestamp 1616071647
<< nwell >>
rect -13 170 202 297
rect -13 169 196 170
<< nmos >>
rect 40 20 55 62
rect 91 20 106 62
rect 139 20 154 62
<< pmos >>
rect 40 199 55 250
rect 91 199 106 250
rect 139 199 154 250
<< ndiff >>
rect 6 55 40 62
rect 6 36 10 55
rect 30 36 40 55
rect 6 20 40 36
rect 55 51 91 62
rect 55 32 64 51
rect 84 32 91 51
rect 55 20 91 32
rect 106 54 139 62
rect 106 35 113 54
rect 133 35 139 54
rect 106 20 139 35
rect 154 53 190 62
rect 154 34 166 53
rect 186 34 190 53
rect 154 20 190 34
<< pdiff >>
rect 6 236 40 250
rect 6 217 11 236
rect 31 217 40 236
rect 6 199 40 217
rect 55 199 91 250
rect 106 232 139 250
rect 106 213 112 232
rect 132 213 139 232
rect 106 199 139 213
rect 154 239 184 250
rect 154 220 160 239
rect 180 220 184 239
rect 154 199 184 220
<< ndiffc >>
rect 10 36 30 55
rect 64 32 84 51
rect 113 35 133 54
rect 166 34 186 53
<< pdiffc >>
rect 11 217 31 236
rect 112 213 132 232
rect 160 220 180 239
<< poly >>
rect 40 250 55 263
rect 91 250 106 264
rect 139 250 154 264
rect 40 152 55 199
rect 91 153 106 199
rect 139 154 154 199
rect 20 144 55 152
rect 20 126 28 144
rect 45 126 55 144
rect 20 118 55 126
rect 76 145 109 153
rect 76 127 82 145
rect 99 127 109 145
rect 76 119 109 127
rect 130 146 160 154
rect 130 128 137 146
rect 154 128 160 146
rect 130 120 160 128
rect 40 62 55 118
rect 91 62 106 119
rect 139 62 154 120
rect 40 7 55 20
rect 91 7 106 20
rect 139 7 154 20
<< polycont >>
rect 28 126 45 144
rect 82 127 99 145
rect 137 128 154 146
<< locali >>
rect 5 290 181 292
rect 5 273 18 290
rect 36 289 181 290
rect 36 273 144 289
rect 5 272 144 273
rect 162 272 181 289
rect 5 268 181 272
rect 11 236 31 268
rect 11 209 31 217
rect 112 232 132 243
rect 112 191 132 213
rect 160 239 180 268
rect 160 209 180 220
rect 112 171 194 191
rect 20 144 53 152
rect 20 126 28 144
rect 45 126 53 144
rect 20 118 53 126
rect 76 145 109 153
rect 76 127 82 145
rect 99 127 109 145
rect 76 119 109 127
rect 130 146 160 154
rect 130 128 137 146
rect 154 128 160 146
rect 130 120 160 128
rect 10 78 133 101
rect 10 55 30 78
rect 10 27 30 36
rect 64 51 84 60
rect 64 10 84 32
rect 113 54 133 78
rect 177 66 194 171
rect 113 27 133 35
rect 158 53 194 66
rect 158 34 166 53
rect 186 34 194 53
rect 158 27 194 34
rect 4 6 186 10
rect 4 4 166 6
rect 4 -13 16 4
rect 33 -11 166 4
rect 183 -11 186 6
rect 33 -13 186 -11
rect 4 -16 186 -13
<< viali >>
rect 18 273 36 290
rect 144 272 162 289
rect 16 -13 33 4
rect 166 -11 183 6
<< metal1 >>
rect 0 290 190 297
rect 0 273 18 290
rect 36 289 190 290
rect 36 273 144 289
rect 0 272 144 273
rect 162 272 190 289
rect 0 260 190 272
rect 0 6 190 15
rect 0 4 166 6
rect 0 -13 16 4
rect 33 -11 166 4
rect 183 -11 190 6
rect 33 -13 190 -11
rect 0 -20 190 -13
<< labels >>
flabel polycont 82 127 99 145 0 FreeSans 120 0 0 0 A2
port 1 nsew signal input
flabel polycont 137 128 154 146 0 FreeSans 120 0 0 0 B1
port 2 nsew signal input
flabel polycont 28 126 45 144 0 FreeSans 120 0 0 0 A1
port 3 nsew signal input
flabel locali 177 53 194 191 0 FreeSans 120 0 0 0 Y
port 4 nsew signal output
flabel metal1 36 260 144 297 0 FreeSans 120 0 0 0 VPWR
port 5 nsew power bidirectional
flabel locali 33 -16 166 10 0 FreeSans 120 0 0 0 VGND
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180 278
<< end >>
