magic
tech sky130A
timestamp 1614951228
<< nwell >>
rect -20 122 387 305
<< nmos >>
rect 49 41 72 83
rect 159 41 182 83
rect 295 43 316 81
<< pmos >>
rect 49 143 72 234
rect 159 143 182 234
rect 295 181 316 224
<< ndiff >>
rect 10 62 49 83
rect 10 45 19 62
rect 36 45 49 62
rect 10 41 49 45
rect 72 41 159 83
rect 182 62 218 83
rect 182 45 192 62
rect 209 45 218 62
rect 182 41 218 45
rect 250 65 295 81
rect 250 48 258 65
rect 275 48 295 65
rect 250 43 295 48
rect 316 70 369 81
rect 316 53 347 70
rect 364 53 369 70
rect 316 43 369 53
<< pdiff >>
rect 7 228 49 234
rect 7 203 18 228
rect 36 203 49 228
rect 7 143 49 203
rect 72 227 159 234
rect 72 202 102 227
rect 120 202 159 227
rect 72 143 159 202
rect 182 228 219 234
rect 182 203 193 228
rect 211 203 219 228
rect 182 196 219 203
rect 250 224 285 225
rect 250 221 295 224
rect 250 198 259 221
rect 277 198 295 221
rect 182 143 218 196
rect 250 181 295 198
rect 316 215 369 224
rect 316 192 346 215
rect 364 192 369 215
rect 316 181 369 192
<< ndiffc >>
rect 19 45 36 62
rect 192 45 209 62
rect 258 48 275 65
rect 347 53 364 70
<< pdiffc >>
rect 18 203 36 228
rect 102 202 120 227
rect 193 203 211 228
rect 259 198 277 221
rect 346 192 364 215
<< psubdiff >>
rect -21 13 129 14
rect -21 -7 85 13
rect 12 -8 85 -7
rect 102 -8 119 13
rect 136 -8 242 13
rect 112 -9 129 -8
<< nsubdiff >>
rect 12 285 130 286
rect 12 261 84 285
rect 102 261 119 285
rect 137 261 203 285
<< psubdiffcont >>
rect 85 -8 102 13
rect 119 -8 136 13
<< nsubdiffcont >>
rect 84 261 102 285
rect 119 261 137 285
<< poly >>
rect 49 234 72 250
rect 159 234 182 250
rect 295 224 316 241
rect 241 151 274 154
rect 295 151 316 181
rect 241 145 316 151
rect 49 125 72 143
rect 15 119 72 125
rect 15 102 25 119
rect 42 102 72 119
rect 15 91 72 102
rect 49 83 72 91
rect 159 124 182 143
rect 241 128 249 145
rect 266 128 316 145
rect 159 119 215 124
rect 241 122 316 128
rect 241 120 274 122
rect 159 102 190 119
rect 207 102 215 119
rect 159 96 215 102
rect 159 83 182 96
rect 295 81 316 122
rect 49 27 72 41
rect 159 26 182 41
rect 295 30 316 43
<< polycont >>
rect 25 102 42 119
rect 249 128 266 145
rect 190 102 207 119
<< locali >>
rect -20 285 372 290
rect -20 281 84 285
rect -20 264 62 281
rect 79 264 84 281
rect -20 261 84 264
rect 102 261 119 285
rect 137 282 372 285
rect 137 265 139 282
rect 156 265 372 282
rect 137 261 372 265
rect -20 258 372 261
rect 18 233 35 258
rect 193 234 210 258
rect 10 228 44 233
rect 10 203 18 228
rect 36 203 44 228
rect 10 197 44 203
rect 94 227 128 233
rect 94 202 102 227
rect 120 202 128 227
rect 94 196 128 202
rect 185 228 219 234
rect 185 203 193 228
rect 211 203 219 228
rect 258 225 278 258
rect 185 197 219 203
rect 250 221 285 225
rect 250 198 259 221
rect 277 198 285 221
rect 106 175 123 196
rect 250 190 285 198
rect 340 215 369 224
rect 340 192 346 215
rect 364 192 369 215
rect 106 169 154 175
rect 106 154 272 169
rect 106 148 274 154
rect 106 143 154 148
rect 241 145 274 148
rect 15 119 50 125
rect 15 102 25 119
rect 42 102 50 119
rect 15 91 50 102
rect 106 76 123 143
rect 241 128 249 145
rect 266 128 274 145
rect 181 119 215 124
rect 241 120 274 128
rect 181 102 190 119
rect 207 102 215 119
rect 181 96 215 102
rect 10 62 45 69
rect 10 45 19 62
rect 36 45 45 62
rect 10 41 45 45
rect 106 62 218 76
rect 106 45 192 62
rect 209 45 218 62
rect 106 41 218 45
rect 250 65 285 71
rect 250 48 258 65
rect 275 48 285 65
rect 250 43 285 48
rect 340 70 369 192
rect 340 53 347 70
rect 364 53 369 70
rect 340 43 369 53
rect 15 21 38 41
rect 256 21 280 43
rect -21 13 383 21
rect -21 8 85 13
rect -21 -9 60 8
rect 77 -8 85 8
rect 102 -8 119 13
rect 136 9 383 13
rect 136 -8 139 9
rect 156 -8 383 9
rect 77 -9 383 -8
rect -21 -14 383 -9
rect -21 -15 242 -14
<< viali >>
rect 62 264 79 281
rect 139 265 156 282
rect 60 -9 77 8
rect 139 -8 156 9
<< metal1 >>
rect -20 282 379 296
rect -20 281 139 282
rect -20 264 62 281
rect 79 265 139 281
rect 156 265 379 282
rect 79 264 379 265
rect -20 248 379 264
rect 241 120 274 154
rect 256 24 383 25
rect -21 9 383 24
rect -21 8 139 9
rect -21 -9 60 8
rect 77 -8 139 8
rect 156 -8 383 9
rect 77 -9 383 -8
rect -21 -18 383 -9
rect 242 -19 383 -18
<< labels >>
flabel locali s 82 -11 138 16 0 FreeSans 120 0 0 0 VGND
port 3 nsew
flabel locali s 82 259 139 287 0 FreeSans 120 0 0 0 VPWR
port 6 nsew
flabel locali 21 96 46 122 0 FreeSans 120 0 0 0 A
port 1 nsew
flabel locali 186 97 211 123 0 FreeSans 120 0 0 0 B
port 2 nsew
flabel locali s 347 112 365 145 0 FreeSans 120 0 0 0 Y
port 8 nsew
rlabel nwell 119 125 182 137 1 erase
rlabel nwell -20 122 387 305 1 erase
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 232 272
string LEFsource USER
string LEForigin 0 0
<< end >>
