.subckt vsdcell_nand4_2x A B C D VGND VPWR Y
X0 Y A NET1 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X1 Y A NET1 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X2 NET3 B NET1 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X3 NET3 B NET1 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X4 NET2 C NET3 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X5 NET2 C NET3 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X6 NET2 D VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X7 NET2 D VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X8 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X9 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X10 Y B VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X11 Y B VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X12 Y C VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X13 Y C VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X14 Y D VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X15 Y D VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
.ends