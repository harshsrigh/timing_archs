* Function: not ((A1 or A2) and B1)
.subckt vsdcell_o21ai A1 A2 B1 VGND VPWR Y
X0 Y B1 NET1 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X1 NET1 A1 VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X2 NET1 A2 VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X3 NET2 A1 VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X4 Y A2 NET2 VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X5 Y B1 VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
.ends