magic
tech sky130A
timestamp 1616166792
<< nwell >>
rect -13 156 154 293
<< nmos >>
rect 37 33 52 75
rect 85 33 100 75
<< pmos >>
rect 37 179 52 239
rect 85 179 100 239
<< ndiff >>
rect 10 61 37 75
rect 10 40 14 61
rect 31 40 37 61
rect 10 33 37 40
rect 52 65 85 75
rect 52 41 60 65
rect 77 41 85 65
rect 52 33 85 41
rect 100 62 135 75
rect 100 38 107 62
rect 124 38 135 62
rect 100 33 135 38
<< pdiff >>
rect 6 228 37 239
rect 6 197 10 228
rect 29 197 37 228
rect 6 179 37 197
rect 52 221 85 239
rect 52 190 60 221
rect 77 190 85 221
rect 52 179 85 190
rect 100 235 136 239
rect 100 197 110 235
rect 130 197 136 235
rect 100 179 136 197
<< ndiffc >>
rect 14 40 31 61
rect 60 41 77 65
rect 107 38 124 62
<< pdiffc >>
rect 10 197 29 228
rect 60 190 77 221
rect 110 197 130 235
<< poly >>
rect 37 239 52 252
rect 85 239 100 254
rect 37 157 52 179
rect 13 148 52 157
rect 13 123 21 148
rect 39 123 52 148
rect 13 115 52 123
rect 37 75 52 115
rect 85 130 100 179
rect 85 122 125 130
rect 85 97 99 122
rect 117 97 125 122
rect 85 88 125 97
rect 85 75 100 88
rect 37 11 52 33
rect 85 13 100 33
<< polycont >>
rect 21 123 39 148
rect 99 97 117 122
<< locali >>
rect 9 261 14 280
rect 31 262 113 280
rect 130 262 140 280
rect 31 261 140 262
rect 9 260 140 261
rect 10 228 29 260
rect 110 235 130 260
rect 10 183 29 197
rect 60 221 77 231
rect 60 159 77 190
rect 110 189 130 197
rect 13 148 77 159
rect 13 123 21 148
rect 39 142 77 148
rect 39 123 43 142
rect 13 115 43 123
rect 94 122 125 130
rect 94 106 99 122
rect 60 97 99 106
rect 117 97 125 122
rect 60 88 125 97
rect 14 61 31 70
rect 14 12 31 40
rect 60 65 77 88
rect 60 33 77 41
rect 107 62 124 70
rect 107 12 124 38
rect 4 8 136 12
rect 4 -11 15 8
rect 32 7 136 8
rect 32 -11 109 7
rect 4 -12 109 -11
rect 126 -12 136 7
rect 4 -16 136 -12
<< viali >>
rect 14 261 31 280
rect 113 262 130 281
rect 15 -11 32 8
rect 109 -12 126 7
<< metal1 >>
rect 0 281 150 290
rect 0 280 113 281
rect 0 261 14 280
rect 31 262 113 280
rect 130 262 150 281
rect 31 261 150 262
rect 0 249 150 261
rect 0 8 141 20
rect 0 -11 15 8
rect 32 7 141 8
rect 32 -11 109 7
rect 0 -12 109 -11
rect 126 -12 141 7
rect 0 -21 141 -12
<< labels >>
flabel polycont 21 123 39 148 0 FreeSans 120 0 0 0 HI
port 0 nsew signal input
flabel polycont 99 97 117 122 0 FreeSans 120 0 0 0 LO
port 1 nsew signal output
flabel locali 4 -16 136 12 0 FreeSans 120 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali 9 260 140 280 0 FreeSans 120 0 0 0 VPWR
port 3 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 200 272
<< end >>
