* SPICE3 file created from nand_3.ext - technology: sky130A

.option scale=10000u

.subckt nand_3 A VPWR VGND B C Y
X0 a_67_30# A VGND SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X1 Y C a_127_30# SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X2 VPWR B Y w_n10_170# sky130_fd_pr__pfet_01v8 w=50 l=15
X3 Y A VPWR w_n10_170# sky130_fd_pr__pfet_01v8 w=50 l=15
X4 a_127_30# B a_67_30# SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X5 Y C VPWR w_n10_170# sky130_fd_pr__pfet_01v8 w=50 l=15
.ends
