magic
tech sky130A
timestamp 1616045808
<< nwell >>
rect -13 146 142 288
<< nmos >>
rect 63 40 78 83
<< pmos >>
rect 63 166 78 236
<< ndiff >>
rect 6 71 63 83
rect 6 53 10 71
rect 27 53 63 71
rect 6 40 63 53
rect 78 70 123 83
rect 78 52 102 70
rect 119 52 123 70
rect 78 40 123 52
<< pdiff >>
rect 6 228 63 236
rect 6 210 10 228
rect 27 210 63 228
rect 6 193 63 210
rect 6 175 10 193
rect 27 175 63 193
rect 6 166 63 175
rect 78 228 123 236
rect 78 210 102 228
rect 119 210 123 228
rect 78 193 123 210
rect 78 175 102 193
rect 119 175 123 193
rect 78 166 123 175
<< ndiffc >>
rect 10 53 27 71
rect 102 52 119 70
<< pdiffc >>
rect 10 210 27 228
rect 10 175 27 193
rect 102 210 119 228
rect 102 175 119 193
<< poly >>
rect 63 236 78 249
rect 63 149 78 166
rect 41 140 78 149
rect 41 122 46 140
rect 63 122 78 140
rect 41 114 78 122
rect 63 83 78 114
rect 63 27 78 40
<< polycont >>
rect 46 122 63 140
<< locali >>
rect 2 282 135 287
rect 2 281 105 282
rect 2 263 17 281
rect 34 264 105 281
rect 122 264 135 282
rect 34 263 135 264
rect 2 257 135 263
rect 6 228 30 257
rect 6 210 10 228
rect 27 210 30 228
rect 6 193 30 210
rect 6 175 10 193
rect 27 175 30 193
rect 6 166 30 175
rect 100 228 120 236
rect 100 210 102 228
rect 119 210 120 228
rect 100 193 120 210
rect 100 175 102 193
rect 119 175 120 193
rect 41 140 65 149
rect 41 122 46 140
rect 63 122 65 140
rect 41 114 65 122
rect 6 71 30 83
rect 6 53 10 71
rect 27 53 30 71
rect 6 18 30 53
rect 100 70 120 175
rect 100 52 102 70
rect 119 52 120 70
rect 100 40 120 52
rect 0 8 135 18
rect 0 -10 14 8
rect 31 -10 104 8
rect 121 -10 135 8
rect 0 -12 135 -10
<< viali >>
rect 17 263 34 281
rect 105 264 122 282
rect 14 -10 31 8
rect 104 -10 121 8
<< metal1 >>
rect -7 282 135 290
rect -7 281 105 282
rect -7 263 17 281
rect 34 264 105 281
rect 122 264 135 282
rect 34 263 135 264
rect -7 250 135 263
rect -8 8 143 24
rect -8 -10 14 8
rect 31 -10 104 8
rect 121 -10 143 8
rect -8 -17 143 -10
<< labels >>
flabel locali s 100 70 120 205 0 FreeSans 120 0 0 0 Y
port 2 nsew signal output
flabel metal1 31 -17 104 24 0 FreeSans 120 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 34 257 105 287 0 FreeSans 120 0 0 0 VPWR
port 4 nsew power bidirectional
flabel locali s 46 122 63 140 0 FreeSans 120 0 0 0 A
port 1 nsew signal input
flabel pwell 31 -17 104 24 0 FreeSans 120 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell 34 257 105 287 0 FreeSans 120 0 0 0 VPB
port 6 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 138 272
<< end >>
