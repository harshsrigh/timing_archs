magic
tech sky130A
timestamp 1616142855
<< nwell >>
rect -13 146 163 288
<< nmos >>
rect 37 40 52 83
rect 102 40 117 83
<< pmos >>
rect 37 166 52 236
rect 102 166 117 236
<< ndiff >>
rect 6 71 37 83
rect 6 53 10 71
rect 27 53 37 71
rect 6 40 37 53
rect 52 40 102 83
rect 117 70 145 83
rect 117 52 124 70
rect 141 52 145 70
rect 117 40 145 52
<< pdiff >>
rect 63 236 88 239
rect 6 228 37 236
rect 6 210 10 228
rect 27 210 37 228
rect 6 193 37 210
rect 6 175 10 193
rect 27 175 37 193
rect 6 166 37 175
rect 52 228 102 236
rect 52 210 67 228
rect 84 210 102 228
rect 52 192 102 210
rect 52 174 67 192
rect 84 174 102 192
rect 52 166 102 174
rect 117 228 145 236
rect 117 210 124 228
rect 141 210 145 228
rect 117 192 145 210
rect 117 174 124 192
rect 141 174 145 192
rect 117 166 145 174
<< ndiffc >>
rect 10 53 27 71
rect 124 52 141 70
<< pdiffc >>
rect 10 210 27 228
rect 10 175 27 193
rect 67 210 84 228
rect 67 174 84 192
rect 124 210 141 228
rect 124 174 141 192
<< psubdiff >>
rect 2 8 149 10
rect 2 -10 14 8
rect 31 -10 70 8
rect 87 -10 120 8
rect 137 -10 149 8
rect 3 -11 142 -10
<< psubdiffcont >>
rect 14 -10 31 8
rect 70 -10 87 8
rect 120 -10 137 8
<< poly >>
rect 37 236 52 249
rect 102 236 117 249
rect 37 140 52 166
rect 15 131 52 140
rect 15 113 20 131
rect 37 113 52 131
rect 15 105 52 113
rect 37 83 52 105
rect 102 137 117 166
rect 102 129 134 137
rect 102 111 109 129
rect 126 111 134 129
rect 102 103 134 111
rect 102 83 117 103
rect 37 27 52 40
rect 102 27 117 40
<< polycont >>
rect 20 113 37 131
rect 109 111 126 129
<< locali >>
rect 2 282 149 287
rect 2 281 70 282
rect 2 263 17 281
rect 34 264 70 281
rect 87 264 121 282
rect 138 264 149 282
rect 34 263 149 264
rect 2 257 149 263
rect 6 228 30 257
rect 6 210 10 228
rect 27 210 30 228
rect 6 193 30 210
rect 6 175 10 193
rect 27 175 30 193
rect 6 166 30 175
rect 63 228 88 239
rect 63 210 67 228
rect 84 210 88 228
rect 63 192 88 210
rect 63 174 67 192
rect 84 174 88 192
rect 63 166 88 174
rect 121 228 145 257
rect 121 210 124 228
rect 141 210 145 228
rect 121 192 145 210
rect 121 174 124 192
rect 141 174 145 192
rect 121 166 145 174
rect 15 131 39 140
rect 63 133 87 166
rect 15 113 20 131
rect 37 113 39 131
rect 15 105 39 113
rect 62 105 87 133
rect 6 71 30 83
rect 6 53 10 71
rect 27 53 30 71
rect 6 18 30 53
rect 64 67 87 105
rect 104 129 134 137
rect 104 111 109 129
rect 126 111 134 129
rect 104 103 134 111
rect 121 70 145 83
rect 121 67 124 70
rect 64 52 124 67
rect 141 52 145 70
rect 64 49 145 52
rect 121 40 145 49
rect 0 8 150 18
rect 0 -10 14 8
rect 31 -10 70 8
rect 87 -10 120 8
rect 137 -10 150 8
rect 0 -12 150 -10
<< viali >>
rect 17 263 34 281
rect 70 264 87 282
rect 121 264 138 282
rect 14 -10 31 8
rect 70 -10 87 8
rect 120 -10 137 8
<< metal1 >>
rect 0 282 151 290
rect 0 281 70 282
rect 0 263 17 281
rect 34 264 70 281
rect 87 264 121 282
rect 138 264 151 282
rect 34 263 151 264
rect 0 250 151 263
rect 0 8 152 24
rect 0 -10 14 8
rect 31 -10 70 8
rect 87 -10 120 8
rect 137 -10 152 8
rect 0 -17 152 -10
<< labels >>
flabel metal1 34 257 105 287 0 FreeSans 120 0 0 0 VPWR
port 4 nsew power bidirectional
flabel nwell 34 257 105 287 0 FreeSans 120 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 31 -17 104 24 0 FreeSans 120 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 109 112 126 130 0 FreeSans 120 0 0 0 B
port 2 nsew signal input
flabel locali s 20 113 37 131 0 FreeSans 120 0 0 0 A
port 1 nsew signal input
flabel locali s 62 105 87 133 0 FreeSans 120 0 0 0 Y
port 7 nsew signal output
flabel locali s 63 169 88 197 0 FreeSans 120 0 0 0 Y
port 7 nsew signal output
flabel locali s 63 205 88 233 0 FreeSans 120 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 151 272
string LEFsymmetry X Y R90
<< end >>
