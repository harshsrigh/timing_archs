* Function: not ((A1 or A2) and (B1 or B2) and C1)
.subckt vsdcell_o221ai A1 A2 B1 B2 C1 VGND VPWR Y
X0 NET4 A1 VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X1 NET4 A2 VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X2 NET1 B1 NET4 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X3 NET1 B2 NET4 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X4 Y C1 NET1 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X5 Y A2 NET2 VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X6 NET2 A1 VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u

X7 NET3 B1 VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X8 Y B2 NET3 VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u

X9 Y C1 VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
.ends