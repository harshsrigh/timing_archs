* SPICE3 file created from sky130_fd_sc_hd__dfxtp_4.ext - technology: sky130A

.option scale=0.005u

.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
X0 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X1 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 w=130 l=30
X2 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 w=130 l=30
X3 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X4 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8 w=200 l=30
X5 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8 w=200 l=30
X6 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X7 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8 w=200 l=30
X8 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 w=130 l=30
X9 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X10 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X11 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8 w=150 l=30
X12 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8 w=200 l=30
X13 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X14 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X15 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X16 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X17 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 w=128 l=30
X18 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X19 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X20 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 w=130 l=30
X21 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X22 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X23 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8 w=128 l=30
X24 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 w=130 l=30
X25 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8 w=128 l=30
X26 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X27 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X28 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8 w=200 l=30
C0 a_1062_300# VGND 0.35fF
C1 D CLK 0.04fF
C2 a_634_183# VGND 0.23fF
C3 a_27_47# D 0.18fF
C4 a_381_47# VPB 0.00fF
C5 a_475_413# a_27_47# 0.37fF
C6 Q VPB 0.00fF
C7 VGND VPWR 0.03fF
C8 a_475_413# a_1062_300# 0.02fF
C9 a_634_183# D 0.03fF
C10 a_193_47# a_381_47# 0.37fF
C11 a_634_183# a_475_413# 0.60fF
C12 D VPWR 0.03fF
C13 a_891_413# VPB 0.00fF
C14 a_475_413# VPWR 0.35fF
C15 a_381_47# CLK 0.01fF
C16 a_27_47# a_381_47# 0.11fF
C17 a_891_413# a_1020_47# 0.03fF
C18 a_975_413# VPWR 0.02fF
C19 a_193_47# a_891_413# 0.27fF
C20 VGND D 0.03fF
C21 a_1062_300# Q 0.99fF
C22 a_475_413# VGND 0.18fF
C23 a_634_183# a_381_47# 0.04fF
C24 VGND a_572_47# 0.01fF
C25 a_891_413# a_27_47# 0.09fF
C26 a_381_47# VPWR 0.12fF
C27 Q VPWR 0.75fF
C28 a_475_413# D 0.03fF
C29 a_193_47# VPB 0.01fF
C30 a_1062_300# a_891_413# 0.59fF
C31 a_634_183# a_891_413# 0.10fF
C32 a_475_413# a_572_47# 0.05fF
C33 VGND a_381_47# 0.09fF
C34 VGND Q 0.51fF
C35 VPB CLK 0.00fF
C36 a_27_47# VPB 0.01fF
C37 a_891_413# VPWR 0.21fF
C38 a_568_413# VPWR 0.01fF
C39 a_1062_300# VPB 0.01fF
C40 a_381_47# D 0.26fF
C41 a_193_47# CLK 0.05fF
C42 a_193_47# a_27_47# 1.31fF
C43 a_634_183# VPB 0.00fF
C44 a_475_413# a_381_47# 0.11fF
C45 a_891_413# VGND 0.18fF
C46 a_193_47# a_1062_300# 0.10fF
C47 VPB VPWR 0.11fF
C48 a_634_183# a_193_47# 0.43fF
C49 a_27_47# CLK 0.41fF
C50 a_475_413# a_891_413# 0.05fF
C51 a_193_47# VPWR 0.33fF
C52 a_1062_300# a_27_47# 0.11fF
C53 a_475_413# a_568_413# 0.04fF
C54 a_634_183# a_27_47# 0.37fF
C55 a_891_413# a_975_413# 0.05fF
C56 VGND a_1020_47# 0.01fF
C57 VPWR CLK 0.06fF
C58 a_634_183# a_1062_300# 0.03fF
C59 a_193_47# VGND 0.50fF
C60 a_27_47# VPWR 0.75fF
C61 D VPB 0.00fF
C62 a_475_413# VPB 0.01fF
C63 a_1062_300# VPWR 0.35fF
C64 a_891_413# Q 0.03fF
C65 a_634_183# VPWR 0.22fF
C66 a_193_47# D 0.22fF
C67 VGND CLK 0.05fF
C68 a_27_47# VGND 0.36fF
C69 a_193_47# a_475_413# 0.39fF
C70 Q VNB 0.07fF
C71 VGND VNB 0.34fF
C72 VPWR VNB 0.35fF
C73 VPB VNB 0.31fF
C74 a_381_47# VNB 0.08fF
C75 a_891_413# VNB 0.37fF
C76 a_1062_300# VNB 0.95fF
C77 a_475_413# VNB 0.36fF
C78 a_634_183# VNB 0.36fF
C79 a_193_47# VNB 0.26fF
C80 a_27_47# VNB 0.35fF
.ends
