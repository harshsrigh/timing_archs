module picorv32a (clk,
    resetn,
    trap,
    mem_valid,
    mem_instr,
    mem_ready,
    mem_addr,
    mem_wdata,
    mem_wstrb,
    mem_rdata,
    mem_la_read,
    mem_la_write,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    pcpi_valid,
    pcpi_insn,
    pcpi_rs1,
    pcpi_rs2,
    pcpi_wr,
    pcpi_rd,
    pcpi_wait,
    pcpi_ready,
    irq,
    eoi,
    trace_valid,
    trace_data);
 input clk;
 input resetn;
 output trap;
 output mem_valid;
 output mem_instr;
 input mem_ready;
 output [31:0] mem_addr;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 input [31:0] mem_rdata;
 output mem_la_read;
 output mem_la_write;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 output pcpi_valid;
 output [31:0] pcpi_insn;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 input pcpi_wr;
 input [31:0] pcpi_rd;
 input pcpi_wait;
 input pcpi_ready;
 input [31:0] irq;
 output [31:0] eoi;
 output trace_valid;
 output [35:0] trace_data;

 sky130_fd_sc_hd__nand2_4 _24349_ (.A(mem_ready),
    .B(mem_valid),
    .Y(_18188_));
 sky130_fd_sc_hd__buf_1 _24350_ (.A(_18188_),
    .X(_18189_));
 sky130_fd_sc_hd__buf_1 _24351_ (.A(_18189_),
    .X(_18190_));
 sky130_fd_sc_hd__buf_1 _24352_ (.A(_18190_),
    .X(_18191_));
 sky130_fd_sc_hd__buf_1 _24353_ (.A(mem_ready),
    .X(_18192_));
 sky130_fd_sc_hd__buf_1 _24354_ (.A(_18192_),
    .X(_18193_));
 sky130_fd_sc_hd__buf_1 _24355_ (.A(mem_valid),
    .X(_18194_));
 sky130_fd_sc_hd__buf_1 _24356_ (.A(_18194_),
    .X(_18195_));
 sky130_fd_sc_hd__nand3_4 _24357_ (.A(mem_rdata[2]),
    .B(_18193_),
    .C(_18195_),
    .Y(_18196_));
 sky130_fd_sc_hd__a21boi_4 _24358_ (.A1(\mem_rdata_q[2] ),
    .A2(_18191_),
    .B1_N(_18196_),
    .Y(_18197_));
 sky130_vsdinv _24359_ (.A(_18197_),
    .Y(\mem_rdata_latched[2] ));
 sky130_fd_sc_hd__buf_1 _24360_ (.A(\mem_rdata_q[26] ),
    .X(_18198_));
 sky130_fd_sc_hd__buf_1 _24361_ (.A(_18191_),
    .X(_18199_));
 sky130_fd_sc_hd__buf_1 _24362_ (.A(_18193_),
    .X(_18200_));
 sky130_fd_sc_hd__buf_1 _24363_ (.A(_18195_),
    .X(_18201_));
 sky130_fd_sc_hd__nand3_4 _24364_ (.A(mem_rdata[26]),
    .B(_18200_),
    .C(_18201_),
    .Y(_18202_));
 sky130_fd_sc_hd__a21boi_4 _24365_ (.A1(_18198_),
    .A2(_18199_),
    .B1_N(_18202_),
    .Y(_18203_));
 sky130_vsdinv _24366_ (.A(_18203_),
    .Y(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__nand3_4 _24367_ (.A(mem_rdata[3]),
    .B(_18192_),
    .C(_18194_),
    .Y(_18204_));
 sky130_fd_sc_hd__a21boi_4 _24368_ (.A1(\mem_rdata_q[3] ),
    .A2(_18190_),
    .B1_N(_18204_),
    .Y(_18205_));
 sky130_vsdinv _24369_ (.A(_18205_),
    .Y(\mem_rdata_latched[3] ));
 sky130_fd_sc_hd__buf_1 _24370_ (.A(_18193_),
    .X(_18206_));
 sky130_fd_sc_hd__buf_1 _24371_ (.A(_18195_),
    .X(_18207_));
 sky130_fd_sc_hd__nand3_4 _24372_ (.A(mem_rdata[27]),
    .B(_18206_),
    .C(_18207_),
    .Y(_18208_));
 sky130_fd_sc_hd__a21boi_4 _24373_ (.A1(\mem_rdata_q[27] ),
    .A2(_18191_),
    .B1_N(_18208_),
    .Y(_18209_));
 sky130_vsdinv _24374_ (.A(_18209_),
    .Y(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__buf_1 _24375_ (.A(_18189_),
    .X(_18210_));
 sky130_fd_sc_hd__buf_1 _24376_ (.A(mem_ready),
    .X(_18211_));
 sky130_fd_sc_hd__buf_1 _24377_ (.A(mem_valid),
    .X(_18212_));
 sky130_fd_sc_hd__nand3_4 _24378_ (.A(mem_rdata[5]),
    .B(_18211_),
    .C(_18212_),
    .Y(_18213_));
 sky130_fd_sc_hd__a21boi_4 _24379_ (.A1(\mem_rdata_q[5] ),
    .A2(_18210_),
    .B1_N(_18213_),
    .Y(_18214_));
 sky130_vsdinv _24380_ (.A(_18214_),
    .Y(_18215_));
 sky130_fd_sc_hd__buf_1 _24381_ (.A(_18215_),
    .X(\mem_rdata_latched[5] ));
 sky130_fd_sc_hd__nand3_4 _24382_ (.A(mem_rdata[4]),
    .B(mem_ready),
    .C(mem_valid),
    .Y(_18216_));
 sky130_fd_sc_hd__a21boi_4 _24383_ (.A1(\mem_rdata_q[4] ),
    .A2(_18189_),
    .B1_N(_18216_),
    .Y(_18217_));
 sky130_vsdinv _24384_ (.A(_18217_),
    .Y(\mem_rdata_latched[4] ));
 sky130_fd_sc_hd__nand3_4 _24385_ (.A(mem_rdata[1]),
    .B(_18211_),
    .C(_18212_),
    .Y(_18218_));
 sky130_fd_sc_hd__a21bo_4 _24386_ (.A1(\mem_rdata_q[1] ),
    .A2(_18210_),
    .B1_N(_18218_),
    .X(\mem_rdata_latched[1] ));
 sky130_fd_sc_hd__nand3_4 _24387_ (.A(mem_rdata[0]),
    .B(_18211_),
    .C(_18212_),
    .Y(_18219_));
 sky130_fd_sc_hd__a21bo_4 _24388_ (.A1(\mem_rdata_q[0] ),
    .A2(_18189_),
    .B1_N(_18219_),
    .X(\mem_rdata_latched[0] ));
 sky130_fd_sc_hd__nand3_4 _24389_ (.A(mem_rdata[6]),
    .B(_18211_),
    .C(_18212_),
    .Y(_18220_));
 sky130_fd_sc_hd__a21boi_4 _24390_ (.A1(\mem_rdata_q[6] ),
    .A2(_18210_),
    .B1_N(_18220_),
    .Y(_18221_));
 sky130_fd_sc_hd__buf_1 _24391_ (.A(_18221_),
    .X(_18222_));
 sky130_vsdinv _24392_ (.A(_18222_),
    .Y(\mem_rdata_latched[6] ));
 sky130_fd_sc_hd__buf_1 _24393_ (.A(resetn),
    .X(_18223_));
 sky130_vsdinv _24394_ (.A(_18223_),
    .Y(_18224_));
 sky130_fd_sc_hd__buf_1 _24395_ (.A(_18224_),
    .X(_18225_));
 sky130_fd_sc_hd__buf_1 _24396_ (.A(_18225_),
    .X(_18226_));
 sky130_fd_sc_hd__buf_1 _24397_ (.A(_18226_),
    .X(_18227_));
 sky130_fd_sc_hd__buf_1 _24398_ (.A(_18227_),
    .X(_18228_));
 sky130_fd_sc_hd__buf_1 _24399_ (.A(_18228_),
    .X(_18229_));
 sky130_fd_sc_hd__buf_1 _24400_ (.A(resetn),
    .X(_18230_));
 sky130_fd_sc_hd__buf_1 _24401_ (.A(_18230_),
    .X(_18231_));
 sky130_fd_sc_hd__buf_1 _24402_ (.A(_18231_),
    .X(_18232_));
 sky130_fd_sc_hd__buf_1 _24403_ (.A(_18232_),
    .X(_18233_));
 sky130_fd_sc_hd__buf_1 _24404_ (.A(_18233_),
    .X(_18234_));
 sky130_fd_sc_hd__buf_1 _24405_ (.A(mem_do_rdata),
    .X(_18235_));
 sky130_vsdinv _24406_ (.A(_18235_),
    .Y(_18236_));
 sky130_fd_sc_hd__buf_1 _24407_ (.A(_18236_),
    .X(_18237_));
 sky130_fd_sc_hd__buf_1 _24408_ (.A(\cpu_state[6] ),
    .X(_18238_));
 sky130_fd_sc_hd__buf_1 _24409_ (.A(_18238_),
    .X(_18239_));
 sky130_fd_sc_hd__buf_1 _24410_ (.A(_18239_),
    .X(_18240_));
 sky130_fd_sc_hd__nand4_4 _24411_ (.A(_18234_),
    .B(_18237_),
    .C(_18240_),
    .D(instr_lw),
    .Y(_18241_));
 sky130_fd_sc_hd__buf_1 _24412_ (.A(\cpu_state[5] ),
    .X(_18242_));
 sky130_fd_sc_hd__buf_1 _24413_ (.A(_18242_),
    .X(_18243_));
 sky130_fd_sc_hd__buf_1 _24414_ (.A(mem_do_wdata),
    .X(_18244_));
 sky130_vsdinv _24415_ (.A(_18244_),
    .Y(_18245_));
 sky130_fd_sc_hd__buf_1 _24416_ (.A(_18245_),
    .X(_18246_));
 sky130_fd_sc_hd__buf_1 _24417_ (.A(_18231_),
    .X(_18247_));
 sky130_fd_sc_hd__buf_1 _24418_ (.A(_18247_),
    .X(_18248_));
 sky130_fd_sc_hd__buf_1 _24419_ (.A(_18248_),
    .X(_18249_));
 sky130_fd_sc_hd__nand4_4 _24420_ (.A(_18243_),
    .B(_18246_),
    .C(_18249_),
    .D(instr_sw),
    .Y(_18250_));
 sky130_fd_sc_hd__nor2_4 _24421_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .Y(_18251_));
 sky130_fd_sc_hd__nor3_4 _24422_ (.A(mem_do_wdata),
    .B(mem_do_rinst),
    .C(mem_do_rdata),
    .Y(_18252_));
 sky130_vsdinv _24423_ (.A(mem_do_rinst),
    .Y(_18253_));
 sky130_fd_sc_hd__nand2_4 _24424_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .Y(_18254_));
 sky130_fd_sc_hd__o32ai_4 _24425_ (.A1(_18188_),
    .A2(_18251_),
    .A3(_18252_),
    .B1(_18253_),
    .B2(_18254_),
    .Y(_18255_));
 sky130_vsdinv _24426_ (.A(mem_do_prefetch),
    .Y(_18256_));
 sky130_fd_sc_hd__a21oi_4 _24427_ (.A1(_18255_),
    .A2(_18230_),
    .B1(_18256_),
    .Y(_18257_));
 sky130_fd_sc_hd__buf_1 _24428_ (.A(_18257_),
    .X(_18258_));
 sky130_fd_sc_hd__buf_1 _24429_ (.A(_18258_),
    .X(_18259_));
 sky130_fd_sc_hd__a21oi_4 _24430_ (.A1(_18241_),
    .A2(_18250_),
    .B1(_18259_),
    .Y(_18260_));
 sky130_fd_sc_hd__nand2_4 _24431_ (.A(resetn),
    .B(\cpu_state[1] ),
    .Y(_18261_));
 sky130_vsdinv _24432_ (.A(_18261_),
    .Y(_18262_));
 sky130_fd_sc_hd__buf_1 _24433_ (.A(_18225_),
    .X(_18263_));
 sky130_fd_sc_hd__buf_1 _24434_ (.A(_18263_),
    .X(_18264_));
 sky130_vsdinv _24435_ (.A(_18242_),
    .Y(_18265_));
 sky130_fd_sc_hd__buf_1 _24436_ (.A(\cpu_state[1] ),
    .X(_18266_));
 sky130_vsdinv _24437_ (.A(_18266_),
    .Y(_18267_));
 sky130_fd_sc_hd__buf_1 _24438_ (.A(_18267_),
    .X(_18268_));
 sky130_vsdinv _24439_ (.A(_18238_),
    .Y(_18269_));
 sky130_fd_sc_hd__buf_1 _24440_ (.A(_18269_),
    .X(_18270_));
 sky130_fd_sc_hd__nand3_4 _24441_ (.A(_18265_),
    .B(_18268_),
    .C(_18270_),
    .Y(_18271_));
 sky130_fd_sc_hd__nor2_4 _24442_ (.A(\cpu_state[5] ),
    .B(\cpu_state[6] ),
    .Y(_18272_));
 sky130_fd_sc_hd__buf_1 _24443_ (.A(_18272_),
    .X(_18273_));
 sky130_fd_sc_hd__buf_1 _24444_ (.A(_18256_),
    .X(_18274_));
 sky130_fd_sc_hd__buf_1 _24445_ (.A(_18255_),
    .X(_18275_));
 sky130_fd_sc_hd__or3_4 _24446_ (.A(_18274_),
    .B(_18226_),
    .C(_18275_),
    .X(_18276_));
 sky130_fd_sc_hd__o22a_4 _24447_ (.A1(_18264_),
    .A2(_18271_),
    .B1(_18273_),
    .B2(_18276_),
    .X(_18277_));
 sky130_fd_sc_hd__o21a_4 _24448_ (.A1(_18256_),
    .A2(_18255_),
    .B1(_18247_),
    .X(_18278_));
 sky130_fd_sc_hd__buf_1 _24449_ (.A(_18278_),
    .X(_18279_));
 sky130_fd_sc_hd__buf_1 _24450_ (.A(_18244_),
    .X(_18280_));
 sky130_fd_sc_hd__a2bb2o_4 _24451_ (.A1_N(_18237_),
    .A2_N(_18269_),
    .B1(_18243_),
    .B2(_18280_),
    .X(_18281_));
 sky130_fd_sc_hd__nand2_4 _24452_ (.A(_18279_),
    .B(_18281_),
    .Y(_18282_));
 sky130_fd_sc_hd__a21boi_4 _24453_ (.A1(_18277_),
    .A2(_18282_),
    .B1_N(\mem_wordsize[0] ),
    .Y(_18283_));
 sky130_fd_sc_hd__a2111o_4 _24454_ (.A1(_18229_),
    .A2(\mem_wordsize[0] ),
    .B1(_18260_),
    .C1(_18262_),
    .D1(_18283_),
    .X(_00666_));
 sky130_fd_sc_hd__buf_1 _24455_ (.A(_18263_),
    .X(_18284_));
 sky130_fd_sc_hd__buf_1 _24456_ (.A(_18284_),
    .X(_18285_));
 sky130_fd_sc_hd__buf_1 _24457_ (.A(_18285_),
    .X(_18286_));
 sky130_vsdinv _24458_ (.A(is_lb_lh_lw_lbu_lhu),
    .Y(_18287_));
 sky130_vsdinv _24459_ (.A(\cpu_state[2] ),
    .Y(_18288_));
 sky130_fd_sc_hd__buf_1 _24460_ (.A(_18288_),
    .X(_18289_));
 sky130_fd_sc_hd__buf_1 _24461_ (.A(_18289_),
    .X(_18290_));
 sky130_fd_sc_hd__buf_1 _24462_ (.A(_18290_),
    .X(_18291_));
 sky130_fd_sc_hd__buf_1 _24463_ (.A(_18291_),
    .X(_18292_));
 sky130_fd_sc_hd__o21a_4 _24464_ (.A1(_18244_),
    .A2(mem_do_rdata),
    .B1(_18223_),
    .X(_18293_));
 sky130_vsdinv _24465_ (.A(_18293_),
    .Y(_18294_));
 sky130_fd_sc_hd__buf_1 _24466_ (.A(\mem_wordsize[2] ),
    .X(_18295_));
 sky130_fd_sc_hd__buf_1 _24467_ (.A(pcpi_rs1[0]),
    .X(_18296_));
 sky130_fd_sc_hd__buf_1 _24468_ (.A(_18296_),
    .X(_18297_));
 sky130_fd_sc_hd__nand2_4 _24469_ (.A(_18295_),
    .B(_18297_),
    .Y(_18298_));
 sky130_vsdinv _24470_ (.A(_18298_),
    .Y(_18299_));
 sky130_fd_sc_hd__buf_1 _24471_ (.A(_18297_),
    .X(_18300_));
 sky130_fd_sc_hd__buf_1 _24472_ (.A(pcpi_rs1[1]),
    .X(_18301_));
 sky130_fd_sc_hd__o21a_4 _24473_ (.A1(_18300_),
    .A2(_18301_),
    .B1(\mem_wordsize[0] ),
    .X(_18302_));
 sky130_fd_sc_hd__nor2_4 _24474_ (.A(_18299_),
    .B(_18302_),
    .Y(_18303_));
 sky130_fd_sc_hd__buf_1 _24475_ (.A(\reg_pc[1] ),
    .X(_18304_));
 sky130_fd_sc_hd__o21a_4 _24476_ (.A1(_18304_),
    .A2(\reg_pc[0] ),
    .B1(mem_do_rinst),
    .X(_18305_));
 sky130_fd_sc_hd__buf_1 _24477_ (.A(_18305_),
    .X(_18306_));
 sky130_fd_sc_hd__and2_4 _24478_ (.A(_18306_),
    .B(_18223_),
    .X(_18307_));
 sky130_vsdinv _24479_ (.A(_18307_),
    .Y(_18308_));
 sky130_fd_sc_hd__o21ai_4 _24480_ (.A1(_18294_),
    .A2(_18303_),
    .B1(_18308_),
    .Y(_18309_));
 sky130_fd_sc_hd__buf_1 _24481_ (.A(_18309_),
    .X(_18310_));
 sky130_fd_sc_hd__buf_1 _24482_ (.A(\irq_mask[2] ),
    .X(_18311_));
 sky130_fd_sc_hd__nor2_4 _24483_ (.A(_18311_),
    .B(irq_active),
    .Y(_18312_));
 sky130_fd_sc_hd__buf_1 _24484_ (.A(_18312_),
    .X(_18313_));
 sky130_vsdinv _24485_ (.A(_18313_),
    .Y(_18314_));
 sky130_fd_sc_hd__buf_1 _24486_ (.A(_18314_),
    .X(_18315_));
 sky130_fd_sc_hd__and2_4 _24487_ (.A(_18310_),
    .B(_18315_),
    .X(_18316_));
 sky130_fd_sc_hd__buf_1 _24488_ (.A(_18316_),
    .X(_18317_));
 sky130_vsdinv _24489_ (.A(instr_rdinstr),
    .Y(_18318_));
 sky130_vsdinv _24490_ (.A(instr_rdinstrh),
    .Y(_18319_));
 sky130_vsdinv _24491_ (.A(instr_rdcycleh),
    .Y(_18320_));
 sky130_vsdinv _24492_ (.A(instr_rdcycle),
    .Y(_18321_));
 sky130_fd_sc_hd__nand4_4 _24493_ (.A(_18318_),
    .B(_18319_),
    .C(_18320_),
    .D(_18321_),
    .Y(_18322_));
 sky130_fd_sc_hd__nor2_4 _24494_ (.A(instr_lbu),
    .B(instr_lb),
    .Y(_18323_));
 sky130_fd_sc_hd__nor2_4 _24495_ (.A(instr_lhu),
    .B(instr_lh),
    .Y(_18324_));
 sky130_fd_sc_hd__nor2_4 _24496_ (.A(instr_slt),
    .B(instr_slti),
    .Y(_18325_));
 sky130_fd_sc_hd__nor2_4 _24497_ (.A(instr_maskirq),
    .B(instr_retirq),
    .Y(_18326_));
 sky130_fd_sc_hd__nand4_4 _24498_ (.A(_18323_),
    .B(_18324_),
    .C(_18325_),
    .D(_18326_),
    .Y(_18327_));
 sky130_fd_sc_hd__nor2_4 _24499_ (.A(instr_setq),
    .B(instr_getq),
    .Y(_18328_));
 sky130_vsdinv _24500_ (.A(instr_bgeu),
    .Y(_18329_));
 sky130_vsdinv _24501_ (.A(instr_bge),
    .Y(_18330_));
 sky130_fd_sc_hd__and3_4 _24502_ (.A(_18328_),
    .B(_18329_),
    .C(_18330_),
    .X(_18331_));
 sky130_fd_sc_hd__nor2_4 _24503_ (.A(instr_sltu),
    .B(instr_sltiu),
    .Y(_18332_));
 sky130_fd_sc_hd__nor2_4 _24504_ (.A(instr_xor),
    .B(instr_xori),
    .Y(_18333_));
 sky130_fd_sc_hd__nand3_4 _24505_ (.A(_18331_),
    .B(_18332_),
    .C(_18333_),
    .Y(_18334_));
 sky130_fd_sc_hd__nor3_4 _24506_ (.A(_18322_),
    .B(_18327_),
    .C(_18334_),
    .Y(_18335_));
 sky130_fd_sc_hd__or3_4 _24507_ (.A(instr_auipc),
    .B(instr_jal),
    .C(instr_lui),
    .X(_18336_));
 sky130_fd_sc_hd__buf_1 _24508_ (.A(_18336_),
    .X(_00368_));
 sky130_fd_sc_hd__nor4_4 _24509_ (.A(instr_srl),
    .B(instr_sra),
    .C(instr_srli),
    .D(instr_srai),
    .Y(_18337_));
 sky130_vsdinv _24510_ (.A(_18337_),
    .Y(_18338_));
 sky130_fd_sc_hd__or4_4 _24511_ (.A(instr_blt),
    .B(instr_bne),
    .C(instr_beq),
    .D(instr_jalr),
    .X(_18339_));
 sky130_fd_sc_hd__nor3_4 _24512_ (.A(_00368_),
    .B(_18338_),
    .C(_18339_),
    .Y(_18340_));
 sky130_fd_sc_hd__nor4_4 _24513_ (.A(instr_or),
    .B(instr_and),
    .C(instr_sll),
    .D(instr_add),
    .Y(_18341_));
 sky130_fd_sc_hd__buf_1 _24514_ (.A(instr_waitirq),
    .X(_18342_));
 sky130_fd_sc_hd__nor4_4 _24515_ (.A(instr_sw),
    .B(instr_lw),
    .C(_18342_),
    .D(instr_timer),
    .Y(_18343_));
 sky130_fd_sc_hd__and2_4 _24516_ (.A(_18341_),
    .B(_18343_),
    .X(_18344_));
 sky130_fd_sc_hd__nor4_4 _24517_ (.A(instr_addi),
    .B(instr_sb),
    .C(instr_sh),
    .D(instr_bltu),
    .Y(_18345_));
 sky130_fd_sc_hd__buf_1 _24518_ (.A(instr_sub),
    .X(_18346_));
 sky130_fd_sc_hd__buf_1 _24519_ (.A(_18346_),
    .X(_18347_));
 sky130_fd_sc_hd__buf_1 _24520_ (.A(_18347_),
    .X(_18348_));
 sky130_fd_sc_hd__buf_1 _24521_ (.A(_18348_),
    .X(_18349_));
 sky130_fd_sc_hd__buf_1 _24522_ (.A(_18349_),
    .X(_18350_));
 sky130_fd_sc_hd__buf_1 _24523_ (.A(_18350_),
    .X(_18351_));
 sky130_fd_sc_hd__buf_1 _24524_ (.A(_18351_),
    .X(_18352_));
 sky130_fd_sc_hd__buf_1 _24525_ (.A(_18352_),
    .X(_18353_));
 sky130_fd_sc_hd__buf_1 _24526_ (.A(_18353_),
    .X(_18354_));
 sky130_fd_sc_hd__nor2_4 _24527_ (.A(_18354_),
    .B(instr_andi),
    .Y(_18355_));
 sky130_fd_sc_hd__nor2_4 _24528_ (.A(instr_slli),
    .B(instr_ori),
    .Y(_18356_));
 sky130_fd_sc_hd__and3_4 _24529_ (.A(_18345_),
    .B(_18355_),
    .C(_18356_),
    .X(_18357_));
 sky130_fd_sc_hd__and4_4 _24530_ (.A(_18335_),
    .B(_18340_),
    .C(_18344_),
    .D(_18357_),
    .X(_18358_));
 sky130_fd_sc_hd__buf_1 _24531_ (.A(_18255_),
    .X(_18359_));
 sky130_fd_sc_hd__buf_1 _24532_ (.A(_18359_),
    .X(_18360_));
 sky130_fd_sc_hd__buf_1 _24533_ (.A(_18274_),
    .X(_18361_));
 sky130_fd_sc_hd__buf_1 _24534_ (.A(_18269_),
    .X(_18362_));
 sky130_fd_sc_hd__a2111o_4 _24535_ (.A1(_18360_),
    .A2(_18233_),
    .B1(_18361_),
    .C1(_18362_),
    .D1(_18310_),
    .X(_18363_));
 sky130_fd_sc_hd__o41a_4 _24536_ (.A1(_18287_),
    .A2(_18292_),
    .A3(_18317_),
    .A4(_18358_),
    .B1(_18363_),
    .X(_18364_));
 sky130_fd_sc_hd__buf_1 _24537_ (.A(_18240_),
    .X(_18365_));
 sky130_fd_sc_hd__and3_4 _24538_ (.A(_18305_),
    .B(_18223_),
    .C(_18312_),
    .X(_18366_));
 sky130_fd_sc_hd__buf_1 _24539_ (.A(_18366_),
    .X(_18367_));
 sky130_vsdinv _24540_ (.A(_18367_),
    .Y(_18368_));
 sky130_fd_sc_hd__buf_1 _24541_ (.A(_18368_),
    .X(_18369_));
 sky130_fd_sc_hd__buf_1 _24542_ (.A(_18293_),
    .X(_18370_));
 sky130_fd_sc_hd__a21oi_4 _24543_ (.A1(_18306_),
    .A2(_18231_),
    .B1(_18370_),
    .Y(_18371_));
 sky130_vsdinv _24544_ (.A(_18371_),
    .Y(_18372_));
 sky130_fd_sc_hd__buf_1 _24545_ (.A(_18372_),
    .X(_18373_));
 sky130_fd_sc_hd__buf_1 _24546_ (.A(_18230_),
    .X(_18374_));
 sky130_fd_sc_hd__buf_1 _24547_ (.A(_18374_),
    .X(_18375_));
 sky130_fd_sc_hd__nand3_4 _24548_ (.A(_18359_),
    .B(_18274_),
    .C(_18375_),
    .Y(_18376_));
 sky130_vsdinv _24549_ (.A(_18376_),
    .Y(_18377_));
 sky130_vsdinv _24550_ (.A(_18278_),
    .Y(_18378_));
 sky130_fd_sc_hd__a211o_4 _24551_ (.A1(_18369_),
    .A2(_18373_),
    .B1(_18377_),
    .C1(_18378_),
    .X(_18379_));
 sky130_vsdinv _24552_ (.A(_18303_),
    .Y(_18380_));
 sky130_vsdinv _24553_ (.A(_18306_),
    .Y(_18381_));
 sky130_fd_sc_hd__nor2_4 _24554_ (.A(_18244_),
    .B(_18235_),
    .Y(_18382_));
 sky130_vsdinv _24555_ (.A(_18382_),
    .Y(_18383_));
 sky130_fd_sc_hd__nand3_4 _24556_ (.A(_18381_),
    .B(_18231_),
    .C(_18383_),
    .Y(_18384_));
 sky130_fd_sc_hd__a21oi_4 _24557_ (.A1(_18380_),
    .A2(_18315_),
    .B1(_18384_),
    .Y(_18385_));
 sky130_fd_sc_hd__nand3_4 _24558_ (.A(_18279_),
    .B(_18376_),
    .C(_18385_),
    .Y(_18386_));
 sky130_fd_sc_hd__buf_1 _24559_ (.A(_18299_),
    .X(_18387_));
 sky130_fd_sc_hd__nand3_4 _24560_ (.A(_18293_),
    .B(_18302_),
    .C(_18313_),
    .Y(_18388_));
 sky130_fd_sc_hd__a211o_4 _24561_ (.A1(_18374_),
    .A2(_18306_),
    .B1(_18387_),
    .C1(_18388_),
    .X(_18389_));
 sky130_fd_sc_hd__and3_4 _24562_ (.A(_18293_),
    .B(_18313_),
    .C(_18299_),
    .X(_18390_));
 sky130_fd_sc_hd__buf_1 _24563_ (.A(_18381_),
    .X(_18391_));
 sky130_fd_sc_hd__buf_1 _24564_ (.A(_18367_),
    .X(_18392_));
 sky130_fd_sc_hd__a21oi_4 _24565_ (.A1(_18390_),
    .A2(_18391_),
    .B1(_18392_),
    .Y(_18393_));
 sky130_fd_sc_hd__or2_4 _24566_ (.A(_18225_),
    .B(_18275_),
    .X(_18394_));
 sky130_fd_sc_hd__buf_1 _24567_ (.A(_18394_),
    .X(_18395_));
 sky130_fd_sc_hd__a211o_4 _24568_ (.A1(_18389_),
    .A2(_18393_),
    .B1(_18361_),
    .C1(_18395_),
    .X(_18396_));
 sky130_fd_sc_hd__nand3_4 _24569_ (.A(_18379_),
    .B(_18386_),
    .C(_18396_),
    .Y(_18397_));
 sky130_fd_sc_hd__a2bb2o_4 _24570_ (.A1_N(_18286_),
    .A2_N(_18364_),
    .B1(_18365_),
    .B2(_18397_),
    .X(_00665_));
 sky130_fd_sc_hd__buf_1 _24571_ (.A(\cpu_state[4] ),
    .X(_18398_));
 sky130_fd_sc_hd__buf_1 _24572_ (.A(_18398_),
    .X(_18399_));
 sky130_fd_sc_hd__buf_1 _24573_ (.A(_18399_),
    .X(_18400_));
 sky130_fd_sc_hd__buf_1 _24574_ (.A(_18359_),
    .X(_18401_));
 sky130_vsdinv _24575_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_18402_));
 sky130_fd_sc_hd__nor2_4 _24576_ (.A(alu_wait),
    .B(_18402_),
    .Y(_18403_));
 sky130_fd_sc_hd__o21a_4 _24577_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .X(_18404_));
 sky130_vsdinv _24578_ (.A(_18404_),
    .Y(_18405_));
 sky130_fd_sc_hd__buf_1 _24579_ (.A(_18405_),
    .X(_18406_));
 sky130_fd_sc_hd__buf_1 _24580_ (.A(_18406_),
    .X(_18407_));
 sky130_fd_sc_hd__buf_1 _24581_ (.A(irq_active),
    .X(_18408_));
 sky130_vsdinv _24582_ (.A(_18408_),
    .Y(_18409_));
 sky130_vsdinv _24583_ (.A(\irq_mask[1] ),
    .Y(_18410_));
 sky130_vsdinv _24584_ (.A(\irq_mask[9] ),
    .Y(_18411_));
 sky130_fd_sc_hd__a22oi_4 _24585_ (.A1(_18410_),
    .A2(\irq_pending[1] ),
    .B1(\irq_pending[9] ),
    .B2(_18411_),
    .Y(_18412_));
 sky130_vsdinv _24586_ (.A(\irq_mask[0] ),
    .Y(_18413_));
 sky130_vsdinv _24587_ (.A(\irq_mask[6] ),
    .Y(_18414_));
 sky130_fd_sc_hd__a22oi_4 _24588_ (.A1(_18413_),
    .A2(\irq_pending[0] ),
    .B1(\irq_pending[6] ),
    .B2(_18414_),
    .Y(_18415_));
 sky130_vsdinv _24589_ (.A(\irq_mask[2] ),
    .Y(_18416_));
 sky130_vsdinv _24590_ (.A(\irq_mask[10] ),
    .Y(_18417_));
 sky130_fd_sc_hd__a22oi_4 _24591_ (.A1(_18416_),
    .A2(\irq_pending[2] ),
    .B1(\irq_pending[10] ),
    .B2(_18417_),
    .Y(_18418_));
 sky130_vsdinv _24592_ (.A(\irq_mask[4] ),
    .Y(_18419_));
 sky130_vsdinv _24593_ (.A(\irq_mask[29] ),
    .Y(_18420_));
 sky130_fd_sc_hd__a22oi_4 _24594_ (.A1(_18419_),
    .A2(\irq_pending[4] ),
    .B1(\irq_pending[29] ),
    .B2(_18420_),
    .Y(_18421_));
 sky130_fd_sc_hd__and4_4 _24595_ (.A(_18412_),
    .B(_18415_),
    .C(_18418_),
    .D(_18421_),
    .X(_18422_));
 sky130_vsdinv _24596_ (.A(\irq_mask[12] ),
    .Y(_18423_));
 sky130_vsdinv _24597_ (.A(\irq_mask[23] ),
    .Y(_18424_));
 sky130_fd_sc_hd__a22oi_4 _24598_ (.A1(_18423_),
    .A2(\irq_pending[12] ),
    .B1(\irq_pending[23] ),
    .B2(_18424_),
    .Y(_18425_));
 sky130_vsdinv _24599_ (.A(\irq_mask[19] ),
    .Y(_18426_));
 sky130_vsdinv _24600_ (.A(\irq_mask[22] ),
    .Y(_18427_));
 sky130_fd_sc_hd__a22oi_4 _24601_ (.A1(_18426_),
    .A2(\irq_pending[19] ),
    .B1(\irq_pending[22] ),
    .B2(_18427_),
    .Y(_18428_));
 sky130_vsdinv _24602_ (.A(\irq_mask[3] ),
    .Y(_18429_));
 sky130_vsdinv _24603_ (.A(\irq_mask[7] ),
    .Y(_18430_));
 sky130_fd_sc_hd__a22oi_4 _24604_ (.A1(_18429_),
    .A2(\irq_pending[3] ),
    .B1(\irq_pending[7] ),
    .B2(_18430_),
    .Y(_18431_));
 sky130_vsdinv _24605_ (.A(\irq_mask[5] ),
    .Y(_18432_));
 sky130_vsdinv _24606_ (.A(\irq_mask[16] ),
    .Y(_18433_));
 sky130_fd_sc_hd__a22oi_4 _24607_ (.A1(_18432_),
    .A2(\irq_pending[5] ),
    .B1(\irq_pending[16] ),
    .B2(_18433_),
    .Y(_18434_));
 sky130_fd_sc_hd__and4_4 _24608_ (.A(_18425_),
    .B(_18428_),
    .C(_18431_),
    .D(_18434_),
    .X(_18435_));
 sky130_vsdinv _24609_ (.A(\irq_mask[8] ),
    .Y(_18436_));
 sky130_vsdinv _24610_ (.A(\irq_mask[14] ),
    .Y(_18437_));
 sky130_fd_sc_hd__a22oi_4 _24611_ (.A1(_18436_),
    .A2(\irq_pending[8] ),
    .B1(\irq_pending[14] ),
    .B2(_18437_),
    .Y(_18438_));
 sky130_vsdinv _24612_ (.A(\irq_mask[11] ),
    .Y(_18439_));
 sky130_vsdinv _24613_ (.A(\irq_mask[20] ),
    .Y(_18440_));
 sky130_fd_sc_hd__a22oi_4 _24614_ (.A1(_18439_),
    .A2(\irq_pending[11] ),
    .B1(\irq_pending[20] ),
    .B2(_18440_),
    .Y(_18441_));
 sky130_vsdinv _24615_ (.A(\irq_mask[15] ),
    .Y(_18442_));
 sky130_vsdinv _24616_ (.A(\irq_mask[21] ),
    .Y(_18443_));
 sky130_fd_sc_hd__a22oi_4 _24617_ (.A1(_18442_),
    .A2(\irq_pending[15] ),
    .B1(\irq_pending[21] ),
    .B2(_18443_),
    .Y(_18444_));
 sky130_vsdinv _24618_ (.A(\irq_mask[13] ),
    .Y(_18445_));
 sky130_vsdinv _24619_ (.A(\irq_mask[28] ),
    .Y(_18446_));
 sky130_fd_sc_hd__a22oi_4 _24620_ (.A1(_18445_),
    .A2(\irq_pending[13] ),
    .B1(\irq_pending[28] ),
    .B2(_18446_),
    .Y(_18447_));
 sky130_fd_sc_hd__and4_4 _24621_ (.A(_18438_),
    .B(_18441_),
    .C(_18444_),
    .D(_18447_),
    .X(_18448_));
 sky130_vsdinv _24622_ (.A(\irq_mask[17] ),
    .Y(_18449_));
 sky130_vsdinv _24623_ (.A(\irq_mask[18] ),
    .Y(_18450_));
 sky130_fd_sc_hd__a22oi_4 _24624_ (.A1(_18449_),
    .A2(\irq_pending[17] ),
    .B1(\irq_pending[18] ),
    .B2(_18450_),
    .Y(_18451_));
 sky130_vsdinv _24625_ (.A(\irq_mask[25] ),
    .Y(_18452_));
 sky130_vsdinv _24626_ (.A(\irq_mask[26] ),
    .Y(_18453_));
 sky130_fd_sc_hd__a22oi_4 _24627_ (.A1(_18452_),
    .A2(\irq_pending[25] ),
    .B1(\irq_pending[26] ),
    .B2(_18453_),
    .Y(_18454_));
 sky130_vsdinv _24628_ (.A(\irq_mask[27] ),
    .Y(_18455_));
 sky130_vsdinv _24629_ (.A(\irq_mask[30] ),
    .Y(_18456_));
 sky130_fd_sc_hd__a22oi_4 _24630_ (.A1(_18455_),
    .A2(\irq_pending[27] ),
    .B1(\irq_pending[30] ),
    .B2(_18456_),
    .Y(_18457_));
 sky130_vsdinv _24631_ (.A(\irq_mask[24] ),
    .Y(_18458_));
 sky130_vsdinv _24632_ (.A(\irq_mask[31] ),
    .Y(_18459_));
 sky130_fd_sc_hd__a22oi_4 _24633_ (.A1(_18458_),
    .A2(\irq_pending[24] ),
    .B1(\irq_pending[31] ),
    .B2(_18459_),
    .Y(_18460_));
 sky130_fd_sc_hd__and4_4 _24634_ (.A(_18451_),
    .B(_18454_),
    .C(_18457_),
    .D(_18460_),
    .X(_18461_));
 sky130_fd_sc_hd__nand4_4 _24635_ (.A(_18422_),
    .B(_18435_),
    .C(_18448_),
    .D(_18461_),
    .Y(_18462_));
 sky130_vsdinv _24636_ (.A(irq_delay),
    .Y(_18463_));
 sky130_fd_sc_hd__nand4_4 _24637_ (.A(_18409_),
    .B(_18462_),
    .C(decoder_trigger),
    .D(_18463_),
    .Y(_18464_));
 sky130_fd_sc_hd__buf_1 _24638_ (.A(_18464_),
    .X(_18465_));
 sky130_fd_sc_hd__buf_1 _24639_ (.A(\irq_state[0] ),
    .X(_18466_));
 sky130_fd_sc_hd__nor2_4 _24640_ (.A(\irq_state[1] ),
    .B(_18466_),
    .Y(_18467_));
 sky130_fd_sc_hd__buf_1 _24641_ (.A(_18467_),
    .X(_18468_));
 sky130_fd_sc_hd__nand3_4 _24642_ (.A(_18465_),
    .B(_18247_),
    .C(_18468_),
    .Y(_18469_));
 sky130_fd_sc_hd__buf_1 _24643_ (.A(_18469_),
    .X(_18470_));
 sky130_fd_sc_hd__nor4_4 _24644_ (.A(_18268_),
    .B(_18369_),
    .C(_18407_),
    .D(_18470_),
    .Y(_18471_));
 sky130_fd_sc_hd__a41o_4 _24645_ (.A1(_18249_),
    .A2(_18400_),
    .A3(_18401_),
    .A4(_18403_),
    .B1(_18471_),
    .X(_18472_));
 sky130_fd_sc_hd__nor3_4 _24646_ (.A(_18311_),
    .B(_18408_),
    .C(_18298_),
    .Y(_18473_));
 sky130_fd_sc_hd__nand3_4 _24647_ (.A(_18381_),
    .B(_18473_),
    .C(_18370_),
    .Y(_18474_));
 sky130_fd_sc_hd__and4_4 _24648_ (.A(_18389_),
    .B(_18310_),
    .C(_18368_),
    .D(_18474_),
    .X(_18475_));
 sky130_vsdinv _24649_ (.A(_18475_),
    .Y(_18476_));
 sky130_fd_sc_hd__buf_1 _24650_ (.A(_18226_),
    .X(_18477_));
 sky130_fd_sc_hd__buf_1 _24651_ (.A(_18477_),
    .X(_18478_));
 sky130_fd_sc_hd__buf_1 _24652_ (.A(_18267_),
    .X(_18479_));
 sky130_fd_sc_hd__buf_1 _24653_ (.A(_18479_),
    .X(_18480_));
 sky130_fd_sc_hd__buf_1 _24654_ (.A(decoder_trigger),
    .X(_18481_));
 sky130_vsdinv _24655_ (.A(_18467_),
    .Y(_18482_));
 sky130_fd_sc_hd__a41oi_4 _24656_ (.A1(_18409_),
    .A2(_18462_),
    .A3(_18481_),
    .A4(_18463_),
    .B1(_18482_),
    .Y(_18483_));
 sky130_fd_sc_hd__buf_1 _24657_ (.A(_18483_),
    .X(_18484_));
 sky130_fd_sc_hd__buf_1 _24658_ (.A(_18484_),
    .X(_18485_));
 sky130_fd_sc_hd__nor4_4 _24659_ (.A(_18478_),
    .B(_18480_),
    .C(_18369_),
    .D(_18485_),
    .Y(_18486_));
 sky130_fd_sc_hd__buf_1 _24660_ (.A(_18302_),
    .X(_18487_));
 sky130_fd_sc_hd__a21o_4 _24661_ (.A1(_18487_),
    .A2(_18314_),
    .B1(_18387_),
    .X(_18488_));
 sky130_fd_sc_hd__o21a_4 _24662_ (.A1(_18384_),
    .A2(_18488_),
    .B1(_18393_),
    .X(_18489_));
 sky130_fd_sc_hd__buf_1 _24663_ (.A(\pcpi_mul.active[1] ),
    .X(_18490_));
 sky130_fd_sc_hd__nor2_4 _24664_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_18491_));
 sky130_fd_sc_hd__nor4_4 _24665_ (.A(_18408_),
    .B(\irq_mask[1] ),
    .C(_18490_),
    .D(_18491_),
    .Y(_18492_));
 sky130_fd_sc_hd__a21boi_4 _24666_ (.A1(_18489_),
    .A2(_18373_),
    .B1_N(_18492_),
    .Y(_18493_));
 sky130_fd_sc_hd__nand3_4 _24667_ (.A(_18389_),
    .B(_18310_),
    .C(_18368_),
    .Y(_18494_));
 sky130_fd_sc_hd__and2_4 _24668_ (.A(_18494_),
    .B(_18490_),
    .X(_18495_));
 sky130_fd_sc_hd__buf_1 _24669_ (.A(_18340_),
    .X(_18496_));
 sky130_fd_sc_hd__and3_4 _24670_ (.A(_18496_),
    .B(_18344_),
    .C(_18357_),
    .X(_18497_));
 sky130_fd_sc_hd__buf_1 _24671_ (.A(\cpu_state[3] ),
    .X(_18498_));
 sky130_fd_sc_hd__buf_1 _24672_ (.A(_18498_),
    .X(_18499_));
 sky130_fd_sc_hd__buf_1 _24673_ (.A(_18499_),
    .X(_18500_));
 sky130_fd_sc_hd__buf_1 _24674_ (.A(_18500_),
    .X(_18501_));
 sky130_fd_sc_hd__buf_1 _24675_ (.A(_18501_),
    .X(_18502_));
 sky130_fd_sc_hd__buf_1 _24676_ (.A(_18335_),
    .X(_18503_));
 sky130_fd_sc_hd__and4_4 _24677_ (.A(_18497_),
    .B(_18248_),
    .C(_18502_),
    .D(_18503_),
    .X(_18504_));
 sky130_fd_sc_hd__o21a_4 _24678_ (.A1(_18493_),
    .A2(_18495_),
    .B1(_18504_),
    .X(_18505_));
 sky130_fd_sc_hd__buf_1 _24679_ (.A(_18375_),
    .X(_18506_));
 sky130_fd_sc_hd__buf_1 _24680_ (.A(_18506_),
    .X(_18507_));
 sky130_fd_sc_hd__nand2_4 _24681_ (.A(_18488_),
    .B(_18383_),
    .Y(_18508_));
 sky130_fd_sc_hd__buf_1 _24682_ (.A(_18374_),
    .X(_18509_));
 sky130_fd_sc_hd__nand3_4 _24683_ (.A(_18508_),
    .B(_18509_),
    .C(_18391_),
    .Y(_18510_));
 sky130_fd_sc_hd__buf_1 _24684_ (.A(_18328_),
    .X(_18511_));
 sky130_vsdinv _24685_ (.A(instr_timer),
    .Y(_18512_));
 sky130_fd_sc_hd__and3_4 _24686_ (.A(_18511_),
    .B(_18326_),
    .C(_18512_),
    .X(_18513_));
 sky130_vsdinv _24687_ (.A(_18513_),
    .Y(_18514_));
 sky130_fd_sc_hd__buf_1 _24688_ (.A(_18514_),
    .X(_18515_));
 sky130_fd_sc_hd__nor2_4 _24689_ (.A(_18322_),
    .B(_18515_),
    .Y(_18516_));
 sky130_fd_sc_hd__a211o_4 _24690_ (.A1(_18510_),
    .A2(_18393_),
    .B1(_18291_),
    .C1(_18516_),
    .X(_18517_));
 sky130_vsdinv _24691_ (.A(_18272_),
    .Y(_18518_));
 sky130_fd_sc_hd__and4_4 _24692_ (.A(_18275_),
    .B(_18274_),
    .C(_18247_),
    .D(_18518_),
    .X(_18519_));
 sky130_fd_sc_hd__buf_1 _24693_ (.A(_18519_),
    .X(_00211_));
 sky130_fd_sc_hd__o21ai_4 _24694_ (.A1(_18392_),
    .A2(_18385_),
    .B1(_00211_),
    .Y(_18520_));
 sky130_fd_sc_hd__buf_1 _24695_ (.A(alu_wait),
    .X(_18521_));
 sky130_vsdinv _24696_ (.A(_18521_),
    .Y(_18522_));
 sky130_fd_sc_hd__nand3_4 _24697_ (.A(_18402_),
    .B(_18522_),
    .C(_18398_),
    .Y(_18523_));
 sky130_fd_sc_hd__o21a_4 _24698_ (.A1(_18387_),
    .A2(_18487_),
    .B1(_18383_),
    .X(_18524_));
 sky130_fd_sc_hd__o21a_4 _24699_ (.A1(_18307_),
    .A2(_18524_),
    .B1(_18315_),
    .X(_18525_));
 sky130_fd_sc_hd__or2_4 _24700_ (.A(_18523_),
    .B(_18525_),
    .X(_18526_));
 sky130_fd_sc_hd__nand4_4 _24701_ (.A(_18507_),
    .B(_18517_),
    .C(_18520_),
    .D(_18526_),
    .Y(_18527_));
 sky130_fd_sc_hd__a2111oi_4 _24702_ (.A1(_18472_),
    .A2(_18476_),
    .B1(_18486_),
    .C1(_18505_),
    .D1(_18527_),
    .Y(_18528_));
 sky130_fd_sc_hd__buf_1 _24703_ (.A(_18477_),
    .X(_18529_));
 sky130_fd_sc_hd__buf_1 _24704_ (.A(_18529_),
    .X(_18530_));
 sky130_fd_sc_hd__buf_1 _24705_ (.A(_18382_),
    .X(_18531_));
 sky130_fd_sc_hd__and2_4 _24706_ (.A(_18357_),
    .B(_18344_),
    .X(_18532_));
 sky130_fd_sc_hd__buf_1 _24707_ (.A(_18500_),
    .X(_18533_));
 sky130_fd_sc_hd__buf_1 _24708_ (.A(_18533_),
    .X(_18534_));
 sky130_fd_sc_hd__and4_4 _24709_ (.A(_18532_),
    .B(_18534_),
    .C(_18503_),
    .D(_18496_),
    .X(_18535_));
 sky130_fd_sc_hd__buf_1 _24710_ (.A(_18509_),
    .X(_18536_));
 sky130_fd_sc_hd__buf_1 _24711_ (.A(_18490_),
    .X(_18537_));
 sky130_fd_sc_hd__and4_4 _24712_ (.A(_18535_),
    .B(_18536_),
    .C(_18537_),
    .D(_18473_),
    .X(_18538_));
 sky130_fd_sc_hd__buf_1 _24713_ (.A(instr_jal),
    .X(_18539_));
 sky130_fd_sc_hd__buf_1 _24714_ (.A(_18539_),
    .X(_18540_));
 sky130_fd_sc_hd__buf_1 _24715_ (.A(_18481_),
    .X(_18541_));
 sky130_fd_sc_hd__buf_1 _24716_ (.A(_18541_),
    .X(_18542_));
 sky130_fd_sc_hd__nand4_4 _24717_ (.A(_18375_),
    .B(_18303_),
    .C(_18540_),
    .D(_18542_),
    .Y(_18543_));
 sky130_fd_sc_hd__buf_1 _24718_ (.A(_18468_),
    .X(_18544_));
 sky130_fd_sc_hd__nand3_4 _24719_ (.A(_18465_),
    .B(_18406_),
    .C(_18544_),
    .Y(_18545_));
 sky130_fd_sc_hd__or2_4 _24720_ (.A(_18543_),
    .B(_18545_),
    .X(_18546_));
 sky130_vsdinv _24721_ (.A(_18483_),
    .Y(_18547_));
 sky130_fd_sc_hd__buf_1 _24722_ (.A(_18232_),
    .X(_18548_));
 sky130_fd_sc_hd__nand3_4 _24723_ (.A(_18547_),
    .B(_18548_),
    .C(_18473_),
    .Y(_18549_));
 sky130_fd_sc_hd__buf_1 _24724_ (.A(_18268_),
    .X(_18550_));
 sky130_fd_sc_hd__buf_1 _24725_ (.A(_18550_),
    .X(_18551_));
 sky130_fd_sc_hd__a21oi_4 _24726_ (.A1(_18546_),
    .A2(_18549_),
    .B1(_18551_),
    .Y(_18552_));
 sky130_fd_sc_hd__buf_1 _24727_ (.A(_18406_),
    .X(_18553_));
 sky130_fd_sc_hd__nor3_4 _24728_ (.A(_18550_),
    .B(_18553_),
    .C(_18470_),
    .Y(_18554_));
 sky130_fd_sc_hd__o32a_4 _24729_ (.A1(_18370_),
    .A2(_00211_),
    .A3(_18554_),
    .B1(_18478_),
    .B2(_18391_),
    .X(_18555_));
 sky130_fd_sc_hd__o41ai_4 _24730_ (.A1(_18530_),
    .A2(_18531_),
    .A3(_18538_),
    .A4(_18552_),
    .B1(_18555_),
    .Y(_18556_));
 sky130_fd_sc_hd__buf_1 _24731_ (.A(_18405_),
    .X(_18557_));
 sky130_fd_sc_hd__or3_4 _24732_ (.A(_18388_),
    .B(_18557_),
    .C(_18469_),
    .X(_18558_));
 sky130_fd_sc_hd__o41ai_4 _24733_ (.A1(_18227_),
    .A2(_18531_),
    .A3(_18487_),
    .A4(_18484_),
    .B1(_18558_),
    .Y(_18559_));
 sky130_fd_sc_hd__nand3_4 _24734_ (.A(_18559_),
    .B(_18308_),
    .C(_18298_),
    .Y(_18560_));
 sky130_fd_sc_hd__nor3_4 _24735_ (.A(_18387_),
    .B(_18388_),
    .C(_18307_),
    .Y(_18561_));
 sky130_vsdinv _24736_ (.A(_18342_),
    .Y(_18562_));
 sky130_fd_sc_hd__nand3_4 _24737_ (.A(_18562_),
    .B(_18539_),
    .C(_18541_),
    .Y(_18563_));
 sky130_vsdinv _24738_ (.A(_18563_),
    .Y(_18564_));
 sky130_fd_sc_hd__o41ai_4 _24739_ (.A1(_18392_),
    .A2(_18371_),
    .A3(_18390_),
    .A4(_18561_),
    .B1(_18564_),
    .Y(_18565_));
 sky130_fd_sc_hd__buf_1 _24740_ (.A(_18481_),
    .X(_18566_));
 sky130_fd_sc_hd__a21oi_4 _24741_ (.A1(_18342_),
    .A2(do_waitirq),
    .B1(_18566_),
    .Y(_18567_));
 sky130_fd_sc_hd__nand4_4 _24742_ (.A(_18313_),
    .B(_18370_),
    .C(_18487_),
    .D(_18298_),
    .Y(_18568_));
 sky130_fd_sc_hd__nand4_4 _24743_ (.A(_18309_),
    .B(_18368_),
    .C(_18474_),
    .D(_18568_),
    .Y(_18569_));
 sky130_vsdinv _24744_ (.A(_18473_),
    .Y(_18570_));
 sky130_fd_sc_hd__a211o_4 _24745_ (.A1(_18380_),
    .A2(_18570_),
    .B1(_18384_),
    .C1(_18405_),
    .X(_18571_));
 sky130_fd_sc_hd__a21boi_4 _24746_ (.A1(_18567_),
    .A2(_18569_),
    .B1_N(_18571_),
    .Y(_18572_));
 sky130_fd_sc_hd__a21oi_4 _24747_ (.A1(_18565_),
    .A2(_18572_),
    .B1(_18470_),
    .Y(_18573_));
 sky130_fd_sc_hd__buf_1 _24748_ (.A(_18263_),
    .X(_18574_));
 sky130_fd_sc_hd__and2_4 _24749_ (.A(_18389_),
    .B(_18372_),
    .X(_18575_));
 sky130_fd_sc_hd__buf_1 _24750_ (.A(_18484_),
    .X(_18576_));
 sky130_fd_sc_hd__nor3_4 _24751_ (.A(_18574_),
    .B(_18575_),
    .C(_18576_),
    .Y(_18577_));
 sky130_fd_sc_hd__nor2_4 _24752_ (.A(_18573_),
    .B(_18577_),
    .Y(_18578_));
 sky130_fd_sc_hd__buf_1 _24753_ (.A(_18480_),
    .X(_18579_));
 sky130_fd_sc_hd__a21o_4 _24754_ (.A1(_18560_),
    .A2(_18578_),
    .B1(_18579_),
    .X(_18580_));
 sky130_fd_sc_hd__nand3_4 _24755_ (.A(_18528_),
    .B(_18556_),
    .C(_18580_),
    .Y(_00660_));
 sky130_fd_sc_hd__buf_1 _24756_ (.A(pcpi_rs1[5]),
    .X(_18581_));
 sky130_fd_sc_hd__buf_1 _24757_ (.A(_18581_),
    .X(_18582_));
 sky130_fd_sc_hd__buf_1 _24758_ (.A(mem_la_wdata[5]),
    .X(_18583_));
 sky130_fd_sc_hd__nor2_4 _24759_ (.A(_18582_),
    .B(_18583_),
    .Y(_18584_));
 sky130_fd_sc_hd__nand2_4 _24760_ (.A(_18582_),
    .B(_18583_),
    .Y(_18585_));
 sky130_vsdinv _24761_ (.A(_18585_),
    .Y(_18586_));
 sky130_fd_sc_hd__buf_1 _24762_ (.A(pcpi_rs1[7]),
    .X(_18587_));
 sky130_fd_sc_hd__buf_1 _24763_ (.A(_18587_),
    .X(_18588_));
 sky130_fd_sc_hd__buf_1 _24764_ (.A(mem_la_wdata[7]),
    .X(_18589_));
 sky130_fd_sc_hd__nand2_4 _24765_ (.A(_18588_),
    .B(_18589_),
    .Y(_18590_));
 sky130_vsdinv _24766_ (.A(_18590_),
    .Y(_18591_));
 sky130_fd_sc_hd__nor2_4 _24767_ (.A(_18588_),
    .B(_18589_),
    .Y(_18592_));
 sky130_fd_sc_hd__o22a_4 _24768_ (.A1(_18584_),
    .A2(_18586_),
    .B1(_18591_),
    .B2(_18592_),
    .X(_18593_));
 sky130_fd_sc_hd__buf_1 _24769_ (.A(pcpi_rs1[6]),
    .X(_18594_));
 sky130_fd_sc_hd__buf_1 _24770_ (.A(mem_la_wdata[6]),
    .X(_18595_));
 sky130_fd_sc_hd__nor2_4 _24771_ (.A(_18594_),
    .B(_18595_),
    .Y(_18596_));
 sky130_fd_sc_hd__nand2_4 _24772_ (.A(_18594_),
    .B(_18595_),
    .Y(_18597_));
 sky130_vsdinv _24773_ (.A(_18597_),
    .Y(_18598_));
 sky130_fd_sc_hd__buf_1 _24774_ (.A(pcpi_rs1[4]),
    .X(_18599_));
 sky130_fd_sc_hd__buf_1 _24775_ (.A(_18599_),
    .X(_18600_));
 sky130_fd_sc_hd__buf_1 _24776_ (.A(mem_la_wdata[4]),
    .X(_18601_));
 sky130_fd_sc_hd__buf_1 _24777_ (.A(_18601_),
    .X(_18602_));
 sky130_fd_sc_hd__nor2_4 _24778_ (.A(_18600_),
    .B(_18602_),
    .Y(_18603_));
 sky130_fd_sc_hd__nand2_4 _24779_ (.A(_18600_),
    .B(_18601_),
    .Y(_18604_));
 sky130_vsdinv _24780_ (.A(_18604_),
    .Y(_18605_));
 sky130_fd_sc_hd__o22a_4 _24781_ (.A1(_18596_),
    .A2(_18598_),
    .B1(_18603_),
    .B2(_18605_),
    .X(_18606_));
 sky130_fd_sc_hd__buf_1 _24782_ (.A(pcpi_rs1[3]),
    .X(_18607_));
 sky130_fd_sc_hd__buf_1 _24783_ (.A(mem_la_wdata[3]),
    .X(_18608_));
 sky130_fd_sc_hd__nor2_4 _24784_ (.A(_18607_),
    .B(_18608_),
    .Y(_18609_));
 sky130_fd_sc_hd__nand2_4 _24785_ (.A(_18607_),
    .B(mem_la_wdata[3]),
    .Y(_18610_));
 sky130_vsdinv _24786_ (.A(_18610_),
    .Y(_18611_));
 sky130_fd_sc_hd__buf_1 _24787_ (.A(pcpi_rs1[2]),
    .X(_18612_));
 sky130_fd_sc_hd__buf_1 _24788_ (.A(_18612_),
    .X(_18613_));
 sky130_fd_sc_hd__buf_1 _24789_ (.A(mem_la_wdata[2]),
    .X(_18614_));
 sky130_fd_sc_hd__nor2_4 _24790_ (.A(_18613_),
    .B(_18614_),
    .Y(_18615_));
 sky130_fd_sc_hd__nand2_4 _24791_ (.A(_18613_),
    .B(_18614_),
    .Y(_18616_));
 sky130_vsdinv _24792_ (.A(_18616_),
    .Y(_18617_));
 sky130_fd_sc_hd__o22a_4 _24793_ (.A1(_18609_),
    .A2(_18611_),
    .B1(_18615_),
    .B2(_18617_),
    .X(_18618_));
 sky130_fd_sc_hd__buf_1 _24794_ (.A(_18301_),
    .X(_18619_));
 sky130_fd_sc_hd__buf_1 _24795_ (.A(_18619_),
    .X(_18620_));
 sky130_fd_sc_hd__buf_1 _24796_ (.A(mem_la_wdata[1]),
    .X(_18621_));
 sky130_fd_sc_hd__buf_1 _24797_ (.A(_18621_),
    .X(_18622_));
 sky130_fd_sc_hd__buf_1 _24798_ (.A(_18622_),
    .X(_18623_));
 sky130_fd_sc_hd__nor2_4 _24799_ (.A(_18620_),
    .B(_18623_),
    .Y(_18624_));
 sky130_fd_sc_hd__nand2_4 _24800_ (.A(_18620_),
    .B(_18622_),
    .Y(_18625_));
 sky130_vsdinv _24801_ (.A(_18625_),
    .Y(_18626_));
 sky130_fd_sc_hd__buf_1 _24802_ (.A(mem_la_wdata[0]),
    .X(_18627_));
 sky130_fd_sc_hd__buf_1 _24803_ (.A(_18627_),
    .X(_18628_));
 sky130_fd_sc_hd__buf_1 _24804_ (.A(_18628_),
    .X(_18629_));
 sky130_fd_sc_hd__buf_1 _24805_ (.A(_18629_),
    .X(_18630_));
 sky130_fd_sc_hd__buf_1 _24806_ (.A(_18630_),
    .X(_18631_));
 sky130_fd_sc_hd__nor2_4 _24807_ (.A(_18300_),
    .B(_18631_),
    .Y(_18632_));
 sky130_fd_sc_hd__nand2_4 _24808_ (.A(pcpi_rs1[0]),
    .B(_18627_),
    .Y(_18633_));
 sky130_vsdinv _24809_ (.A(_18633_),
    .Y(_18634_));
 sky130_fd_sc_hd__o22a_4 _24810_ (.A1(_18624_),
    .A2(_18626_),
    .B1(_18632_),
    .B2(_18634_),
    .X(_18635_));
 sky130_fd_sc_hd__and4_4 _24811_ (.A(_18593_),
    .B(_18606_),
    .C(_18618_),
    .D(_18635_),
    .X(_18636_));
 sky130_fd_sc_hd__buf_1 _24812_ (.A(pcpi_rs1[14]),
    .X(_18637_));
 sky130_fd_sc_hd__buf_1 _24813_ (.A(_18637_),
    .X(_18638_));
 sky130_fd_sc_hd__xnor2_4 _24814_ (.A(_18638_),
    .B(pcpi_rs2[14]),
    .Y(_18639_));
 sky130_fd_sc_hd__buf_1 _24815_ (.A(pcpi_rs1[13]),
    .X(_18640_));
 sky130_fd_sc_hd__xnor2_4 _24816_ (.A(_18640_),
    .B(pcpi_rs2[13]),
    .Y(_18641_));
 sky130_fd_sc_hd__buf_1 _24817_ (.A(pcpi_rs1[15]),
    .X(_18642_));
 sky130_fd_sc_hd__buf_1 _24818_ (.A(pcpi_rs2[15]),
    .X(_18643_));
 sky130_fd_sc_hd__xnor2_4 _24819_ (.A(_18642_),
    .B(_18643_),
    .Y(_18644_));
 sky130_fd_sc_hd__buf_1 _24820_ (.A(pcpi_rs1[12]),
    .X(_18645_));
 sky130_fd_sc_hd__buf_1 _24821_ (.A(_18645_),
    .X(_18646_));
 sky130_fd_sc_hd__buf_1 _24822_ (.A(pcpi_rs2[12]),
    .X(_18647_));
 sky130_fd_sc_hd__xnor2_4 _24823_ (.A(_18646_),
    .B(_18647_),
    .Y(_18648_));
 sky130_fd_sc_hd__and4_4 _24824_ (.A(_18639_),
    .B(_18641_),
    .C(_18644_),
    .D(_18648_),
    .X(_18649_));
 sky130_fd_sc_hd__buf_1 _24825_ (.A(pcpi_rs1[9]),
    .X(_18650_));
 sky130_fd_sc_hd__buf_1 _24826_ (.A(_18650_),
    .X(_18651_));
 sky130_fd_sc_hd__xnor2_4 _24827_ (.A(_18651_),
    .B(pcpi_rs2[9]),
    .Y(_18652_));
 sky130_fd_sc_hd__buf_1 _24828_ (.A(pcpi_rs1[10]),
    .X(_18653_));
 sky130_fd_sc_hd__buf_1 _24829_ (.A(pcpi_rs2[10]),
    .X(_18654_));
 sky130_fd_sc_hd__xnor2_4 _24830_ (.A(_18653_),
    .B(_18654_),
    .Y(_18655_));
 sky130_fd_sc_hd__buf_1 _24831_ (.A(pcpi_rs1[11]),
    .X(_18656_));
 sky130_fd_sc_hd__buf_1 _24832_ (.A(_18656_),
    .X(_18657_));
 sky130_fd_sc_hd__buf_1 _24833_ (.A(pcpi_rs2[11]),
    .X(_18658_));
 sky130_fd_sc_hd__xnor2_4 _24834_ (.A(_18657_),
    .B(_18658_),
    .Y(_18659_));
 sky130_fd_sc_hd__buf_1 _24835_ (.A(pcpi_rs1[8]),
    .X(_18660_));
 sky130_fd_sc_hd__buf_1 _24836_ (.A(pcpi_rs2[8]),
    .X(_18661_));
 sky130_fd_sc_hd__xnor2_4 _24837_ (.A(_18660_),
    .B(_18661_),
    .Y(_18662_));
 sky130_fd_sc_hd__and4_4 _24838_ (.A(_18652_),
    .B(_18655_),
    .C(_18659_),
    .D(_18662_),
    .X(_18663_));
 sky130_fd_sc_hd__nand3_4 _24839_ (.A(_18636_),
    .B(_18649_),
    .C(_18663_),
    .Y(_18664_));
 sky130_fd_sc_hd__buf_1 _24840_ (.A(pcpi_rs1[20]),
    .X(_18665_));
 sky130_fd_sc_hd__buf_1 _24841_ (.A(_18665_),
    .X(_18666_));
 sky130_fd_sc_hd__buf_1 _24842_ (.A(pcpi_rs2[20]),
    .X(_18667_));
 sky130_fd_sc_hd__buf_1 _24843_ (.A(_18667_),
    .X(_18668_));
 sky130_fd_sc_hd__nor2_4 _24844_ (.A(_18666_),
    .B(_18668_),
    .Y(_18669_));
 sky130_fd_sc_hd__nand2_4 _24845_ (.A(_18665_),
    .B(_18667_),
    .Y(_18670_));
 sky130_vsdinv _24846_ (.A(_18670_),
    .Y(_18671_));
 sky130_fd_sc_hd__buf_1 _24847_ (.A(pcpi_rs1[22]),
    .X(_18672_));
 sky130_vsdinv _24848_ (.A(_18672_),
    .Y(_18673_));
 sky130_vsdinv _24849_ (.A(pcpi_rs2[22]),
    .Y(_18674_));
 sky130_fd_sc_hd__nand2_4 _24850_ (.A(_18673_),
    .B(_18674_),
    .Y(_18675_));
 sky130_fd_sc_hd__buf_1 _24851_ (.A(_18672_),
    .X(_18676_));
 sky130_fd_sc_hd__buf_1 _24852_ (.A(pcpi_rs2[22]),
    .X(_18677_));
 sky130_fd_sc_hd__nand2_4 _24853_ (.A(_18676_),
    .B(_18677_),
    .Y(_18678_));
 sky130_fd_sc_hd__a2bb2oi_4 _24854_ (.A1_N(_18669_),
    .A2_N(_18671_),
    .B1(_18675_),
    .B2(_18678_),
    .Y(_18679_));
 sky130_fd_sc_hd__buf_1 _24855_ (.A(pcpi_rs1[21]),
    .X(_18680_));
 sky130_fd_sc_hd__buf_1 _24856_ (.A(pcpi_rs2[21]),
    .X(_18681_));
 sky130_fd_sc_hd__buf_1 _24857_ (.A(_18681_),
    .X(_18682_));
 sky130_fd_sc_hd__nor2_4 _24858_ (.A(_18680_),
    .B(_18682_),
    .Y(_18683_));
 sky130_fd_sc_hd__nand2_4 _24859_ (.A(pcpi_rs1[21]),
    .B(_18681_),
    .Y(_18684_));
 sky130_vsdinv _24860_ (.A(_18684_),
    .Y(_18685_));
 sky130_fd_sc_hd__nand2_4 _24861_ (.A(pcpi_rs1[23]),
    .B(pcpi_rs2[23]),
    .Y(_18686_));
 sky130_vsdinv _24862_ (.A(_18686_),
    .Y(_18687_));
 sky130_fd_sc_hd__buf_1 _24863_ (.A(pcpi_rs1[23]),
    .X(_18688_));
 sky130_fd_sc_hd__buf_1 _24864_ (.A(pcpi_rs2[23]),
    .X(_18689_));
 sky130_fd_sc_hd__nor2_4 _24865_ (.A(_18688_),
    .B(_18689_),
    .Y(_18690_));
 sky130_fd_sc_hd__o22a_4 _24866_ (.A1(_18683_),
    .A2(_18685_),
    .B1(_18687_),
    .B2(_18690_),
    .X(_18691_));
 sky130_fd_sc_hd__and2_4 _24867_ (.A(_18679_),
    .B(_18691_),
    .X(_18692_));
 sky130_fd_sc_hd__buf_1 _24868_ (.A(pcpi_rs1[19]),
    .X(_18693_));
 sky130_fd_sc_hd__buf_1 _24869_ (.A(_18693_),
    .X(_18694_));
 sky130_fd_sc_hd__buf_1 _24870_ (.A(pcpi_rs2[19]),
    .X(_18695_));
 sky130_fd_sc_hd__buf_1 _24871_ (.A(_18695_),
    .X(_18696_));
 sky130_fd_sc_hd__nor2_4 _24872_ (.A(_18694_),
    .B(_18696_),
    .Y(_18697_));
 sky130_fd_sc_hd__nand2_4 _24873_ (.A(_18693_),
    .B(_18695_),
    .Y(_18698_));
 sky130_vsdinv _24874_ (.A(_18698_),
    .Y(_18699_));
 sky130_fd_sc_hd__buf_1 _24875_ (.A(pcpi_rs1[18]),
    .X(_18700_));
 sky130_vsdinv _24876_ (.A(_18700_),
    .Y(_18701_));
 sky130_vsdinv _24877_ (.A(pcpi_rs2[18]),
    .Y(_18702_));
 sky130_fd_sc_hd__buf_1 _24878_ (.A(_18702_),
    .X(_18703_));
 sky130_fd_sc_hd__nand2_4 _24879_ (.A(_18701_),
    .B(_18703_),
    .Y(_18704_));
 sky130_fd_sc_hd__buf_1 _24880_ (.A(_18700_),
    .X(_18705_));
 sky130_fd_sc_hd__buf_1 _24881_ (.A(pcpi_rs2[18]),
    .X(_18706_));
 sky130_fd_sc_hd__nand2_4 _24882_ (.A(_18705_),
    .B(_18706_),
    .Y(_18707_));
 sky130_fd_sc_hd__a2bb2oi_4 _24883_ (.A1_N(_18697_),
    .A2_N(_18699_),
    .B1(_18704_),
    .B2(_18707_),
    .Y(_18708_));
 sky130_fd_sc_hd__buf_1 _24884_ (.A(pcpi_rs1[16]),
    .X(_18709_));
 sky130_fd_sc_hd__buf_1 _24885_ (.A(_18709_),
    .X(_18710_));
 sky130_fd_sc_hd__buf_1 _24886_ (.A(pcpi_rs2[16]),
    .X(_18711_));
 sky130_fd_sc_hd__buf_1 _24887_ (.A(_18711_),
    .X(_18712_));
 sky130_fd_sc_hd__xnor2_4 _24888_ (.A(_18710_),
    .B(_18712_),
    .Y(_18713_));
 sky130_fd_sc_hd__buf_1 _24889_ (.A(pcpi_rs1[17]),
    .X(_18714_));
 sky130_fd_sc_hd__buf_1 _24890_ (.A(_18714_),
    .X(_18715_));
 sky130_fd_sc_hd__buf_1 _24891_ (.A(pcpi_rs2[17]),
    .X(_18716_));
 sky130_fd_sc_hd__buf_1 _24892_ (.A(_18716_),
    .X(_18717_));
 sky130_fd_sc_hd__xnor2_4 _24893_ (.A(_18715_),
    .B(_18717_),
    .Y(_18718_));
 sky130_fd_sc_hd__and4_4 _24894_ (.A(_18692_),
    .B(_18708_),
    .C(_18713_),
    .D(_18718_),
    .X(_18719_));
 sky130_fd_sc_hd__buf_1 _24895_ (.A(pcpi_rs1[26]),
    .X(_18720_));
 sky130_fd_sc_hd__buf_1 _24896_ (.A(_18720_),
    .X(_18721_));
 sky130_fd_sc_hd__buf_1 _24897_ (.A(pcpi_rs2[26]),
    .X(_18722_));
 sky130_fd_sc_hd__nor2_4 _24898_ (.A(_18721_),
    .B(_18722_),
    .Y(_18723_));
 sky130_fd_sc_hd__buf_1 _24899_ (.A(_18720_),
    .X(_18724_));
 sky130_fd_sc_hd__nand2_4 _24900_ (.A(_18724_),
    .B(_18722_),
    .Y(_18725_));
 sky130_vsdinv _24901_ (.A(_18725_),
    .Y(_18726_));
 sky130_vsdinv _24902_ (.A(pcpi_rs1[24]),
    .Y(_18727_));
 sky130_fd_sc_hd__buf_1 _24903_ (.A(_18727_),
    .X(_18728_));
 sky130_vsdinv _24904_ (.A(pcpi_rs2[24]),
    .Y(_18729_));
 sky130_fd_sc_hd__nand2_4 _24905_ (.A(_18728_),
    .B(_18729_),
    .Y(_18730_));
 sky130_fd_sc_hd__buf_1 _24906_ (.A(pcpi_rs1[24]),
    .X(_18731_));
 sky130_fd_sc_hd__buf_1 _24907_ (.A(_18731_),
    .X(_18732_));
 sky130_fd_sc_hd__buf_1 _24908_ (.A(pcpi_rs2[24]),
    .X(_18733_));
 sky130_fd_sc_hd__buf_1 _24909_ (.A(_18733_),
    .X(_18734_));
 sky130_fd_sc_hd__nand2_4 _24910_ (.A(_18732_),
    .B(_18734_),
    .Y(_18735_));
 sky130_fd_sc_hd__a2bb2oi_4 _24911_ (.A1_N(_18723_),
    .A2_N(_18726_),
    .B1(_18730_),
    .B2(_18735_),
    .Y(_18736_));
 sky130_fd_sc_hd__buf_1 _24912_ (.A(pcpi_rs2[30]),
    .X(_18737_));
 sky130_fd_sc_hd__nor2_4 _24913_ (.A(pcpi_rs1[30]),
    .B(_18737_),
    .Y(_18738_));
 sky130_fd_sc_hd__nand2_4 _24914_ (.A(pcpi_rs1[30]),
    .B(pcpi_rs2[30]),
    .Y(_18739_));
 sky130_vsdinv _24915_ (.A(_18739_),
    .Y(_18740_));
 sky130_fd_sc_hd__buf_1 _24916_ (.A(pcpi_rs1[31]),
    .X(_18741_));
 sky130_fd_sc_hd__nand2_4 _24917_ (.A(_18741_),
    .B(pcpi_rs2[31]),
    .Y(_18742_));
 sky130_vsdinv _24918_ (.A(_18742_),
    .Y(_18743_));
 sky130_fd_sc_hd__nor2_4 _24919_ (.A(_18741_),
    .B(pcpi_rs2[31]),
    .Y(_18744_));
 sky130_fd_sc_hd__o22a_4 _24920_ (.A1(_18738_),
    .A2(_18740_),
    .B1(_18743_),
    .B2(_18744_),
    .X(_18745_));
 sky130_fd_sc_hd__buf_1 _24921_ (.A(pcpi_rs1[28]),
    .X(_18746_));
 sky130_fd_sc_hd__buf_1 _24922_ (.A(pcpi_rs2[28]),
    .X(_18747_));
 sky130_fd_sc_hd__nor2_4 _24923_ (.A(_18746_),
    .B(_18747_),
    .Y(_18748_));
 sky130_fd_sc_hd__nand2_4 _24924_ (.A(_18746_),
    .B(pcpi_rs2[28]),
    .Y(_18749_));
 sky130_vsdinv _24925_ (.A(_18749_),
    .Y(_18750_));
 sky130_fd_sc_hd__buf_1 _24926_ (.A(pcpi_rs1[29]),
    .X(_18751_));
 sky130_fd_sc_hd__buf_1 _24927_ (.A(pcpi_rs2[29]),
    .X(_18752_));
 sky130_fd_sc_hd__nand2_4 _24928_ (.A(_18751_),
    .B(_18752_),
    .Y(_18753_));
 sky130_vsdinv _24929_ (.A(_18753_),
    .Y(_18754_));
 sky130_fd_sc_hd__nor2_4 _24930_ (.A(_18751_),
    .B(_18752_),
    .Y(_18755_));
 sky130_fd_sc_hd__o22a_4 _24931_ (.A1(_18748_),
    .A2(_18750_),
    .B1(_18754_),
    .B2(_18755_),
    .X(_18756_));
 sky130_fd_sc_hd__buf_1 _24932_ (.A(pcpi_rs1[27]),
    .X(_18757_));
 sky130_vsdinv _24933_ (.A(_18757_),
    .Y(_18758_));
 sky130_vsdinv _24934_ (.A(pcpi_rs2[27]),
    .Y(_18759_));
 sky130_fd_sc_hd__buf_1 _24935_ (.A(_18759_),
    .X(_18760_));
 sky130_fd_sc_hd__nand2_4 _24936_ (.A(_18758_),
    .B(_18760_),
    .Y(_18761_));
 sky130_fd_sc_hd__buf_1 _24937_ (.A(pcpi_rs2[27]),
    .X(_18762_));
 sky130_fd_sc_hd__nand2_4 _24938_ (.A(_18757_),
    .B(_18762_),
    .Y(_18763_));
 sky130_fd_sc_hd__buf_1 _24939_ (.A(pcpi_rs1[25]),
    .X(_18764_));
 sky130_fd_sc_hd__buf_1 _24940_ (.A(_18764_),
    .X(_18765_));
 sky130_fd_sc_hd__buf_1 _24941_ (.A(_18765_),
    .X(_18766_));
 sky130_fd_sc_hd__buf_1 _24942_ (.A(pcpi_rs2[25]),
    .X(_18767_));
 sky130_fd_sc_hd__nor2_4 _24943_ (.A(_18766_),
    .B(_18767_),
    .Y(_18768_));
 sky130_vsdinv _24944_ (.A(_18768_),
    .Y(_18769_));
 sky130_fd_sc_hd__nand2_4 _24945_ (.A(_18766_),
    .B(_18767_),
    .Y(_18770_));
 sky130_fd_sc_hd__a22oi_4 _24946_ (.A1(_18761_),
    .A2(_18763_),
    .B1(_18769_),
    .B2(_18770_),
    .Y(_18771_));
 sky130_fd_sc_hd__and4_4 _24947_ (.A(_18736_),
    .B(_18745_),
    .C(_18756_),
    .D(_18771_),
    .X(_18772_));
 sky130_fd_sc_hd__nand2_4 _24948_ (.A(_18719_),
    .B(_18772_),
    .Y(_18773_));
 sky130_fd_sc_hd__nor2_4 _24949_ (.A(_18664_),
    .B(_18773_),
    .Y(_00000_));
 sky130_fd_sc_hd__buf_1 _24950_ (.A(_18539_),
    .X(_18774_));
 sky130_fd_sc_hd__buf_1 _24951_ (.A(_18774_),
    .X(_18775_));
 sky130_fd_sc_hd__buf_1 _24952_ (.A(_18775_),
    .X(_18776_));
 sky130_fd_sc_hd__buf_1 _24953_ (.A(_18776_),
    .X(_18777_));
 sky130_fd_sc_hd__buf_1 _24954_ (.A(_18465_),
    .X(_18778_));
 sky130_fd_sc_hd__and4_4 _24955_ (.A(_18778_),
    .B(_18566_),
    .C(_18406_),
    .D(_18544_),
    .X(_18779_));
 sky130_fd_sc_hd__buf_1 _24956_ (.A(_18779_),
    .X(_18780_));
 sky130_fd_sc_hd__buf_1 _24957_ (.A(_18780_),
    .X(_18781_));
 sky130_vsdinv _24958_ (.A(_18781_),
    .Y(_18782_));
 sky130_fd_sc_hd__nor4_4 _24959_ (.A(_18777_),
    .B(_18261_),
    .C(_18525_),
    .D(_18782_),
    .Y(_00661_));
 sky130_fd_sc_hd__buf_1 _24960_ (.A(_18529_),
    .X(_18783_));
 sky130_fd_sc_hd__buf_1 _24961_ (.A(_18783_),
    .X(_18784_));
 sky130_fd_sc_hd__nor2_4 _24962_ (.A(\cpu_state[0] ),
    .B(_18525_),
    .Y(_18785_));
 sky130_fd_sc_hd__buf_1 _24963_ (.A(_18226_),
    .X(_18786_));
 sky130_vsdinv _24964_ (.A(_18533_),
    .Y(_18787_));
 sky130_fd_sc_hd__buf_1 _24965_ (.A(_18787_),
    .X(_18788_));
 sky130_vsdinv _24966_ (.A(_18358_),
    .Y(_18789_));
 sky130_fd_sc_hd__or4_4 _24967_ (.A(_18786_),
    .B(_18537_),
    .C(_18788_),
    .D(_18789_),
    .X(_18790_));
 sky130_fd_sc_hd__a2111o_4 _24968_ (.A1(_18409_),
    .A2(_18410_),
    .B1(_18475_),
    .C1(_18491_),
    .D1(_18790_),
    .X(_18791_));
 sky130_fd_sc_hd__o21ai_4 _24969_ (.A1(_18784_),
    .A2(_18785_),
    .B1(_18791_),
    .Y(_00659_));
 sky130_vsdinv _24970_ (.A(_18491_),
    .Y(_18792_));
 sky130_vsdinv _24971_ (.A(_18504_),
    .Y(_18793_));
 sky130_fd_sc_hd__buf_1 _24972_ (.A(is_lui_auipc_jal),
    .X(_18794_));
 sky130_fd_sc_hd__buf_1 _24973_ (.A(_18794_),
    .X(_18795_));
 sky130_fd_sc_hd__nor3_4 _24974_ (.A(_18795_),
    .B(is_slli_srli_srai),
    .C(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .Y(_18796_));
 sky130_fd_sc_hd__buf_1 _24975_ (.A(\cpu_state[2] ),
    .X(_18797_));
 sky130_fd_sc_hd__buf_1 _24976_ (.A(_18797_),
    .X(_18798_));
 sky130_fd_sc_hd__nand3_4 _24977_ (.A(_18796_),
    .B(_18248_),
    .C(_18798_),
    .Y(_18799_));
 sky130_fd_sc_hd__buf_1 _24978_ (.A(_18514_),
    .X(_18800_));
 sky130_fd_sc_hd__or3_4 _24979_ (.A(_18322_),
    .B(_18799_),
    .C(_18800_),
    .X(_18801_));
 sky130_fd_sc_hd__a41oi_4 _24980_ (.A1(_18335_),
    .A2(_18496_),
    .A3(_18344_),
    .A4(_18357_),
    .B1(_18287_),
    .Y(_18802_));
 sky130_fd_sc_hd__a211o_4 _24981_ (.A1(_18373_),
    .A2(_18489_),
    .B1(_18801_),
    .C1(_18802_),
    .X(_18803_));
 sky130_fd_sc_hd__o41ai_4 _24982_ (.A1(_18537_),
    .A2(_18317_),
    .A3(_18792_),
    .A4(_18793_),
    .B1(_18803_),
    .Y(_00662_));
 sky130_fd_sc_hd__o32a_4 _24983_ (.A1(_18317_),
    .A2(_18377_),
    .A3(_18378_),
    .B1(_18276_),
    .B2(_18475_),
    .X(_18804_));
 sky130_fd_sc_hd__buf_1 _24984_ (.A(_18574_),
    .X(_18805_));
 sky130_fd_sc_hd__buf_1 _24985_ (.A(_18788_),
    .X(_18806_));
 sky130_vsdinv _24986_ (.A(is_sb_sh_sw),
    .Y(_18807_));
 sky130_fd_sc_hd__buf_1 _24987_ (.A(_18807_),
    .X(_18808_));
 sky130_fd_sc_hd__a2111o_4 _24988_ (.A1(_18489_),
    .A2(_18373_),
    .B1(_18805_),
    .C1(_18806_),
    .D1(_18808_),
    .X(_18809_));
 sky130_fd_sc_hd__o21ai_4 _24989_ (.A1(_18265_),
    .A2(_18804_),
    .B1(_18809_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand2_4 _24990_ (.A(_18230_),
    .B(pcpi_valid),
    .Y(_18810_));
 sky130_vsdinv _24991_ (.A(pcpi_insn[3]),
    .Y(_18811_));
 sky130_vsdinv _24992_ (.A(pcpi_insn[2]),
    .Y(_18812_));
 sky130_fd_sc_hd__nand4_4 _24993_ (.A(pcpi_insn[1]),
    .B(_18811_),
    .C(_18812_),
    .D(pcpi_insn[0]),
    .Y(_18813_));
 sky130_vsdinv _24994_ (.A(pcpi_insn[29]),
    .Y(_18814_));
 sky130_vsdinv _24995_ (.A(pcpi_insn[6]),
    .Y(_18815_));
 sky130_vsdinv _24996_ (.A(pcpi_insn[26]),
    .Y(_18816_));
 sky130_fd_sc_hd__nand4_4 _24997_ (.A(pcpi_insn[5]),
    .B(_18815_),
    .C(_18816_),
    .D(pcpi_insn[4]),
    .Y(_18817_));
 sky130_vsdinv _24998_ (.A(pcpi_insn[28]),
    .Y(_18818_));
 sky130_vsdinv _24999_ (.A(pcpi_insn[27]),
    .Y(_18819_));
 sky130_vsdinv _25000_ (.A(pcpi_insn[30]),
    .Y(_18820_));
 sky130_fd_sc_hd__nand4_4 _25001_ (.A(pcpi_insn[25]),
    .B(_18818_),
    .C(_18819_),
    .D(_18820_),
    .Y(_18821_));
 sky130_fd_sc_hd__nor2_4 _25002_ (.A(_18817_),
    .B(_18821_),
    .Y(_18822_));
 sky130_vsdinv _25003_ (.A(pcpi_insn[31]),
    .Y(_18823_));
 sky130_vsdinv _25004_ (.A(pcpi_insn[14]),
    .Y(_18824_));
 sky130_fd_sc_hd__nand4_4 _25005_ (.A(_18814_),
    .B(_18822_),
    .C(_18823_),
    .D(_18824_),
    .Y(_18825_));
 sky130_fd_sc_hd__nor3_4 _25006_ (.A(_18810_),
    .B(_18813_),
    .C(_18825_),
    .Y(_18826_));
 sky130_fd_sc_hd__o21a_4 _25007_ (.A1(pcpi_insn[13]),
    .A2(pcpi_insn[12]),
    .B1(_18826_),
    .X(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__or3_4 _25008_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_00371_));
 sky130_fd_sc_hd__or3_4 _25009_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_00372_));
 sky130_vsdinv _25010_ (.A(\mem_rdata_q[25] ),
    .Y(_18827_));
 sky130_vsdinv _25011_ (.A(_18210_),
    .Y(_18828_));
 sky130_fd_sc_hd__nand3_4 _25012_ (.A(mem_rdata[25]),
    .B(_18206_),
    .C(_18207_),
    .Y(_18829_));
 sky130_fd_sc_hd__o21ai_4 _25013_ (.A1(_18827_),
    .A2(_18828_),
    .B1(_18829_),
    .Y(\mem_rdata_latched[25] ));
 sky130_vsdinv _25014_ (.A(\mem_rdata_q[28] ),
    .Y(_18830_));
 sky130_fd_sc_hd__buf_1 _25015_ (.A(_18828_),
    .X(_18831_));
 sky130_fd_sc_hd__nand3_4 _25016_ (.A(mem_rdata[28]),
    .B(_18206_),
    .C(_18207_),
    .Y(_18832_));
 sky130_fd_sc_hd__o21ai_4 _25017_ (.A1(_18830_),
    .A2(_18831_),
    .B1(_18832_),
    .Y(\mem_rdata_latched[28] ));
 sky130_vsdinv _25018_ (.A(instr_sh),
    .Y(_18833_));
 sky130_fd_sc_hd__buf_1 _25019_ (.A(_18246_),
    .X(_18834_));
 sky130_fd_sc_hd__buf_1 _25020_ (.A(_18233_),
    .X(_18835_));
 sky130_fd_sc_hd__nand3_4 _25021_ (.A(_18834_),
    .B(_18243_),
    .C(_18835_),
    .Y(_18836_));
 sky130_fd_sc_hd__buf_1 _25022_ (.A(_18237_),
    .X(_18837_));
 sky130_fd_sc_hd__buf_1 _25023_ (.A(_18240_),
    .X(_18838_));
 sky130_fd_sc_hd__nand3_4 _25024_ (.A(_18837_),
    .B(_18234_),
    .C(_18838_),
    .Y(_18839_));
 sky130_fd_sc_hd__o22a_4 _25025_ (.A1(_18833_),
    .A2(_18836_),
    .B1(_18839_),
    .B2(_18324_),
    .X(_18840_));
 sky130_fd_sc_hd__buf_1 _25026_ (.A(_18295_),
    .X(_18841_));
 sky130_fd_sc_hd__buf_1 _25027_ (.A(_18841_),
    .X(_18842_));
 sky130_fd_sc_hd__buf_1 _25028_ (.A(_18234_),
    .X(_18843_));
 sky130_fd_sc_hd__nand3_4 _25029_ (.A(_18277_),
    .B(_18843_),
    .C(_18282_),
    .Y(_18844_));
 sky130_fd_sc_hd__a2bb2o_4 _25030_ (.A1_N(_18259_),
    .A2_N(_18840_),
    .B1(_18842_),
    .B2(_18844_),
    .X(_00668_));
 sky130_vsdinv _25031_ (.A(instr_sb),
    .Y(_18845_));
 sky130_fd_sc_hd__o22a_4 _25032_ (.A1(_18845_),
    .A2(_18836_),
    .B1(_18839_),
    .B2(_18323_),
    .X(_18846_));
 sky130_fd_sc_hd__buf_1 _25033_ (.A(\mem_wordsize[1] ),
    .X(_18847_));
 sky130_fd_sc_hd__buf_1 _25034_ (.A(_18258_),
    .X(_18848_));
 sky130_fd_sc_hd__buf_1 _25035_ (.A(_18266_),
    .X(_18849_));
 sky130_fd_sc_hd__buf_1 _25036_ (.A(_18849_),
    .X(_18850_));
 sky130_fd_sc_hd__buf_1 _25037_ (.A(_18850_),
    .X(_18851_));
 sky130_fd_sc_hd__nor3_4 _25038_ (.A(_18243_),
    .B(_18851_),
    .C(_18240_),
    .Y(_18852_));
 sky130_fd_sc_hd__and2_4 _25039_ (.A(_18279_),
    .B(_18281_),
    .X(_18853_));
 sky130_fd_sc_hd__a2111o_4 _25040_ (.A1(_18848_),
    .A2(_18518_),
    .B1(_18228_),
    .C1(_18852_),
    .D1(_18853_),
    .X(_18854_));
 sky130_fd_sc_hd__a2bb2o_4 _25041_ (.A1_N(_18259_),
    .A2_N(_18846_),
    .B1(_18847_),
    .B2(_18854_),
    .X(_00667_));
 sky130_fd_sc_hd__buf_1 _25042_ (.A(_18534_),
    .X(_18855_));
 sky130_fd_sc_hd__nand3_4 _25043_ (.A(_18789_),
    .B(_18855_),
    .C(_18808_),
    .Y(_18856_));
 sky130_fd_sc_hd__buf_1 _25044_ (.A(_18521_),
    .X(_18857_));
 sky130_fd_sc_hd__nor2_4 _25045_ (.A(_18290_),
    .B(_18796_),
    .Y(_18858_));
 sky130_fd_sc_hd__a32o_4 _25046_ (.A1(_18857_),
    .A2(_18399_),
    .A3(_18531_),
    .B1(_18508_),
    .B2(_18858_),
    .X(_18859_));
 sky130_fd_sc_hd__a2bb2o_4 _25047_ (.A1_N(_18317_),
    .A2_N(_18856_),
    .B1(_18391_),
    .B2(_18859_),
    .X(_18860_));
 sky130_fd_sc_hd__buf_1 _25048_ (.A(_18548_),
    .X(_18861_));
 sky130_fd_sc_hd__buf_1 _25049_ (.A(_18861_),
    .X(_18862_));
 sky130_fd_sc_hd__nor3_4 _25050_ (.A(_18529_),
    .B(_18522_),
    .C(_18489_),
    .Y(_18863_));
 sky130_fd_sc_hd__buf_1 _25051_ (.A(_18402_),
    .X(_18864_));
 sky130_fd_sc_hd__nor4_4 _25052_ (.A(_18864_),
    .B(_18857_),
    .C(_18394_),
    .D(_18475_),
    .Y(_18865_));
 sky130_fd_sc_hd__buf_1 _25053_ (.A(_18400_),
    .X(_18866_));
 sky130_fd_sc_hd__o21a_4 _25054_ (.A1(_18863_),
    .A2(_18865_),
    .B1(_18866_),
    .X(_18867_));
 sky130_vsdinv _25055_ (.A(_18858_),
    .Y(_18868_));
 sky130_fd_sc_hd__a21oi_4 _25056_ (.A1(_18369_),
    .A2(_18474_),
    .B1(_18868_),
    .Y(_18869_));
 sky130_fd_sc_hd__a211o_4 _25057_ (.A1(_18860_),
    .A2(_18862_),
    .B1(_18867_),
    .C1(_18869_),
    .X(_00663_));
 sky130_vsdinv _25058_ (.A(\mem_rdata_q[12] ),
    .Y(_18870_));
 sky130_fd_sc_hd__buf_1 _25059_ (.A(_18831_),
    .X(_18871_));
 sky130_fd_sc_hd__buf_1 _25060_ (.A(_18200_),
    .X(_18872_));
 sky130_fd_sc_hd__buf_1 _25061_ (.A(_18201_),
    .X(_18873_));
 sky130_fd_sc_hd__nand3_4 _25062_ (.A(mem_rdata[12]),
    .B(_18872_),
    .C(_18873_),
    .Y(_18874_));
 sky130_fd_sc_hd__o21ai_4 _25063_ (.A1(_18870_),
    .A2(_18871_),
    .B1(_18874_),
    .Y(\mem_rdata_latched[12] ));
 sky130_vsdinv _25064_ (.A(\mem_rdata_q[13] ),
    .Y(_18875_));
 sky130_fd_sc_hd__buf_1 _25065_ (.A(_18831_),
    .X(_18876_));
 sky130_fd_sc_hd__nand3_4 _25066_ (.A(mem_rdata[13]),
    .B(_18872_),
    .C(_18873_),
    .Y(_18877_));
 sky130_fd_sc_hd__o21ai_4 _25067_ (.A1(_18875_),
    .A2(_18876_),
    .B1(_18877_),
    .Y(\mem_rdata_latched[13] ));
 sky130_vsdinv _25068_ (.A(\mem_rdata_q[14] ),
    .Y(_18878_));
 sky130_fd_sc_hd__nand3_4 _25069_ (.A(mem_rdata[14]),
    .B(_18872_),
    .C(_18873_),
    .Y(_18879_));
 sky130_fd_sc_hd__o21ai_4 _25070_ (.A1(_18878_),
    .A2(_18876_),
    .B1(_18879_),
    .Y(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__nand3_4 _25071_ (.A(mem_rdata[29]),
    .B(_18193_),
    .C(_18195_),
    .Y(_18880_));
 sky130_fd_sc_hd__a21boi_4 _25072_ (.A1(\mem_rdata_q[29] ),
    .A2(_18191_),
    .B1_N(_18880_),
    .Y(_18881_));
 sky130_vsdinv _25073_ (.A(_18881_),
    .Y(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__nand3_4 _25074_ (.A(mem_rdata[30]),
    .B(_18192_),
    .C(_18194_),
    .Y(_18882_));
 sky130_fd_sc_hd__a21boi_4 _25075_ (.A1(\mem_rdata_q[30] ),
    .A2(_18190_),
    .B1_N(_18882_),
    .Y(_18883_));
 sky130_vsdinv _25076_ (.A(_18883_),
    .Y(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__nand3_4 _25077_ (.A(mem_rdata[31]),
    .B(_18192_),
    .C(_18194_),
    .Y(_18884_));
 sky130_fd_sc_hd__a21boi_4 _25078_ (.A1(\mem_rdata_q[31] ),
    .A2(_18190_),
    .B1_N(_18884_),
    .Y(_18885_));
 sky130_vsdinv _25079_ (.A(_18885_),
    .Y(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__buf_1 _25080_ (.A(\mem_state[0] ),
    .X(_18886_));
 sky130_vsdinv _25081_ (.A(_18886_),
    .Y(_18887_));
 sky130_vsdinv _25082_ (.A(\mem_state[1] ),
    .Y(_18888_));
 sky130_fd_sc_hd__nand4_4 _25083_ (.A(_18509_),
    .B(_18887_),
    .C(_18888_),
    .D(_18280_),
    .Y(_18889_));
 sky130_vsdinv _25084_ (.A(_18889_),
    .Y(_18890_));
 sky130_fd_sc_hd__buf_1 _25085_ (.A(_18890_),
    .X(mem_la_write));
 sky130_fd_sc_hd__buf_1 _25086_ (.A(mem_do_prefetch),
    .X(_18891_));
 sky130_fd_sc_hd__buf_1 _25087_ (.A(mem_do_rinst),
    .X(_18892_));
 sky130_fd_sc_hd__nor2_4 _25088_ (.A(_18891_),
    .B(_18892_),
    .Y(_18893_));
 sky130_fd_sc_hd__buf_1 _25089_ (.A(_18529_),
    .X(_18894_));
 sky130_fd_sc_hd__buf_1 _25090_ (.A(_18251_),
    .X(_18895_));
 sky130_vsdinv _25091_ (.A(_18895_),
    .Y(_18896_));
 sky130_fd_sc_hd__buf_1 _25092_ (.A(_18896_),
    .X(_18897_));
 sky130_fd_sc_hd__a211o_4 _25093_ (.A1(_18893_),
    .A2(_18837_),
    .B1(_18894_),
    .C1(_18897_),
    .X(_18898_));
 sky130_vsdinv _25094_ (.A(_18898_),
    .Y(mem_la_read));
 sky130_fd_sc_hd__nor3_4 _25095_ (.A(_18242_),
    .B(_18239_),
    .C(_18797_),
    .Y(_18899_));
 sky130_fd_sc_hd__buf_1 _25096_ (.A(_18899_),
    .X(_18900_));
 sky130_fd_sc_hd__nor3_4 _25097_ (.A(\cpu_state[4] ),
    .B(_18501_),
    .C(\cpu_state[0] ),
    .Y(_18901_));
 sky130_fd_sc_hd__buf_1 _25098_ (.A(_18901_),
    .X(_18902_));
 sky130_fd_sc_hd__buf_1 _25099_ (.A(\irq_state[1] ),
    .X(_18903_));
 sky130_fd_sc_hd__buf_1 _25100_ (.A(_18903_),
    .X(_18904_));
 sky130_fd_sc_hd__buf_1 _25101_ (.A(_18904_),
    .X(_18905_));
 sky130_fd_sc_hd__and4_4 _25102_ (.A(_18900_),
    .B(_18902_),
    .C(_18413_),
    .D(_18905_),
    .X(_18906_));
 sky130_fd_sc_hd__buf_1 _25103_ (.A(\irq_pending[0] ),
    .X(_18907_));
 sky130_fd_sc_hd__buf_1 _25104_ (.A(\timer[13] ),
    .X(_18908_));
 sky130_fd_sc_hd__nor4_4 _25105_ (.A(\timer[8] ),
    .B(\timer[11] ),
    .C(_18908_),
    .D(\timer[12] ),
    .Y(_18909_));
 sky130_fd_sc_hd__nor2_4 _25106_ (.A(\timer[9] ),
    .B(\timer[10] ),
    .Y(_18910_));
 sky130_fd_sc_hd__nor2_4 _25107_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .Y(_18911_));
 sky130_fd_sc_hd__buf_1 _25108_ (.A(_18911_),
    .X(_18912_));
 sky130_fd_sc_hd__and3_4 _25109_ (.A(_18909_),
    .B(_18910_),
    .C(_18912_),
    .X(_18913_));
 sky130_vsdinv _25110_ (.A(\timer[1] ),
    .Y(_18914_));
 sky130_vsdinv _25111_ (.A(\timer[2] ),
    .Y(_18915_));
 sky130_vsdinv _25112_ (.A(\timer[3] ),
    .Y(_18916_));
 sky130_fd_sc_hd__buf_1 _25113_ (.A(_18916_),
    .X(_18917_));
 sky130_fd_sc_hd__buf_1 _25114_ (.A(\timer[0] ),
    .X(_18918_));
 sky130_fd_sc_hd__and4_4 _25115_ (.A(_18914_),
    .B(_18915_),
    .C(_18917_),
    .D(_18918_),
    .X(_18919_));
 sky130_fd_sc_hd__nor4_4 _25116_ (.A(\timer[15] ),
    .B(\timer[14] ),
    .C(\timer[7] ),
    .D(\timer[6] ),
    .Y(_18920_));
 sky130_fd_sc_hd__and3_4 _25117_ (.A(_18913_),
    .B(_18919_),
    .C(_18920_),
    .X(_18921_));
 sky130_fd_sc_hd__nor4_4 _25118_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .C(\timer[31] ),
    .D(\timer[30] ),
    .Y(_18922_));
 sky130_fd_sc_hd__nor3_4 _25119_ (.A(\timer[17] ),
    .B(\timer[16] ),
    .C(\timer[18] ),
    .Y(_18923_));
 sky130_fd_sc_hd__nor3_4 _25120_ (.A(\timer[19] ),
    .B(\timer[23] ),
    .C(\timer[22] ),
    .Y(_18924_));
 sky130_fd_sc_hd__nor2_4 _25121_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .Y(_18925_));
 sky130_fd_sc_hd__and3_4 _25122_ (.A(_18923_),
    .B(_18924_),
    .C(_18925_),
    .X(_18926_));
 sky130_vsdinv _25123_ (.A(\timer[24] ),
    .Y(_18927_));
 sky130_vsdinv _25124_ (.A(\timer[27] ),
    .Y(_18928_));
 sky130_fd_sc_hd__nor2_4 _25125_ (.A(\timer[25] ),
    .B(\timer[26] ),
    .Y(_18929_));
 sky130_fd_sc_hd__and4_4 _25126_ (.A(_18926_),
    .B(_18927_),
    .C(_18928_),
    .D(_18929_),
    .X(_18930_));
 sky130_fd_sc_hd__buf_1 _25127_ (.A(_18930_),
    .X(_18931_));
 sky130_fd_sc_hd__and3_4 _25128_ (.A(_18921_),
    .B(_18922_),
    .C(_18931_),
    .X(_18932_));
 sky130_fd_sc_hd__nor3_4 _25129_ (.A(_18907_),
    .B(irq[0]),
    .C(_18932_),
    .Y(_18933_));
 sky130_fd_sc_hd__nor3_4 _25130_ (.A(_18784_),
    .B(_18906_),
    .C(_18933_),
    .Y(_00328_));
 sky130_fd_sc_hd__buf_1 _25131_ (.A(_18783_),
    .X(_18934_));
 sky130_fd_sc_hd__buf_1 _25132_ (.A(\irq_pending[1] ),
    .X(_18935_));
 sky130_fd_sc_hd__buf_1 _25133_ (.A(_18904_),
    .X(_18936_));
 sky130_fd_sc_hd__a2bb2o_4 _25134_ (.A1_N(_18935_),
    .A2_N(irq[1]),
    .B1(_18410_),
    .B2(_18936_),
    .X(_18937_));
 sky130_fd_sc_hd__and3_4 _25135_ (.A(_18937_),
    .B(_18900_),
    .C(_18902_),
    .X(_18938_));
 sky130_fd_sc_hd__and4_4 _25136_ (.A(_18497_),
    .B(_18855_),
    .C(_18503_),
    .D(_18492_),
    .X(_18939_));
 sky130_fd_sc_hd__nor3_4 _25137_ (.A(_18935_),
    .B(irq[1]),
    .C(_18939_),
    .Y(_18940_));
 sky130_fd_sc_hd__nor3_4 _25138_ (.A(_18934_),
    .B(_18938_),
    .C(_18940_),
    .Y(_00339_));
 sky130_fd_sc_hd__buf_1 _25139_ (.A(_18900_),
    .X(_18941_));
 sky130_fd_sc_hd__buf_1 _25140_ (.A(_18902_),
    .X(_18942_));
 sky130_fd_sc_hd__buf_1 _25141_ (.A(_18905_),
    .X(_18943_));
 sky130_fd_sc_hd__nand4_4 _25142_ (.A(_18429_),
    .B(_18941_),
    .C(_18942_),
    .D(_18943_),
    .Y(_18944_));
 sky130_fd_sc_hd__buf_1 _25143_ (.A(_18507_),
    .X(_18945_));
 sky130_fd_sc_hd__buf_1 _25144_ (.A(\irq_pending[3] ),
    .X(_18946_));
 sky130_fd_sc_hd__or2_4 _25145_ (.A(_18946_),
    .B(irq[3]),
    .X(_18947_));
 sky130_fd_sc_hd__and3_4 _25146_ (.A(_18944_),
    .B(_18945_),
    .C(_18947_),
    .X(_00353_));
 sky130_fd_sc_hd__nand4_4 _25147_ (.A(_18419_),
    .B(_18941_),
    .C(_18942_),
    .D(_18943_),
    .Y(_18948_));
 sky130_fd_sc_hd__or2_4 _25148_ (.A(\irq_pending[4] ),
    .B(irq[4]),
    .X(_18949_));
 sky130_fd_sc_hd__and3_4 _25149_ (.A(_18948_),
    .B(_18945_),
    .C(_18949_),
    .X(_00354_));
 sky130_fd_sc_hd__nand4_4 _25150_ (.A(_18432_),
    .B(_18941_),
    .C(_18942_),
    .D(_18943_),
    .Y(_18950_));
 sky130_fd_sc_hd__or2_4 _25151_ (.A(\irq_pending[5] ),
    .B(irq[5]),
    .X(_18951_));
 sky130_fd_sc_hd__and3_4 _25152_ (.A(_18950_),
    .B(_18945_),
    .C(_18951_),
    .X(_00355_));
 sky130_fd_sc_hd__buf_1 _25153_ (.A(_18904_),
    .X(_18952_));
 sky130_fd_sc_hd__buf_1 _25154_ (.A(_18952_),
    .X(_18953_));
 sky130_fd_sc_hd__nand4_4 _25155_ (.A(_18414_),
    .B(_18941_),
    .C(_18942_),
    .D(_18953_),
    .Y(_18954_));
 sky130_fd_sc_hd__or2_4 _25156_ (.A(\irq_pending[6] ),
    .B(irq[6]),
    .X(_18955_));
 sky130_fd_sc_hd__and3_4 _25157_ (.A(_18954_),
    .B(_18945_),
    .C(_18955_),
    .X(_00356_));
 sky130_fd_sc_hd__buf_1 _25158_ (.A(_18899_),
    .X(_18956_));
 sky130_fd_sc_hd__buf_1 _25159_ (.A(_18956_),
    .X(_18957_));
 sky130_fd_sc_hd__buf_1 _25160_ (.A(_18957_),
    .X(_18958_));
 sky130_fd_sc_hd__buf_1 _25161_ (.A(_18901_),
    .X(_18959_));
 sky130_fd_sc_hd__buf_1 _25162_ (.A(_18959_),
    .X(_18960_));
 sky130_fd_sc_hd__buf_1 _25163_ (.A(_18960_),
    .X(_18961_));
 sky130_fd_sc_hd__nand4_4 _25164_ (.A(_18430_),
    .B(_18958_),
    .C(_18961_),
    .D(_18953_),
    .Y(_18962_));
 sky130_fd_sc_hd__buf_1 _25165_ (.A(_18548_),
    .X(_18963_));
 sky130_fd_sc_hd__buf_1 _25166_ (.A(_18963_),
    .X(_18964_));
 sky130_fd_sc_hd__or2_4 _25167_ (.A(\irq_pending[7] ),
    .B(irq[7]),
    .X(_18965_));
 sky130_fd_sc_hd__and3_4 _25168_ (.A(_18962_),
    .B(_18964_),
    .C(_18965_),
    .X(_00357_));
 sky130_fd_sc_hd__nand4_4 _25169_ (.A(_18436_),
    .B(_18958_),
    .C(_18961_),
    .D(_18953_),
    .Y(_18966_));
 sky130_fd_sc_hd__or2_4 _25170_ (.A(\irq_pending[8] ),
    .B(irq[8]),
    .X(_18967_));
 sky130_fd_sc_hd__and3_4 _25171_ (.A(_18966_),
    .B(_18964_),
    .C(_18967_),
    .X(_00358_));
 sky130_fd_sc_hd__nand4_4 _25172_ (.A(_18411_),
    .B(_18958_),
    .C(_18961_),
    .D(_18953_),
    .Y(_18968_));
 sky130_fd_sc_hd__or2_4 _25173_ (.A(\irq_pending[9] ),
    .B(irq[9]),
    .X(_18969_));
 sky130_fd_sc_hd__and3_4 _25174_ (.A(_18968_),
    .B(_18964_),
    .C(_18969_),
    .X(_00359_));
 sky130_fd_sc_hd__buf_1 _25175_ (.A(_18952_),
    .X(_18970_));
 sky130_fd_sc_hd__nand4_4 _25176_ (.A(_18417_),
    .B(_18958_),
    .C(_18961_),
    .D(_18970_),
    .Y(_18971_));
 sky130_fd_sc_hd__or2_4 _25177_ (.A(\irq_pending[10] ),
    .B(irq[10]),
    .X(_18972_));
 sky130_fd_sc_hd__and3_4 _25178_ (.A(_18971_),
    .B(_18964_),
    .C(_18972_),
    .X(_00329_));
 sky130_fd_sc_hd__buf_1 _25179_ (.A(_18957_),
    .X(_18973_));
 sky130_fd_sc_hd__buf_1 _25180_ (.A(_18960_),
    .X(_18974_));
 sky130_fd_sc_hd__nand4_4 _25181_ (.A(_18439_),
    .B(_18973_),
    .C(_18974_),
    .D(_18970_),
    .Y(_18975_));
 sky130_fd_sc_hd__buf_1 _25182_ (.A(_18963_),
    .X(_18976_));
 sky130_fd_sc_hd__or2_4 _25183_ (.A(\irq_pending[11] ),
    .B(irq[11]),
    .X(_18977_));
 sky130_fd_sc_hd__and3_4 _25184_ (.A(_18975_),
    .B(_18976_),
    .C(_18977_),
    .X(_00330_));
 sky130_fd_sc_hd__nand4_4 _25185_ (.A(_18423_),
    .B(_18973_),
    .C(_18974_),
    .D(_18970_),
    .Y(_18978_));
 sky130_fd_sc_hd__or2_4 _25186_ (.A(\irq_pending[12] ),
    .B(irq[12]),
    .X(_18979_));
 sky130_fd_sc_hd__and3_4 _25187_ (.A(_18978_),
    .B(_18976_),
    .C(_18979_),
    .X(_00331_));
 sky130_fd_sc_hd__nand4_4 _25188_ (.A(_18445_),
    .B(_18973_),
    .C(_18974_),
    .D(_18970_),
    .Y(_18980_));
 sky130_fd_sc_hd__or2_4 _25189_ (.A(\irq_pending[13] ),
    .B(irq[13]),
    .X(_18981_));
 sky130_fd_sc_hd__and3_4 _25190_ (.A(_18980_),
    .B(_18976_),
    .C(_18981_),
    .X(_00332_));
 sky130_fd_sc_hd__buf_1 _25191_ (.A(_18952_),
    .X(_18982_));
 sky130_fd_sc_hd__nand4_4 _25192_ (.A(_18437_),
    .B(_18973_),
    .C(_18974_),
    .D(_18982_),
    .Y(_18983_));
 sky130_fd_sc_hd__or2_4 _25193_ (.A(\irq_pending[14] ),
    .B(irq[14]),
    .X(_18984_));
 sky130_fd_sc_hd__and3_4 _25194_ (.A(_18983_),
    .B(_18976_),
    .C(_18984_),
    .X(_00333_));
 sky130_fd_sc_hd__buf_1 _25195_ (.A(_18957_),
    .X(_18985_));
 sky130_fd_sc_hd__buf_1 _25196_ (.A(_18960_),
    .X(_18986_));
 sky130_fd_sc_hd__nand4_4 _25197_ (.A(_18442_),
    .B(_18985_),
    .C(_18986_),
    .D(_18982_),
    .Y(_18987_));
 sky130_fd_sc_hd__buf_1 _25198_ (.A(_18963_),
    .X(_18988_));
 sky130_fd_sc_hd__or2_4 _25199_ (.A(\irq_pending[15] ),
    .B(irq[15]),
    .X(_18989_));
 sky130_fd_sc_hd__and3_4 _25200_ (.A(_18987_),
    .B(_18988_),
    .C(_18989_),
    .X(_00334_));
 sky130_fd_sc_hd__nand4_4 _25201_ (.A(_18433_),
    .B(_18985_),
    .C(_18986_),
    .D(_18982_),
    .Y(_18990_));
 sky130_fd_sc_hd__or2_4 _25202_ (.A(\irq_pending[16] ),
    .B(irq[16]),
    .X(_18991_));
 sky130_fd_sc_hd__and3_4 _25203_ (.A(_18990_),
    .B(_18988_),
    .C(_18991_),
    .X(_00335_));
 sky130_fd_sc_hd__nand4_4 _25204_ (.A(_18449_),
    .B(_18985_),
    .C(_18986_),
    .D(_18982_),
    .Y(_18992_));
 sky130_fd_sc_hd__or2_4 _25205_ (.A(\irq_pending[17] ),
    .B(irq[17]),
    .X(_18993_));
 sky130_fd_sc_hd__and3_4 _25206_ (.A(_18992_),
    .B(_18988_),
    .C(_18993_),
    .X(_00336_));
 sky130_fd_sc_hd__buf_1 _25207_ (.A(_18952_),
    .X(_18994_));
 sky130_fd_sc_hd__nand4_4 _25208_ (.A(_18450_),
    .B(_18985_),
    .C(_18986_),
    .D(_18994_),
    .Y(_18995_));
 sky130_fd_sc_hd__or2_4 _25209_ (.A(\irq_pending[18] ),
    .B(irq[18]),
    .X(_18996_));
 sky130_fd_sc_hd__and3_4 _25210_ (.A(_18995_),
    .B(_18988_),
    .C(_18996_),
    .X(_00337_));
 sky130_fd_sc_hd__buf_1 _25211_ (.A(_18957_),
    .X(_18997_));
 sky130_fd_sc_hd__buf_1 _25212_ (.A(_18960_),
    .X(_18998_));
 sky130_fd_sc_hd__nand4_4 _25213_ (.A(_18426_),
    .B(_18997_),
    .C(_18998_),
    .D(_18994_),
    .Y(_18999_));
 sky130_fd_sc_hd__buf_1 _25214_ (.A(_18963_),
    .X(_19000_));
 sky130_fd_sc_hd__or2_4 _25215_ (.A(\irq_pending[19] ),
    .B(irq[19]),
    .X(_19001_));
 sky130_fd_sc_hd__and3_4 _25216_ (.A(_18999_),
    .B(_19000_),
    .C(_19001_),
    .X(_00338_));
 sky130_fd_sc_hd__nand4_4 _25217_ (.A(_18440_),
    .B(_18997_),
    .C(_18998_),
    .D(_18994_),
    .Y(_19002_));
 sky130_fd_sc_hd__or2_4 _25218_ (.A(\irq_pending[20] ),
    .B(irq[20]),
    .X(_19003_));
 sky130_fd_sc_hd__and3_4 _25219_ (.A(_19002_),
    .B(_19000_),
    .C(_19003_),
    .X(_00340_));
 sky130_fd_sc_hd__nand4_4 _25220_ (.A(_18443_),
    .B(_18997_),
    .C(_18998_),
    .D(_18994_),
    .Y(_19004_));
 sky130_fd_sc_hd__or2_4 _25221_ (.A(\irq_pending[21] ),
    .B(irq[21]),
    .X(_19005_));
 sky130_fd_sc_hd__and3_4 _25222_ (.A(_19004_),
    .B(_19000_),
    .C(_19005_),
    .X(_00341_));
 sky130_fd_sc_hd__buf_1 _25223_ (.A(_18936_),
    .X(_19006_));
 sky130_fd_sc_hd__nand4_4 _25224_ (.A(_18427_),
    .B(_18997_),
    .C(_18998_),
    .D(_19006_),
    .Y(_19007_));
 sky130_fd_sc_hd__or2_4 _25225_ (.A(\irq_pending[22] ),
    .B(irq[22]),
    .X(_19008_));
 sky130_fd_sc_hd__and3_4 _25226_ (.A(_19007_),
    .B(_19000_),
    .C(_19008_),
    .X(_00342_));
 sky130_fd_sc_hd__buf_1 _25227_ (.A(_18956_),
    .X(_19009_));
 sky130_fd_sc_hd__buf_1 _25228_ (.A(_18959_),
    .X(_19010_));
 sky130_fd_sc_hd__nand4_4 _25229_ (.A(_18424_),
    .B(_19009_),
    .C(_19010_),
    .D(_19006_),
    .Y(_19011_));
 sky130_fd_sc_hd__buf_1 _25230_ (.A(_18506_),
    .X(_19012_));
 sky130_fd_sc_hd__buf_1 _25231_ (.A(_19012_),
    .X(_19013_));
 sky130_fd_sc_hd__or2_4 _25232_ (.A(\irq_pending[23] ),
    .B(irq[23]),
    .X(_19014_));
 sky130_fd_sc_hd__and3_4 _25233_ (.A(_19011_),
    .B(_19013_),
    .C(_19014_),
    .X(_00343_));
 sky130_fd_sc_hd__nand4_4 _25234_ (.A(_18458_),
    .B(_19009_),
    .C(_19010_),
    .D(_19006_),
    .Y(_19015_));
 sky130_fd_sc_hd__or2_4 _25235_ (.A(\irq_pending[24] ),
    .B(irq[24]),
    .X(_19016_));
 sky130_fd_sc_hd__and3_4 _25236_ (.A(_19015_),
    .B(_19013_),
    .C(_19016_),
    .X(_00344_));
 sky130_fd_sc_hd__nand4_4 _25237_ (.A(_18452_),
    .B(_19009_),
    .C(_19010_),
    .D(_19006_),
    .Y(_19017_));
 sky130_fd_sc_hd__or2_4 _25238_ (.A(\irq_pending[25] ),
    .B(irq[25]),
    .X(_19018_));
 sky130_fd_sc_hd__and3_4 _25239_ (.A(_19017_),
    .B(_19013_),
    .C(_19018_),
    .X(_00345_));
 sky130_fd_sc_hd__buf_1 _25240_ (.A(_18936_),
    .X(_19019_));
 sky130_fd_sc_hd__nand4_4 _25241_ (.A(_18453_),
    .B(_19009_),
    .C(_19010_),
    .D(_19019_),
    .Y(_19020_));
 sky130_fd_sc_hd__or2_4 _25242_ (.A(\irq_pending[26] ),
    .B(irq[26]),
    .X(_19021_));
 sky130_fd_sc_hd__and3_4 _25243_ (.A(_19020_),
    .B(_19013_),
    .C(_19021_),
    .X(_00346_));
 sky130_fd_sc_hd__buf_1 _25244_ (.A(_18956_),
    .X(_19022_));
 sky130_fd_sc_hd__buf_1 _25245_ (.A(_18959_),
    .X(_19023_));
 sky130_fd_sc_hd__nand4_4 _25246_ (.A(_18455_),
    .B(_19022_),
    .C(_19023_),
    .D(_19019_),
    .Y(_19024_));
 sky130_fd_sc_hd__buf_1 _25247_ (.A(_19012_),
    .X(_19025_));
 sky130_fd_sc_hd__or2_4 _25248_ (.A(\irq_pending[27] ),
    .B(irq[27]),
    .X(_19026_));
 sky130_fd_sc_hd__and3_4 _25249_ (.A(_19024_),
    .B(_19025_),
    .C(_19026_),
    .X(_00347_));
 sky130_fd_sc_hd__nand4_4 _25250_ (.A(_18446_),
    .B(_19022_),
    .C(_19023_),
    .D(_19019_),
    .Y(_19027_));
 sky130_fd_sc_hd__or2_4 _25251_ (.A(\irq_pending[28] ),
    .B(irq[28]),
    .X(_19028_));
 sky130_fd_sc_hd__and3_4 _25252_ (.A(_19027_),
    .B(_19025_),
    .C(_19028_),
    .X(_00348_));
 sky130_fd_sc_hd__nand4_4 _25253_ (.A(_18420_),
    .B(_19022_),
    .C(_19023_),
    .D(_19019_),
    .Y(_19029_));
 sky130_fd_sc_hd__or2_4 _25254_ (.A(\irq_pending[29] ),
    .B(irq[29]),
    .X(_19030_));
 sky130_fd_sc_hd__and3_4 _25255_ (.A(_19029_),
    .B(_19025_),
    .C(_19030_),
    .X(_00349_));
 sky130_fd_sc_hd__nand4_4 _25256_ (.A(_18456_),
    .B(_19022_),
    .C(_19023_),
    .D(_18905_),
    .Y(_19031_));
 sky130_fd_sc_hd__or2_4 _25257_ (.A(\irq_pending[30] ),
    .B(irq[30]),
    .X(_19032_));
 sky130_fd_sc_hd__and3_4 _25258_ (.A(_19031_),
    .B(_19025_),
    .C(_19032_),
    .X(_00351_));
 sky130_fd_sc_hd__nand4_4 _25259_ (.A(_18459_),
    .B(_18900_),
    .C(_18902_),
    .D(_18905_),
    .Y(_19033_));
 sky130_fd_sc_hd__buf_1 _25260_ (.A(_19012_),
    .X(_19034_));
 sky130_fd_sc_hd__or2_4 _25261_ (.A(\irq_pending[31] ),
    .B(irq[31]),
    .X(_19035_));
 sky130_fd_sc_hd__and3_4 _25262_ (.A(_19033_),
    .B(_19034_),
    .C(_19035_),
    .X(_00352_));
 sky130_vsdinv _25263_ (.A(_18398_),
    .Y(_19036_));
 sky130_fd_sc_hd__buf_1 _25264_ (.A(_19036_),
    .X(_19037_));
 sky130_fd_sc_hd__buf_1 _25265_ (.A(_19037_),
    .X(_19038_));
 sky130_vsdinv _25266_ (.A(instr_bne),
    .Y(_19039_));
 sky130_fd_sc_hd__nand2_4 _25267_ (.A(_19039_),
    .B(alu_eq),
    .Y(_19040_));
 sky130_fd_sc_hd__nand2_4 _25268_ (.A(_18329_),
    .B(_18330_),
    .Y(_19041_));
 sky130_fd_sc_hd__or4_4 _25269_ (.A(is_slti_blt_slt),
    .B(is_sltiu_bltu_sltu),
    .C(_19040_),
    .D(_19041_),
    .X(_19042_));
 sky130_fd_sc_hd__a2bb2oi_4 _25270_ (.A1_N(alu_lts),
    .A2_N(_18330_),
    .B1(is_sltiu_bltu_sltu),
    .B2(alu_ltu),
    .Y(_19043_));
 sky130_fd_sc_hd__or2_4 _25271_ (.A(alu_ltu),
    .B(_18329_),
    .X(_19044_));
 sky130_fd_sc_hd__a2bb2oi_4 _25272_ (.A1_N(alu_eq),
    .A2_N(_19039_),
    .B1(is_slti_blt_slt),
    .B2(alu_lts),
    .Y(_19045_));
 sky130_fd_sc_hd__nand4_4 _25273_ (.A(_19042_),
    .B(_19043_),
    .C(_19044_),
    .D(_19045_),
    .Y(_19046_));
 sky130_fd_sc_hd__nand2_4 _25274_ (.A(_19046_),
    .B(_18403_),
    .Y(_19047_));
 sky130_fd_sc_hd__buf_1 _25275_ (.A(_18892_),
    .X(_19048_));
 sky130_fd_sc_hd__nand3_4 _25276_ (.A(_18275_),
    .B(_18232_),
    .C(_19048_),
    .Y(_19049_));
 sky130_vsdinv _25277_ (.A(_19049_),
    .Y(_19050_));
 sky130_fd_sc_hd__buf_1 _25278_ (.A(_19050_),
    .X(_19051_));
 sky130_fd_sc_hd__buf_1 _25279_ (.A(_19051_),
    .X(_19052_));
 sky130_fd_sc_hd__o32a_4 _25280_ (.A1(_19038_),
    .A2(_18518_),
    .A3(_19047_),
    .B1(_00211_),
    .B2(_19052_),
    .X(_00212_));
 sky130_fd_sc_hd__buf_1 _25281_ (.A(\pcpi_timeout_counter[0] ),
    .X(_19053_));
 sky130_fd_sc_hd__nor3_4 _25282_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .C(\pcpi_timeout_counter[2] ),
    .Y(_19054_));
 sky130_vsdinv _25283_ (.A(\pcpi_timeout_counter[3] ),
    .Y(_19055_));
 sky130_fd_sc_hd__nand2_4 _25284_ (.A(_19054_),
    .B(_19055_),
    .Y(_19056_));
 sky130_vsdinv _25285_ (.A(_19056_),
    .Y(_19057_));
 sky130_vsdinv _25286_ (.A(_18810_),
    .Y(_19058_));
 sky130_fd_sc_hd__o21a_4 _25287_ (.A1(_19053_),
    .A2(_19057_),
    .B1(_19058_),
    .X(_19059_));
 sky130_fd_sc_hd__buf_1 _25288_ (.A(_19055_),
    .X(_19060_));
 sky130_fd_sc_hd__nand3_4 _25289_ (.A(_19054_),
    .B(_19053_),
    .C(_19060_),
    .Y(_19061_));
 sky130_fd_sc_hd__nand2_4 _25290_ (.A(_19059_),
    .B(_19061_),
    .Y(_00493_));
 sky130_fd_sc_hd__buf_1 _25291_ (.A(\pcpi_timeout_counter[1] ),
    .X(_19062_));
 sky130_fd_sc_hd__nor2_4 _25292_ (.A(_19062_),
    .B(_19053_),
    .Y(_19063_));
 sky130_fd_sc_hd__a21oi_4 _25293_ (.A1(_19062_),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_18810_),
    .Y(_19064_));
 sky130_fd_sc_hd__a21bo_4 _25294_ (.A1(_19056_),
    .A2(_19063_),
    .B1_N(_19064_),
    .X(_00494_));
 sky130_fd_sc_hd__or4_4 _25295_ (.A(_19062_),
    .B(\pcpi_timeout_counter[0] ),
    .C(\pcpi_timeout_counter[2] ),
    .D(_19060_),
    .X(_19065_));
 sky130_fd_sc_hd__o21ai_4 _25296_ (.A1(_19062_),
    .A2(_19053_),
    .B1(\pcpi_timeout_counter[2] ),
    .Y(_19066_));
 sky130_fd_sc_hd__nand3_4 _25297_ (.A(_19065_),
    .B(_19058_),
    .C(_19066_),
    .Y(_00495_));
 sky130_fd_sc_hd__o21ai_4 _25298_ (.A1(_19060_),
    .A2(_19054_),
    .B1(_19058_),
    .Y(_00496_));
 sky130_vsdinv _25299_ (.A(\latched_rd[0] ),
    .Y(_19067_));
 sky130_fd_sc_hd__buf_1 _25300_ (.A(_19067_),
    .X(_19068_));
 sky130_fd_sc_hd__buf_1 _25301_ (.A(_19068_),
    .X(_19069_));
 sky130_fd_sc_hd__buf_1 _25302_ (.A(_18849_),
    .X(_19070_));
 sky130_fd_sc_hd__o21a_4 _25303_ (.A1(_19070_),
    .A2(_18398_),
    .B1(_18289_),
    .X(_19071_));
 sky130_fd_sc_hd__o21a_4 _25304_ (.A1(_19036_),
    .A2(_18403_),
    .B1(_19071_),
    .X(_19072_));
 sky130_fd_sc_hd__and2_4 _25305_ (.A(_19072_),
    .B(_18249_),
    .X(_19073_));
 sky130_fd_sc_hd__buf_1 _25306_ (.A(_19073_),
    .X(_19074_));
 sky130_fd_sc_hd__buf_1 _25307_ (.A(_18576_),
    .X(_19075_));
 sky130_fd_sc_hd__buf_1 _25308_ (.A(_18466_),
    .X(_19076_));
 sky130_fd_sc_hd__buf_1 _25309_ (.A(_19076_),
    .X(_19077_));
 sky130_fd_sc_hd__buf_1 _25310_ (.A(_19077_),
    .X(_19078_));
 sky130_fd_sc_hd__a21o_4 _25311_ (.A1(_19075_),
    .A2(\decoded_rd[0] ),
    .B1(_19078_),
    .X(_19079_));
 sky130_fd_sc_hd__a2bb2o_4 _25312_ (.A1_N(_19069_),
    .A2_N(_19074_),
    .B1(_18262_),
    .B2(_19079_),
    .X(_00377_));
 sky130_fd_sc_hd__buf_1 _25313_ (.A(_18267_),
    .X(_19080_));
 sky130_fd_sc_hd__buf_1 _25314_ (.A(_19080_),
    .X(_19081_));
 sky130_fd_sc_hd__buf_1 _25315_ (.A(_19081_),
    .X(_19082_));
 sky130_vsdinv _25316_ (.A(\decoded_rd[1] ),
    .Y(_19083_));
 sky130_fd_sc_hd__buf_1 _25317_ (.A(_18470_),
    .X(_19084_));
 sky130_vsdinv _25318_ (.A(\latched_rd[1] ),
    .Y(_19085_));
 sky130_fd_sc_hd__buf_1 _25319_ (.A(_19085_),
    .X(_19086_));
 sky130_fd_sc_hd__buf_1 _25320_ (.A(_19086_),
    .X(_19087_));
 sky130_fd_sc_hd__o32ai_4 _25321_ (.A1(_19082_),
    .A2(_19083_),
    .A3(_19084_),
    .B1(_19087_),
    .B2(_19074_),
    .Y(_00378_));
 sky130_vsdinv _25322_ (.A(\decoded_rd[2] ),
    .Y(_19088_));
 sky130_fd_sc_hd__buf_1 _25323_ (.A(\latched_rd[2] ),
    .X(_19089_));
 sky130_vsdinv _25324_ (.A(_19089_),
    .Y(_19090_));
 sky130_fd_sc_hd__o32ai_4 _25325_ (.A1(_19082_),
    .A2(_19088_),
    .A3(_19084_),
    .B1(_19090_),
    .B2(_19074_),
    .Y(_00379_));
 sky130_fd_sc_hd__buf_1 _25326_ (.A(_18479_),
    .X(_19091_));
 sky130_fd_sc_hd__buf_1 _25327_ (.A(_19091_),
    .X(_19092_));
 sky130_vsdinv _25328_ (.A(\decoded_rd[3] ),
    .Y(_19093_));
 sky130_fd_sc_hd__buf_1 _25329_ (.A(\latched_rd[3] ),
    .X(_19094_));
 sky130_vsdinv _25330_ (.A(_19094_),
    .Y(_19095_));
 sky130_fd_sc_hd__o32ai_4 _25331_ (.A1(_19092_),
    .A2(_19093_),
    .A3(_19084_),
    .B1(_19095_),
    .B2(_19074_),
    .Y(_00380_));
 sky130_fd_sc_hd__buf_1 _25332_ (.A(instr_setq),
    .X(_19096_));
 sky130_fd_sc_hd__buf_1 _25333_ (.A(_18798_),
    .X(_19097_));
 sky130_fd_sc_hd__buf_1 _25334_ (.A(\latched_rd[4] ),
    .X(_19098_));
 sky130_fd_sc_hd__a21oi_4 _25335_ (.A1(_19096_),
    .A2(_19097_),
    .B1(_19098_),
    .Y(_19099_));
 sky130_fd_sc_hd__buf_1 _25336_ (.A(_19070_),
    .X(_19100_));
 sky130_fd_sc_hd__buf_1 _25337_ (.A(_19100_),
    .X(_19101_));
 sky130_fd_sc_hd__buf_1 _25338_ (.A(_19101_),
    .X(_19102_));
 sky130_fd_sc_hd__buf_1 _25339_ (.A(_18778_),
    .X(_19103_));
 sky130_fd_sc_hd__buf_1 _25340_ (.A(_19103_),
    .X(_19104_));
 sky130_vsdinv _25341_ (.A(\decoded_rd[4] ),
    .Y(_19105_));
 sky130_fd_sc_hd__buf_1 _25342_ (.A(_18544_),
    .X(_19106_));
 sky130_fd_sc_hd__buf_1 _25343_ (.A(_19106_),
    .X(_19107_));
 sky130_fd_sc_hd__nand3_4 _25344_ (.A(_19104_),
    .B(_19105_),
    .C(_19107_),
    .Y(_19108_));
 sky130_fd_sc_hd__a2bb2oi_4 _25345_ (.A1_N(_19072_),
    .A2_N(_19099_),
    .B1(_19102_),
    .B2(_19108_),
    .Y(_19109_));
 sky130_fd_sc_hd__nand2_4 _25346_ (.A(_18286_),
    .B(_19098_),
    .Y(_19110_));
 sky130_fd_sc_hd__o21ai_4 _25347_ (.A1(_18784_),
    .A2(_19109_),
    .B1(_19110_),
    .Y(_00381_));
 sky130_fd_sc_hd__buf_1 _25348_ (.A(_18249_),
    .X(_19111_));
 sky130_fd_sc_hd__buf_1 _25349_ (.A(_19111_),
    .X(_19112_));
 sky130_fd_sc_hd__buf_1 _25350_ (.A(_19103_),
    .X(_19113_));
 sky130_fd_sc_hd__buf_1 _25351_ (.A(_18850_),
    .X(_19114_));
 sky130_fd_sc_hd__buf_1 _25352_ (.A(_19114_),
    .X(_19115_));
 sky130_fd_sc_hd__buf_1 _25353_ (.A(_19115_),
    .X(_19116_));
 sky130_fd_sc_hd__buf_1 _25354_ (.A(latched_compr),
    .X(_19117_));
 sky130_vsdinv _25355_ (.A(_19117_),
    .Y(_19118_));
 sky130_fd_sc_hd__a41oi_4 _25356_ (.A1(_19112_),
    .A2(_19113_),
    .A3(_19116_),
    .A4(_19107_),
    .B1(_19118_),
    .Y(_00374_));
 sky130_fd_sc_hd__or2_4 _25357_ (.A(_18482_),
    .B(_19113_),
    .X(_19119_));
 sky130_fd_sc_hd__buf_1 _25358_ (.A(_19070_),
    .X(_19120_));
 sky130_fd_sc_hd__buf_1 _25359_ (.A(_19120_),
    .X(_19121_));
 sky130_fd_sc_hd__buf_1 _25360_ (.A(_19121_),
    .X(_19122_));
 sky130_fd_sc_hd__buf_1 _25361_ (.A(_19122_),
    .X(_19123_));
 sky130_fd_sc_hd__buf_1 _25362_ (.A(_18509_),
    .X(_19124_));
 sky130_fd_sc_hd__buf_1 _25363_ (.A(_19124_),
    .X(_19125_));
 sky130_fd_sc_hd__buf_1 _25364_ (.A(_19125_),
    .X(_19126_));
 sky130_fd_sc_hd__o21ai_4 _25365_ (.A1(_19116_),
    .A2(_19078_),
    .B1(_19126_),
    .Y(_19127_));
 sky130_fd_sc_hd__a21oi_4 _25366_ (.A1(_19119_),
    .A2(_19123_),
    .B1(_19127_),
    .Y(_00360_));
 sky130_vsdinv _25367_ (.A(\irq_state[1] ),
    .Y(_19128_));
 sky130_fd_sc_hd__buf_1 _25368_ (.A(_19128_),
    .X(_19129_));
 sky130_fd_sc_hd__nand2_4 _25369_ (.A(_19121_),
    .B(_19078_),
    .Y(_19130_));
 sky130_fd_sc_hd__buf_1 _25370_ (.A(_18478_),
    .X(_19131_));
 sky130_fd_sc_hd__a21o_4 _25371_ (.A1(_19102_),
    .A2(_18943_),
    .B1(_19131_),
    .X(_19132_));
 sky130_fd_sc_hd__a21oi_4 _25372_ (.A1(_19129_),
    .A2(_19130_),
    .B1(_19132_),
    .Y(_00361_));
 sky130_vsdinv _25373_ (.A(decoder_trigger),
    .Y(_19133_));
 sky130_fd_sc_hd__buf_1 _25374_ (.A(_19133_),
    .X(_19134_));
 sky130_fd_sc_hd__buf_1 _25375_ (.A(_19134_),
    .X(_19135_));
 sky130_fd_sc_hd__buf_1 _25376_ (.A(_18404_),
    .X(_19136_));
 sky130_fd_sc_hd__nand3_4 _25377_ (.A(_18464_),
    .B(_18266_),
    .C(_18467_),
    .Y(_19137_));
 sky130_fd_sc_hd__buf_1 _25378_ (.A(_19137_),
    .X(_19138_));
 sky130_fd_sc_hd__nor4_4 _25379_ (.A(_18775_),
    .B(_19135_),
    .C(_19136_),
    .D(_19138_),
    .Y(_19139_));
 sky130_vsdinv _25380_ (.A(_19139_),
    .Y(_19140_));
 sky130_fd_sc_hd__buf_1 _25381_ (.A(instr_retirq),
    .X(_19141_));
 sky130_fd_sc_hd__buf_1 _25382_ (.A(instr_jalr),
    .X(_19142_));
 sky130_fd_sc_hd__o21a_4 _25383_ (.A1(_19141_),
    .A2(_19142_),
    .B1(_19139_),
    .X(_19143_));
 sky130_fd_sc_hd__a211o_4 _25384_ (.A1(_18361_),
    .A2(_19140_),
    .B1(_18395_),
    .C1(_19143_),
    .X(_19144_));
 sky130_vsdinv _25385_ (.A(_19144_),
    .Y(_00416_));
 sky130_fd_sc_hd__buf_1 _25386_ (.A(_18918_),
    .X(_19145_));
 sky130_fd_sc_hd__nor3_4 _25387_ (.A(\timer[0] ),
    .B(\timer[1] ),
    .C(\timer[2] ),
    .Y(_19146_));
 sky130_vsdinv _25388_ (.A(\timer[6] ),
    .Y(_19147_));
 sky130_fd_sc_hd__and4_4 _25389_ (.A(_19146_),
    .B(_19147_),
    .C(_18916_),
    .D(_18911_),
    .X(_19148_));
 sky130_vsdinv _25390_ (.A(\timer[8] ),
    .Y(_19149_));
 sky130_vsdinv _25391_ (.A(\timer[7] ),
    .Y(_19150_));
 sky130_fd_sc_hd__and4_4 _25392_ (.A(_19148_),
    .B(_19149_),
    .C(_19150_),
    .D(_18910_),
    .X(_19151_));
 sky130_fd_sc_hd__buf_1 _25393_ (.A(_19151_),
    .X(_19152_));
 sky130_vsdinv _25394_ (.A(\timer[11] ),
    .Y(_19153_));
 sky130_vsdinv _25395_ (.A(\timer[13] ),
    .Y(_19154_));
 sky130_vsdinv _25396_ (.A(\timer[12] ),
    .Y(_19155_));
 sky130_fd_sc_hd__and4_4 _25397_ (.A(_19152_),
    .B(_19153_),
    .C(_19154_),
    .D(_19155_),
    .X(_19156_));
 sky130_fd_sc_hd__and2_4 _25398_ (.A(_18930_),
    .B(_18922_),
    .X(_19157_));
 sky130_vsdinv _25399_ (.A(\timer[15] ),
    .Y(_19158_));
 sky130_vsdinv _25400_ (.A(\timer[14] ),
    .Y(_19159_));
 sky130_fd_sc_hd__and4_4 _25401_ (.A(_19156_),
    .B(_19157_),
    .C(_19158_),
    .D(_19159_),
    .X(_19160_));
 sky130_fd_sc_hd__buf_1 _25402_ (.A(_19160_),
    .X(_19161_));
 sky130_fd_sc_hd__xor2_4 _25403_ (.A(_19145_),
    .B(_19161_),
    .X(_19162_));
 sky130_fd_sc_hd__buf_1 _25404_ (.A(instr_timer),
    .X(_19163_));
 sky130_fd_sc_hd__nand2_4 _25405_ (.A(_19163_),
    .B(_18797_),
    .Y(_19164_));
 sky130_fd_sc_hd__buf_1 _25406_ (.A(_19164_),
    .X(_19165_));
 sky130_fd_sc_hd__buf_1 _25407_ (.A(_19165_),
    .X(_19166_));
 sky130_vsdinv _25408_ (.A(\decoded_rs2[0] ),
    .Y(_19167_));
 sky130_fd_sc_hd__nand2_4 _25409_ (.A(_19167_),
    .B(\cpu_state[3] ),
    .Y(_19168_));
 sky130_fd_sc_hd__o21a_4 _25410_ (.A1(_18498_),
    .A2(\decoded_rs1[0] ),
    .B1(_19168_),
    .X(_19169_));
 sky130_fd_sc_hd__buf_1 _25411_ (.A(_19169_),
    .X(_19170_));
 sky130_fd_sc_hd__buf_1 _25412_ (.A(_19170_),
    .X(_19171_));
 sky130_fd_sc_hd__buf_1 _25413_ (.A(_19171_),
    .X(_19172_));
 sky130_vsdinv _25414_ (.A(\decoded_rs2[2] ),
    .Y(_19173_));
 sky130_fd_sc_hd__nand2_4 _25415_ (.A(_19173_),
    .B(_18498_),
    .Y(_19174_));
 sky130_fd_sc_hd__o21a_4 _25416_ (.A1(_18499_),
    .A2(\decoded_rs1[2] ),
    .B1(_19174_),
    .X(_19175_));
 sky130_fd_sc_hd__buf_1 _25417_ (.A(_19175_),
    .X(_19176_));
 sky130_fd_sc_hd__nor2_4 _25418_ (.A(_19172_),
    .B(_19176_),
    .Y(_19177_));
 sky130_vsdinv _25419_ (.A(\decoded_rs2[1] ),
    .Y(_19178_));
 sky130_fd_sc_hd__nand2_4 _25420_ (.A(_19178_),
    .B(\cpu_state[3] ),
    .Y(_19179_));
 sky130_fd_sc_hd__o21a_4 _25421_ (.A1(_18498_),
    .A2(\decoded_rs1[1] ),
    .B1(_19179_),
    .X(_19180_));
 sky130_vsdinv _25422_ (.A(_19180_),
    .Y(_19181_));
 sky130_fd_sc_hd__buf_1 _25423_ (.A(_19181_),
    .X(_19182_));
 sky130_fd_sc_hd__buf_1 _25424_ (.A(_19182_),
    .X(_19183_));
 sky130_vsdinv _25425_ (.A(\decoded_rs2[3] ),
    .Y(_19184_));
 sky130_fd_sc_hd__nand2_4 _25426_ (.A(_19184_),
    .B(_18499_),
    .Y(_19185_));
 sky130_fd_sc_hd__o21a_4 _25427_ (.A1(_18499_),
    .A2(\decoded_rs1[3] ),
    .B1(_19185_),
    .X(_19186_));
 sky130_vsdinv _25428_ (.A(_19186_),
    .Y(_19187_));
 sky130_vsdinv _25429_ (.A(\decoded_rs1[4] ),
    .Y(_19188_));
 sky130_fd_sc_hd__nand2_4 _25430_ (.A(_18500_),
    .B(\decoded_rs2[4] ),
    .Y(_19189_));
 sky130_fd_sc_hd__o21a_4 _25431_ (.A1(_18500_),
    .A2(_19188_),
    .B1(_19189_),
    .X(_19190_));
 sky130_fd_sc_hd__and4_4 _25432_ (.A(_19177_),
    .B(_19183_),
    .C(_19187_),
    .D(_19190_),
    .X(_19191_));
 sky130_fd_sc_hd__buf_1 _25433_ (.A(_19191_),
    .X(_19192_));
 sky130_fd_sc_hd__buf_1 _25434_ (.A(_19192_),
    .X(_19193_));
 sky130_fd_sc_hd__buf_1 _25435_ (.A(_19193_),
    .X(_19194_));
 sky130_fd_sc_hd__buf_1 _25436_ (.A(_19170_),
    .X(_19195_));
 sky130_fd_sc_hd__buf_1 _25437_ (.A(_19195_),
    .X(_19196_));
 sky130_fd_sc_hd__buf_1 _25438_ (.A(_19196_),
    .X(_19197_));
 sky130_fd_sc_hd__buf_1 _25439_ (.A(_19197_),
    .X(_19198_));
 sky130_fd_sc_hd__buf_1 _25440_ (.A(_19198_),
    .X(_19199_));
 sky130_fd_sc_hd__buf_1 _25441_ (.A(_19182_),
    .X(_19200_));
 sky130_fd_sc_hd__buf_1 _25442_ (.A(_19200_),
    .X(_19201_));
 sky130_fd_sc_hd__buf_1 _25443_ (.A(_19201_),
    .X(_19202_));
 sky130_fd_sc_hd__buf_1 _25444_ (.A(_19202_),
    .X(_19203_));
 sky130_vsdinv _25445_ (.A(_19170_),
    .Y(_19204_));
 sky130_fd_sc_hd__buf_1 _25446_ (.A(_19204_),
    .X(_19205_));
 sky130_fd_sc_hd__buf_1 _25447_ (.A(_19205_),
    .X(_19206_));
 sky130_fd_sc_hd__buf_1 _25448_ (.A(_19206_),
    .X(_19207_));
 sky130_fd_sc_hd__and2_4 _25449_ (.A(_19207_),
    .B(\cpuregs[18][0] ),
    .X(_19208_));
 sky130_fd_sc_hd__a211o_4 _25450_ (.A1(\cpuregs[19][0] ),
    .A2(_19199_),
    .B1(_19203_),
    .C1(_19208_),
    .X(_19209_));
 sky130_fd_sc_hd__buf_1 _25451_ (.A(_19198_),
    .X(_19210_));
 sky130_fd_sc_hd__buf_1 _25452_ (.A(_19180_),
    .X(_19211_));
 sky130_fd_sc_hd__buf_1 _25453_ (.A(_19211_),
    .X(_19212_));
 sky130_fd_sc_hd__buf_1 _25454_ (.A(_19212_),
    .X(_19213_));
 sky130_fd_sc_hd__buf_1 _25455_ (.A(_19213_),
    .X(_19214_));
 sky130_fd_sc_hd__buf_1 _25456_ (.A(_19214_),
    .X(_19215_));
 sky130_fd_sc_hd__buf_1 _25457_ (.A(_19215_),
    .X(_19216_));
 sky130_fd_sc_hd__buf_1 _25458_ (.A(_19204_),
    .X(_19217_));
 sky130_fd_sc_hd__buf_1 _25459_ (.A(_19217_),
    .X(_19218_));
 sky130_fd_sc_hd__buf_1 _25460_ (.A(_19218_),
    .X(_19219_));
 sky130_fd_sc_hd__and2_4 _25461_ (.A(_19219_),
    .B(\cpuregs[16][0] ),
    .X(_19220_));
 sky130_fd_sc_hd__a211o_4 _25462_ (.A1(\cpuregs[17][0] ),
    .A2(_19210_),
    .B1(_19216_),
    .C1(_19220_),
    .X(_19221_));
 sky130_fd_sc_hd__buf_1 _25463_ (.A(_19190_),
    .X(_19222_));
 sky130_fd_sc_hd__buf_1 _25464_ (.A(_19222_),
    .X(_19223_));
 sky130_fd_sc_hd__buf_1 _25465_ (.A(_19223_),
    .X(_19224_));
 sky130_fd_sc_hd__buf_1 _25466_ (.A(_19224_),
    .X(_19225_));
 sky130_fd_sc_hd__a21oi_4 _25467_ (.A1(_19209_),
    .A2(_19221_),
    .B1(_19225_),
    .Y(_19226_));
 sky130_fd_sc_hd__buf_1 _25468_ (.A(_19206_),
    .X(_19227_));
 sky130_fd_sc_hd__buf_1 _25469_ (.A(_19171_),
    .X(_19228_));
 sky130_fd_sc_hd__buf_1 _25470_ (.A(_19228_),
    .X(_19229_));
 sky130_fd_sc_hd__buf_1 _25471_ (.A(_19182_),
    .X(_19230_));
 sky130_fd_sc_hd__buf_1 _25472_ (.A(_19230_),
    .X(_19231_));
 sky130_fd_sc_hd__o21a_4 _25473_ (.A1(\cpuregs[4][0] ),
    .A2(_19229_),
    .B1(_19231_),
    .X(_19232_));
 sky130_fd_sc_hd__o21ai_4 _25474_ (.A1(\cpuregs[5][0] ),
    .A2(_19227_),
    .B1(_19232_),
    .Y(_19233_));
 sky130_fd_sc_hd__buf_1 _25475_ (.A(_19171_),
    .X(_19234_));
 sky130_fd_sc_hd__buf_1 _25476_ (.A(_19234_),
    .X(_19235_));
 sky130_fd_sc_hd__buf_1 _25477_ (.A(_19212_),
    .X(_19236_));
 sky130_fd_sc_hd__buf_1 _25478_ (.A(_19236_),
    .X(_19237_));
 sky130_fd_sc_hd__o21a_4 _25479_ (.A1(\cpuregs[6][0] ),
    .A2(_19235_),
    .B1(_19237_),
    .X(_19238_));
 sky130_fd_sc_hd__o21ai_4 _25480_ (.A1(\cpuregs[7][0] ),
    .A2(_19227_),
    .B1(_19238_),
    .Y(_19239_));
 sky130_fd_sc_hd__buf_1 _25481_ (.A(_19176_),
    .X(_19240_));
 sky130_fd_sc_hd__buf_1 _25482_ (.A(_19240_),
    .X(_19241_));
 sky130_fd_sc_hd__nand3_4 _25483_ (.A(_19233_),
    .B(_19239_),
    .C(_19241_),
    .Y(_19242_));
 sky130_fd_sc_hd__buf_1 _25484_ (.A(_19200_),
    .X(_19243_));
 sky130_fd_sc_hd__o21a_4 _25485_ (.A1(\cpuregs[0][0] ),
    .A2(_19235_),
    .B1(_19243_),
    .X(_19244_));
 sky130_fd_sc_hd__o21ai_4 _25486_ (.A1(\cpuregs[1][0] ),
    .A2(_19207_),
    .B1(_19244_),
    .Y(_19245_));
 sky130_fd_sc_hd__buf_1 _25487_ (.A(_19234_),
    .X(_19246_));
 sky130_fd_sc_hd__buf_1 _25488_ (.A(_19236_),
    .X(_19247_));
 sky130_fd_sc_hd__o21a_4 _25489_ (.A1(\cpuregs[2][0] ),
    .A2(_19246_),
    .B1(_19247_),
    .X(_19248_));
 sky130_fd_sc_hd__o21ai_4 _25490_ (.A1(\cpuregs[3][0] ),
    .A2(_19219_),
    .B1(_19248_),
    .Y(_19249_));
 sky130_vsdinv _25491_ (.A(_19175_),
    .Y(_19250_));
 sky130_fd_sc_hd__buf_1 _25492_ (.A(_19250_),
    .X(_19251_));
 sky130_fd_sc_hd__buf_1 _25493_ (.A(_19251_),
    .X(_19252_));
 sky130_fd_sc_hd__nand3_4 _25494_ (.A(_19245_),
    .B(_19249_),
    .C(_19252_),
    .Y(_19253_));
 sky130_fd_sc_hd__buf_1 _25495_ (.A(_19187_),
    .X(_19254_));
 sky130_fd_sc_hd__buf_1 _25496_ (.A(_19254_),
    .X(_19255_));
 sky130_fd_sc_hd__nand3_4 _25497_ (.A(_19242_),
    .B(_19253_),
    .C(_19255_),
    .Y(_19256_));
 sky130_fd_sc_hd__buf_1 _25498_ (.A(_19171_),
    .X(_19257_));
 sky130_fd_sc_hd__buf_1 _25499_ (.A(_19257_),
    .X(_19258_));
 sky130_fd_sc_hd__o21a_4 _25500_ (.A1(\cpuregs[12][0] ),
    .A2(_19258_),
    .B1(_19243_),
    .X(_19259_));
 sky130_fd_sc_hd__o21ai_4 _25501_ (.A1(\cpuregs[13][0] ),
    .A2(_19227_),
    .B1(_19259_),
    .Y(_19260_));
 sky130_fd_sc_hd__o21a_4 _25502_ (.A1(\cpuregs[14][0] ),
    .A2(_19246_),
    .B1(_19247_),
    .X(_19261_));
 sky130_fd_sc_hd__o21ai_4 _25503_ (.A1(\cpuregs[15][0] ),
    .A2(_19207_),
    .B1(_19261_),
    .Y(_19262_));
 sky130_fd_sc_hd__buf_1 _25504_ (.A(_19176_),
    .X(_19263_));
 sky130_fd_sc_hd__buf_1 _25505_ (.A(_19263_),
    .X(_19264_));
 sky130_fd_sc_hd__nand3_4 _25506_ (.A(_19260_),
    .B(_19262_),
    .C(_19264_),
    .Y(_19265_));
 sky130_fd_sc_hd__o21a_4 _25507_ (.A1(\cpuregs[8][0] ),
    .A2(_19246_),
    .B1(_19243_),
    .X(_19266_));
 sky130_fd_sc_hd__o21ai_4 _25508_ (.A1(\cpuregs[9][0] ),
    .A2(_19207_),
    .B1(_19266_),
    .Y(_19267_));
 sky130_fd_sc_hd__buf_1 _25509_ (.A(_19195_),
    .X(_19268_));
 sky130_fd_sc_hd__buf_1 _25510_ (.A(_19268_),
    .X(_19269_));
 sky130_fd_sc_hd__buf_1 _25511_ (.A(_19212_),
    .X(_19270_));
 sky130_fd_sc_hd__buf_1 _25512_ (.A(_19270_),
    .X(_19271_));
 sky130_fd_sc_hd__o21a_4 _25513_ (.A1(\cpuregs[10][0] ),
    .A2(_19269_),
    .B1(_19271_),
    .X(_19272_));
 sky130_fd_sc_hd__o21ai_4 _25514_ (.A1(\cpuregs[11][0] ),
    .A2(_19219_),
    .B1(_19272_),
    .Y(_19273_));
 sky130_fd_sc_hd__nand3_4 _25515_ (.A(_19267_),
    .B(_19273_),
    .C(_19252_),
    .Y(_19274_));
 sky130_fd_sc_hd__buf_1 _25516_ (.A(_19186_),
    .X(_19275_));
 sky130_fd_sc_hd__buf_1 _25517_ (.A(_19275_),
    .X(_19276_));
 sky130_fd_sc_hd__nand3_4 _25518_ (.A(_19265_),
    .B(_19274_),
    .C(_19276_),
    .Y(_19277_));
 sky130_fd_sc_hd__buf_1 _25519_ (.A(_19222_),
    .X(_19278_));
 sky130_fd_sc_hd__buf_1 _25520_ (.A(_19278_),
    .X(_19279_));
 sky130_fd_sc_hd__nand3_4 _25521_ (.A(_19256_),
    .B(_19277_),
    .C(_19279_),
    .Y(_19280_));
 sky130_vsdinv _25522_ (.A(_19280_),
    .Y(_19281_));
 sky130_fd_sc_hd__nor3_4 _25523_ (.A(_19194_),
    .B(_19226_),
    .C(_19281_),
    .Y(_19282_));
 sky130_fd_sc_hd__o21ai_4 _25524_ (.A1(_19166_),
    .A2(_19282_),
    .B1(_19126_),
    .Y(_19283_));
 sky130_fd_sc_hd__a21oi_4 _25525_ (.A1(_19162_),
    .A2(_19166_),
    .B1(_19283_),
    .Y(_00626_));
 sky130_fd_sc_hd__buf_1 _25526_ (.A(_19268_),
    .X(_19284_));
 sky130_fd_sc_hd__buf_1 _25527_ (.A(_19181_),
    .X(_19285_));
 sky130_fd_sc_hd__buf_1 _25528_ (.A(_19285_),
    .X(_19286_));
 sky130_fd_sc_hd__buf_1 _25529_ (.A(_19286_),
    .X(_19287_));
 sky130_vsdinv _25530_ (.A(\cpuregs[14][1] ),
    .Y(_19288_));
 sky130_fd_sc_hd__buf_1 _25531_ (.A(_19169_),
    .X(_19289_));
 sky130_fd_sc_hd__buf_1 _25532_ (.A(_19289_),
    .X(_19290_));
 sky130_fd_sc_hd__buf_1 _25533_ (.A(_19290_),
    .X(_19291_));
 sky130_fd_sc_hd__buf_1 _25534_ (.A(_19291_),
    .X(_19292_));
 sky130_fd_sc_hd__nor2_4 _25535_ (.A(_19288_),
    .B(_19292_),
    .Y(_19293_));
 sky130_fd_sc_hd__a211o_4 _25536_ (.A1(\cpuregs[15][1] ),
    .A2(_19284_),
    .B1(_19287_),
    .C1(_19293_),
    .X(_19294_));
 sky130_fd_sc_hd__buf_1 _25537_ (.A(_19289_),
    .X(_19295_));
 sky130_fd_sc_hd__buf_1 _25538_ (.A(_19295_),
    .X(_19296_));
 sky130_fd_sc_hd__buf_1 _25539_ (.A(_19296_),
    .X(_19297_));
 sky130_fd_sc_hd__buf_1 _25540_ (.A(_19211_),
    .X(_19298_));
 sky130_fd_sc_hd__buf_1 _25541_ (.A(_19298_),
    .X(_19299_));
 sky130_vsdinv _25542_ (.A(\cpuregs[12][1] ),
    .Y(_19300_));
 sky130_fd_sc_hd__buf_1 _25543_ (.A(_19295_),
    .X(_19301_));
 sky130_fd_sc_hd__buf_1 _25544_ (.A(_19301_),
    .X(_19302_));
 sky130_fd_sc_hd__nor2_4 _25545_ (.A(_19300_),
    .B(_19302_),
    .Y(_19303_));
 sky130_fd_sc_hd__a211o_4 _25546_ (.A1(\cpuregs[13][1] ),
    .A2(_19297_),
    .B1(_19299_),
    .C1(_19303_),
    .X(_19304_));
 sky130_fd_sc_hd__buf_1 _25547_ (.A(_19250_),
    .X(_19305_));
 sky130_fd_sc_hd__buf_1 _25548_ (.A(_19305_),
    .X(_19306_));
 sky130_fd_sc_hd__a21o_4 _25549_ (.A1(_19294_),
    .A2(_19304_),
    .B1(_19306_),
    .X(_19307_));
 sky130_fd_sc_hd__buf_1 _25550_ (.A(_19289_),
    .X(_19308_));
 sky130_fd_sc_hd__buf_1 _25551_ (.A(_19308_),
    .X(_19309_));
 sky130_fd_sc_hd__buf_1 _25552_ (.A(_19309_),
    .X(_19310_));
 sky130_fd_sc_hd__buf_1 _25553_ (.A(_19211_),
    .X(_19311_));
 sky130_fd_sc_hd__buf_1 _25554_ (.A(_19311_),
    .X(_19312_));
 sky130_vsdinv _25555_ (.A(\cpuregs[8][1] ),
    .Y(_19313_));
 sky130_fd_sc_hd__buf_1 _25556_ (.A(_19170_),
    .X(_19314_));
 sky130_fd_sc_hd__buf_1 _25557_ (.A(_19314_),
    .X(_19315_));
 sky130_fd_sc_hd__nor2_4 _25558_ (.A(_19313_),
    .B(_19315_),
    .Y(_19316_));
 sky130_fd_sc_hd__a211o_4 _25559_ (.A1(\cpuregs[9][1] ),
    .A2(_19310_),
    .B1(_19312_),
    .C1(_19316_),
    .X(_19317_));
 sky130_fd_sc_hd__buf_1 _25560_ (.A(_19290_),
    .X(_19318_));
 sky130_fd_sc_hd__buf_1 _25561_ (.A(_19318_),
    .X(_19319_));
 sky130_fd_sc_hd__buf_1 _25562_ (.A(_19286_),
    .X(_19320_));
 sky130_vsdinv _25563_ (.A(\cpuregs[10][1] ),
    .Y(_19321_));
 sky130_fd_sc_hd__buf_1 _25564_ (.A(_19314_),
    .X(_19322_));
 sky130_fd_sc_hd__nor2_4 _25565_ (.A(_19321_),
    .B(_19322_),
    .Y(_19323_));
 sky130_fd_sc_hd__a211o_4 _25566_ (.A1(\cpuregs[11][1] ),
    .A2(_19319_),
    .B1(_19320_),
    .C1(_19323_),
    .X(_19324_));
 sky130_fd_sc_hd__a21o_4 _25567_ (.A1(_19317_),
    .A2(_19324_),
    .B1(_19240_),
    .X(_19325_));
 sky130_fd_sc_hd__buf_1 _25568_ (.A(_19186_),
    .X(_19326_));
 sky130_fd_sc_hd__buf_1 _25569_ (.A(_19326_),
    .X(_19327_));
 sky130_fd_sc_hd__nand3_4 _25570_ (.A(_19307_),
    .B(_19325_),
    .C(_19327_),
    .Y(_19328_));
 sky130_fd_sc_hd__buf_1 _25571_ (.A(_19222_),
    .X(_19329_));
 sky130_fd_sc_hd__buf_1 _25572_ (.A(_19329_),
    .X(_19330_));
 sky130_fd_sc_hd__and2_4 _25573_ (.A(_19328_),
    .B(_19330_),
    .X(_19331_));
 sky130_fd_sc_hd__buf_1 _25574_ (.A(_19331_),
    .X(_19332_));
 sky130_fd_sc_hd__buf_1 _25575_ (.A(_19290_),
    .X(_19333_));
 sky130_fd_sc_hd__buf_1 _25576_ (.A(_19333_),
    .X(_19334_));
 sky130_fd_sc_hd__buf_1 _25577_ (.A(_19334_),
    .X(_19335_));
 sky130_fd_sc_hd__buf_1 _25578_ (.A(_19312_),
    .X(_19336_));
 sky130_fd_sc_hd__buf_1 _25579_ (.A(_19204_),
    .X(_19337_));
 sky130_fd_sc_hd__buf_1 _25580_ (.A(_19337_),
    .X(_19338_));
 sky130_fd_sc_hd__and2_4 _25581_ (.A(_19338_),
    .B(\cpuregs[0][1] ),
    .X(_19339_));
 sky130_fd_sc_hd__a211o_4 _25582_ (.A1(\cpuregs[1][1] ),
    .A2(_19335_),
    .B1(_19336_),
    .C1(_19339_),
    .X(_19340_));
 sky130_fd_sc_hd__buf_1 _25583_ (.A(_19290_),
    .X(_19341_));
 sky130_fd_sc_hd__buf_1 _25584_ (.A(_19341_),
    .X(_19342_));
 sky130_fd_sc_hd__buf_1 _25585_ (.A(_19342_),
    .X(_19343_));
 sky130_fd_sc_hd__buf_1 _25586_ (.A(_19285_),
    .X(_19344_));
 sky130_fd_sc_hd__buf_1 _25587_ (.A(_19344_),
    .X(_19345_));
 sky130_fd_sc_hd__buf_1 _25588_ (.A(_19345_),
    .X(_19346_));
 sky130_vsdinv _25589_ (.A(\cpuregs[2][1] ),
    .Y(_19347_));
 sky130_fd_sc_hd__buf_1 _25590_ (.A(_19295_),
    .X(_19348_));
 sky130_fd_sc_hd__buf_1 _25591_ (.A(_19348_),
    .X(_19349_));
 sky130_fd_sc_hd__buf_1 _25592_ (.A(_19349_),
    .X(_19350_));
 sky130_fd_sc_hd__nor2_4 _25593_ (.A(_19347_),
    .B(_19350_),
    .Y(_19351_));
 sky130_fd_sc_hd__a211o_4 _25594_ (.A1(\cpuregs[3][1] ),
    .A2(_19343_),
    .B1(_19346_),
    .C1(_19351_),
    .X(_19352_));
 sky130_fd_sc_hd__buf_1 _25595_ (.A(_19175_),
    .X(_19353_));
 sky130_fd_sc_hd__buf_1 _25596_ (.A(_19353_),
    .X(_19354_));
 sky130_fd_sc_hd__buf_1 _25597_ (.A(_19354_),
    .X(_19355_));
 sky130_fd_sc_hd__a21o_4 _25598_ (.A1(_19340_),
    .A2(_19352_),
    .B1(_19355_),
    .X(_19356_));
 sky130_fd_sc_hd__buf_1 _25599_ (.A(_19187_),
    .X(_19357_));
 sky130_fd_sc_hd__buf_1 _25600_ (.A(_19357_),
    .X(_19358_));
 sky130_fd_sc_hd__buf_1 _25601_ (.A(_19333_),
    .X(_19359_));
 sky130_fd_sc_hd__buf_1 _25602_ (.A(_19359_),
    .X(_19360_));
 sky130_fd_sc_hd__buf_1 _25603_ (.A(_19183_),
    .X(_19361_));
 sky130_vsdinv _25604_ (.A(\cpuregs[6][1] ),
    .Y(_19362_));
 sky130_fd_sc_hd__buf_1 _25605_ (.A(_19315_),
    .X(_19363_));
 sky130_fd_sc_hd__nor2_4 _25606_ (.A(_19362_),
    .B(_19363_),
    .Y(_19364_));
 sky130_fd_sc_hd__a211o_4 _25607_ (.A1(\cpuregs[7][1] ),
    .A2(_19360_),
    .B1(_19361_),
    .C1(_19364_),
    .X(_19365_));
 sky130_fd_sc_hd__buf_1 _25608_ (.A(_19289_),
    .X(_19366_));
 sky130_fd_sc_hd__buf_1 _25609_ (.A(_19366_),
    .X(_19367_));
 sky130_fd_sc_hd__buf_1 _25610_ (.A(_19367_),
    .X(_19368_));
 sky130_fd_sc_hd__buf_1 _25611_ (.A(_19368_),
    .X(_19369_));
 sky130_fd_sc_hd__buf_1 _25612_ (.A(_19311_),
    .X(_19370_));
 sky130_fd_sc_hd__buf_1 _25613_ (.A(_19370_),
    .X(_19371_));
 sky130_vsdinv _25614_ (.A(\cpuregs[4][1] ),
    .Y(_19372_));
 sky130_fd_sc_hd__nor2_4 _25615_ (.A(_19372_),
    .B(_19229_),
    .Y(_19373_));
 sky130_fd_sc_hd__a211o_4 _25616_ (.A1(\cpuregs[5][1] ),
    .A2(_19369_),
    .B1(_19371_),
    .C1(_19373_),
    .X(_19374_));
 sky130_fd_sc_hd__buf_1 _25617_ (.A(_19305_),
    .X(_19375_));
 sky130_fd_sc_hd__buf_1 _25618_ (.A(_19375_),
    .X(_19376_));
 sky130_fd_sc_hd__a21o_4 _25619_ (.A1(_19365_),
    .A2(_19374_),
    .B1(_19376_),
    .X(_19377_));
 sky130_fd_sc_hd__nand3_4 _25620_ (.A(_19356_),
    .B(_19358_),
    .C(_19377_),
    .Y(_19378_));
 sky130_fd_sc_hd__buf_1 _25621_ (.A(_19378_),
    .X(_19379_));
 sky130_fd_sc_hd__buf_1 _25622_ (.A(_19165_),
    .X(_19380_));
 sky130_fd_sc_hd__buf_1 _25623_ (.A(_19191_),
    .X(_19381_));
 sky130_fd_sc_hd__buf_1 _25624_ (.A(_19381_),
    .X(_19382_));
 sky130_fd_sc_hd__buf_1 _25625_ (.A(_19382_),
    .X(_19383_));
 sky130_fd_sc_hd__buf_1 _25626_ (.A(_19383_),
    .X(_19384_));
 sky130_fd_sc_hd__buf_1 _25627_ (.A(_19308_),
    .X(_19385_));
 sky130_fd_sc_hd__buf_1 _25628_ (.A(_19385_),
    .X(_19386_));
 sky130_fd_sc_hd__buf_1 _25629_ (.A(_19386_),
    .X(_19387_));
 sky130_fd_sc_hd__buf_1 _25630_ (.A(_19387_),
    .X(_19388_));
 sky130_fd_sc_hd__buf_1 _25631_ (.A(_19344_),
    .X(_19389_));
 sky130_fd_sc_hd__buf_1 _25632_ (.A(_19389_),
    .X(_19390_));
 sky130_fd_sc_hd__buf_1 _25633_ (.A(_19390_),
    .X(_19391_));
 sky130_vsdinv _25634_ (.A(\cpuregs[18][1] ),
    .Y(_19392_));
 sky130_fd_sc_hd__buf_1 _25635_ (.A(_19295_),
    .X(_19393_));
 sky130_fd_sc_hd__buf_1 _25636_ (.A(_19393_),
    .X(_19394_));
 sky130_fd_sc_hd__buf_1 _25637_ (.A(_19394_),
    .X(_19395_));
 sky130_fd_sc_hd__buf_1 _25638_ (.A(_19395_),
    .X(_19396_));
 sky130_fd_sc_hd__nor2_4 _25639_ (.A(_19392_),
    .B(_19396_),
    .Y(_19397_));
 sky130_fd_sc_hd__a211o_4 _25640_ (.A1(\cpuregs[19][1] ),
    .A2(_19388_),
    .B1(_19391_),
    .C1(_19397_),
    .X(_19398_));
 sky130_fd_sc_hd__buf_1 _25641_ (.A(_19314_),
    .X(_19399_));
 sky130_fd_sc_hd__buf_1 _25642_ (.A(_19399_),
    .X(_19400_));
 sky130_fd_sc_hd__buf_1 _25643_ (.A(_19400_),
    .X(_19401_));
 sky130_fd_sc_hd__buf_1 _25644_ (.A(_19371_),
    .X(_19402_));
 sky130_vsdinv _25645_ (.A(\cpuregs[16][1] ),
    .Y(_19403_));
 sky130_fd_sc_hd__buf_1 _25646_ (.A(_19348_),
    .X(_19404_));
 sky130_fd_sc_hd__buf_1 _25647_ (.A(_19404_),
    .X(_19405_));
 sky130_fd_sc_hd__buf_1 _25648_ (.A(_19405_),
    .X(_19406_));
 sky130_fd_sc_hd__nor2_4 _25649_ (.A(_19403_),
    .B(_19406_),
    .Y(_19407_));
 sky130_fd_sc_hd__a211o_4 _25650_ (.A1(\cpuregs[17][1] ),
    .A2(_19401_),
    .B1(_19402_),
    .C1(_19407_),
    .X(_19408_));
 sky130_fd_sc_hd__buf_1 _25651_ (.A(_19222_),
    .X(_19409_));
 sky130_fd_sc_hd__buf_1 _25652_ (.A(_19409_),
    .X(_19410_));
 sky130_fd_sc_hd__a21oi_4 _25653_ (.A1(_19398_),
    .A2(_19408_),
    .B1(_19410_),
    .Y(_19411_));
 sky130_fd_sc_hd__buf_1 _25654_ (.A(_19411_),
    .X(_19412_));
 sky130_fd_sc_hd__a2111o_4 _25655_ (.A1(_19332_),
    .A2(_19379_),
    .B1(_19380_),
    .C1(_19384_),
    .D1(_19412_),
    .X(_19413_));
 sky130_fd_sc_hd__buf_1 _25656_ (.A(_19158_),
    .X(_19414_));
 sky130_fd_sc_hd__buf_1 _25657_ (.A(_19414_),
    .X(_19415_));
 sky130_fd_sc_hd__buf_1 _25658_ (.A(_19156_),
    .X(_19416_));
 sky130_fd_sc_hd__buf_1 _25659_ (.A(_19159_),
    .X(_19417_));
 sky130_vsdinv _25660_ (.A(_19164_),
    .Y(_19418_));
 sky130_fd_sc_hd__a41oi_4 _25661_ (.A1(_19415_),
    .A2(_19416_),
    .A3(_19417_),
    .A4(_19157_),
    .B1(_19418_),
    .Y(_19419_));
 sky130_fd_sc_hd__buf_1 _25662_ (.A(_19419_),
    .X(_19420_));
 sky130_fd_sc_hd__buf_1 _25663_ (.A(_19420_),
    .X(_19421_));
 sky130_fd_sc_hd__buf_1 _25664_ (.A(\timer[1] ),
    .X(_19422_));
 sky130_fd_sc_hd__xnor2_4 _25665_ (.A(_19145_),
    .B(_19422_),
    .Y(_19423_));
 sky130_fd_sc_hd__nand2_4 _25666_ (.A(_19421_),
    .B(_19423_),
    .Y(_19424_));
 sky130_fd_sc_hd__buf_1 _25667_ (.A(_18786_),
    .X(_19425_));
 sky130_fd_sc_hd__buf_1 _25668_ (.A(_19425_),
    .X(_19426_));
 sky130_fd_sc_hd__buf_1 _25669_ (.A(_19426_),
    .X(_19427_));
 sky130_fd_sc_hd__a21oi_4 _25670_ (.A1(_19413_),
    .A2(_19424_),
    .B1(_19427_),
    .Y(_00637_));
 sky130_fd_sc_hd__buf_1 _25671_ (.A(_19366_),
    .X(_19428_));
 sky130_fd_sc_hd__buf_1 _25672_ (.A(_19428_),
    .X(_19429_));
 sky130_fd_sc_hd__buf_1 _25673_ (.A(_19429_),
    .X(_19430_));
 sky130_fd_sc_hd__and2_4 _25674_ (.A(_19205_),
    .B(\cpuregs[12][2] ),
    .X(_19431_));
 sky130_fd_sc_hd__a211o_4 _25675_ (.A1(\cpuregs[13][2] ),
    .A2(_19430_),
    .B1(_19237_),
    .C1(_19431_),
    .X(_19432_));
 sky130_fd_sc_hd__buf_1 _25676_ (.A(_19341_),
    .X(_19433_));
 sky130_fd_sc_hd__buf_1 _25677_ (.A(_19433_),
    .X(_19434_));
 sky130_vsdinv _25678_ (.A(\cpuregs[14][2] ),
    .Y(_19435_));
 sky130_fd_sc_hd__nor2_4 _25679_ (.A(_19435_),
    .B(_19246_),
    .Y(_19436_));
 sky130_fd_sc_hd__a211o_4 _25680_ (.A1(\cpuregs[15][2] ),
    .A2(_19434_),
    .B1(_19231_),
    .C1(_19436_),
    .X(_19437_));
 sky130_fd_sc_hd__buf_1 _25681_ (.A(_19251_),
    .X(_19438_));
 sky130_fd_sc_hd__a21o_4 _25682_ (.A1(_19432_),
    .A2(_19437_),
    .B1(_19438_),
    .X(_19439_));
 sky130_fd_sc_hd__buf_1 _25683_ (.A(_19302_),
    .X(_19440_));
 sky130_fd_sc_hd__and2_4 _25684_ (.A(_19205_),
    .B(\cpuregs[8][2] ),
    .X(_19441_));
 sky130_fd_sc_hd__a211o_4 _25685_ (.A1(\cpuregs[9][2] ),
    .A2(_19440_),
    .B1(_19237_),
    .C1(_19441_),
    .X(_19442_));
 sky130_vsdinv _25686_ (.A(\cpuregs[10][2] ),
    .Y(_19443_));
 sky130_fd_sc_hd__buf_1 _25687_ (.A(_19195_),
    .X(_19444_));
 sky130_fd_sc_hd__buf_1 _25688_ (.A(_19444_),
    .X(_19445_));
 sky130_fd_sc_hd__nor2_4 _25689_ (.A(_19443_),
    .B(_19445_),
    .Y(_19446_));
 sky130_fd_sc_hd__a211o_4 _25690_ (.A1(\cpuregs[11][2] ),
    .A2(_19363_),
    .B1(_19231_),
    .C1(_19446_),
    .X(_19447_));
 sky130_fd_sc_hd__a21o_4 _25691_ (.A1(_19442_),
    .A2(_19447_),
    .B1(_19264_),
    .X(_19448_));
 sky130_fd_sc_hd__nand3_4 _25692_ (.A(_19439_),
    .B(_19448_),
    .C(_19276_),
    .Y(_19449_));
 sky130_fd_sc_hd__and2_4 _25693_ (.A(_19449_),
    .B(_19410_),
    .X(_19450_));
 sky130_fd_sc_hd__buf_1 _25694_ (.A(_19235_),
    .X(_19451_));
 sky130_fd_sc_hd__buf_1 _25695_ (.A(_19214_),
    .X(_19452_));
 sky130_fd_sc_hd__and2_4 _25696_ (.A(_19206_),
    .B(\cpuregs[4][2] ),
    .X(_19453_));
 sky130_fd_sc_hd__a211o_4 _25697_ (.A1(\cpuregs[5][2] ),
    .A2(_19451_),
    .B1(_19452_),
    .C1(_19453_),
    .X(_19454_));
 sky130_fd_sc_hd__buf_1 _25698_ (.A(_19285_),
    .X(_19455_));
 sky130_fd_sc_hd__buf_1 _25699_ (.A(_19455_),
    .X(_19456_));
 sky130_fd_sc_hd__buf_1 _25700_ (.A(_19456_),
    .X(_19457_));
 sky130_vsdinv _25701_ (.A(\cpuregs[6][2] ),
    .Y(_19458_));
 sky130_fd_sc_hd__buf_1 _25702_ (.A(_19269_),
    .X(_19459_));
 sky130_fd_sc_hd__nor2_4 _25703_ (.A(_19458_),
    .B(_19459_),
    .Y(_19460_));
 sky130_fd_sc_hd__a211o_4 _25704_ (.A1(\cpuregs[7][2] ),
    .A2(_19451_),
    .B1(_19457_),
    .C1(_19460_),
    .X(_19461_));
 sky130_fd_sc_hd__buf_1 _25705_ (.A(_19305_),
    .X(_19462_));
 sky130_fd_sc_hd__buf_1 _25706_ (.A(_19462_),
    .X(_19463_));
 sky130_fd_sc_hd__a21o_4 _25707_ (.A1(_19454_),
    .A2(_19461_),
    .B1(_19463_),
    .X(_19464_));
 sky130_fd_sc_hd__and2_4 _25708_ (.A(_19206_),
    .B(\cpuregs[0][2] ),
    .X(_19465_));
 sky130_fd_sc_hd__a211o_4 _25709_ (.A1(\cpuregs[1][2] ),
    .A2(_19451_),
    .B1(_19452_),
    .C1(_19465_),
    .X(_19466_));
 sky130_vsdinv _25710_ (.A(\cpuregs[2][2] ),
    .Y(_19467_));
 sky130_fd_sc_hd__buf_1 _25711_ (.A(_19196_),
    .X(_19468_));
 sky130_fd_sc_hd__buf_1 _25712_ (.A(_19468_),
    .X(_19469_));
 sky130_fd_sc_hd__nor2_4 _25713_ (.A(_19467_),
    .B(_19469_),
    .Y(_19470_));
 sky130_fd_sc_hd__a211o_4 _25714_ (.A1(\cpuregs[3][2] ),
    .A2(_19451_),
    .B1(_19457_),
    .C1(_19470_),
    .X(_19471_));
 sky130_fd_sc_hd__buf_1 _25715_ (.A(_19176_),
    .X(_19472_));
 sky130_fd_sc_hd__buf_1 _25716_ (.A(_19472_),
    .X(_19473_));
 sky130_fd_sc_hd__buf_1 _25717_ (.A(_19473_),
    .X(_19474_));
 sky130_fd_sc_hd__a21o_4 _25718_ (.A1(_19466_),
    .A2(_19471_),
    .B1(_19474_),
    .X(_19475_));
 sky130_fd_sc_hd__buf_1 _25719_ (.A(_19254_),
    .X(_19476_));
 sky130_fd_sc_hd__buf_1 _25720_ (.A(_19476_),
    .X(_19477_));
 sky130_fd_sc_hd__nand3_4 _25721_ (.A(_19464_),
    .B(_19475_),
    .C(_19477_),
    .Y(_19478_));
 sky130_fd_sc_hd__buf_1 _25722_ (.A(_19165_),
    .X(_19479_));
 sky130_fd_sc_hd__buf_1 _25723_ (.A(_19195_),
    .X(_19480_));
 sky130_fd_sc_hd__buf_1 _25724_ (.A(_19480_),
    .X(_19481_));
 sky130_fd_sc_hd__buf_1 _25725_ (.A(_19481_),
    .X(_19482_));
 sky130_fd_sc_hd__buf_1 _25726_ (.A(_19482_),
    .X(_19483_));
 sky130_fd_sc_hd__and2_4 _25727_ (.A(_19227_),
    .B(\cpuregs[16][2] ),
    .X(_19484_));
 sky130_fd_sc_hd__a211o_4 _25728_ (.A1(\cpuregs[17][2] ),
    .A2(_19483_),
    .B1(_19216_),
    .C1(_19484_),
    .X(_19485_));
 sky130_vsdinv _25729_ (.A(\cpuregs[18][2] ),
    .Y(_19486_));
 sky130_fd_sc_hd__nor2_4 _25730_ (.A(_19486_),
    .B(_19483_),
    .Y(_19487_));
 sky130_fd_sc_hd__a211o_4 _25731_ (.A1(\cpuregs[19][2] ),
    .A2(_19483_),
    .B1(_19203_),
    .C1(_19487_),
    .X(_19488_));
 sky130_fd_sc_hd__a21oi_4 _25732_ (.A1(_19485_),
    .A2(_19488_),
    .B1(_19225_),
    .Y(_19489_));
 sky130_fd_sc_hd__a2111o_4 _25733_ (.A1(_19450_),
    .A2(_19478_),
    .B1(_19479_),
    .C1(_19384_),
    .D1(_19489_),
    .X(_19490_));
 sky130_fd_sc_hd__o21a_4 _25734_ (.A1(_19145_),
    .A2(_19422_),
    .B1(\timer[2] ),
    .X(_19491_));
 sky130_fd_sc_hd__buf_1 _25735_ (.A(_19420_),
    .X(_19492_));
 sky130_fd_sc_hd__o21ai_4 _25736_ (.A1(_19146_),
    .A2(_19491_),
    .B1(_19492_),
    .Y(_19493_));
 sky130_fd_sc_hd__buf_1 _25737_ (.A(_18786_),
    .X(_19494_));
 sky130_fd_sc_hd__buf_1 _25738_ (.A(_19494_),
    .X(_19495_));
 sky130_fd_sc_hd__buf_1 _25739_ (.A(_19495_),
    .X(_19496_));
 sky130_fd_sc_hd__a21oi_4 _25740_ (.A1(_19490_),
    .A2(_19493_),
    .B1(_19496_),
    .Y(_00648_));
 sky130_fd_sc_hd__buf_1 _25741_ (.A(_19309_),
    .X(_19497_));
 sky130_fd_sc_hd__buf_1 _25742_ (.A(_19204_),
    .X(_19498_));
 sky130_fd_sc_hd__and2_4 _25743_ (.A(_19498_),
    .B(\cpuregs[12][3] ),
    .X(_19499_));
 sky130_fd_sc_hd__a211o_4 _25744_ (.A1(\cpuregs[13][3] ),
    .A2(_19497_),
    .B1(_19214_),
    .C1(_19499_),
    .X(_19500_));
 sky130_fd_sc_hd__buf_1 _25745_ (.A(_19367_),
    .X(_19501_));
 sky130_vsdinv _25746_ (.A(\cpuregs[14][3] ),
    .Y(_19502_));
 sky130_fd_sc_hd__buf_1 _25747_ (.A(_19341_),
    .X(_19503_));
 sky130_fd_sc_hd__nor2_4 _25748_ (.A(_19502_),
    .B(_19503_),
    .Y(_19504_));
 sky130_fd_sc_hd__a211o_4 _25749_ (.A1(\cpuregs[15][3] ),
    .A2(_19501_),
    .B1(_19287_),
    .C1(_19504_),
    .X(_19505_));
 sky130_fd_sc_hd__a21o_4 _25750_ (.A1(_19500_),
    .A2(_19505_),
    .B1(_19462_),
    .X(_19506_));
 sky130_fd_sc_hd__buf_1 _25751_ (.A(_19385_),
    .X(_19507_));
 sky130_fd_sc_hd__buf_1 _25752_ (.A(_19298_),
    .X(_19508_));
 sky130_fd_sc_hd__and2_4 _25753_ (.A(_19498_),
    .B(\cpuregs[8][3] ),
    .X(_19509_));
 sky130_fd_sc_hd__a211o_4 _25754_ (.A1(\cpuregs[9][3] ),
    .A2(_19507_),
    .B1(_19508_),
    .C1(_19509_),
    .X(_19510_));
 sky130_fd_sc_hd__buf_1 _25755_ (.A(_19366_),
    .X(_19511_));
 sky130_fd_sc_hd__buf_1 _25756_ (.A(_19511_),
    .X(_19512_));
 sky130_fd_sc_hd__buf_1 _25757_ (.A(_19344_),
    .X(_19513_));
 sky130_vsdinv _25758_ (.A(\cpuregs[10][3] ),
    .Y(_19514_));
 sky130_fd_sc_hd__buf_1 _25759_ (.A(_19393_),
    .X(_19515_));
 sky130_fd_sc_hd__nor2_4 _25760_ (.A(_19514_),
    .B(_19515_),
    .Y(_19516_));
 sky130_fd_sc_hd__a211o_4 _25761_ (.A1(\cpuregs[11][3] ),
    .A2(_19512_),
    .B1(_19513_),
    .C1(_19516_),
    .X(_19517_));
 sky130_fd_sc_hd__buf_1 _25762_ (.A(_19353_),
    .X(_19518_));
 sky130_fd_sc_hd__a21o_4 _25763_ (.A1(_19510_),
    .A2(_19517_),
    .B1(_19518_),
    .X(_19519_));
 sky130_fd_sc_hd__buf_1 _25764_ (.A(_19326_),
    .X(_19520_));
 sky130_fd_sc_hd__nand3_4 _25765_ (.A(_19506_),
    .B(_19519_),
    .C(_19520_),
    .Y(_19521_));
 sky130_fd_sc_hd__buf_1 _25766_ (.A(_19329_),
    .X(_19522_));
 sky130_fd_sc_hd__and2_4 _25767_ (.A(_19521_),
    .B(_19522_),
    .X(_19523_));
 sky130_fd_sc_hd__buf_1 _25768_ (.A(_19366_),
    .X(_19524_));
 sky130_fd_sc_hd__buf_1 _25769_ (.A(_19524_),
    .X(_19525_));
 sky130_fd_sc_hd__buf_1 _25770_ (.A(_19525_),
    .X(_19526_));
 sky130_fd_sc_hd__buf_1 _25771_ (.A(_19370_),
    .X(_19527_));
 sky130_fd_sc_hd__buf_1 _25772_ (.A(_19217_),
    .X(_19528_));
 sky130_fd_sc_hd__and2_4 _25773_ (.A(_19528_),
    .B(\cpuregs[4][3] ),
    .X(_19529_));
 sky130_fd_sc_hd__a211o_4 _25774_ (.A1(\cpuregs[5][3] ),
    .A2(_19526_),
    .B1(_19527_),
    .C1(_19529_),
    .X(_19530_));
 sky130_fd_sc_hd__buf_1 _25775_ (.A(_19348_),
    .X(_19531_));
 sky130_fd_sc_hd__buf_1 _25776_ (.A(_19531_),
    .X(_19532_));
 sky130_fd_sc_hd__buf_1 _25777_ (.A(_19182_),
    .X(_19533_));
 sky130_fd_sc_hd__buf_1 _25778_ (.A(_19533_),
    .X(_19534_));
 sky130_vsdinv _25779_ (.A(\cpuregs[6][3] ),
    .Y(_19535_));
 sky130_fd_sc_hd__buf_1 _25780_ (.A(_19515_),
    .X(_19536_));
 sky130_fd_sc_hd__nor2_4 _25781_ (.A(_19535_),
    .B(_19536_),
    .Y(_19537_));
 sky130_fd_sc_hd__a211o_4 _25782_ (.A1(\cpuregs[7][3] ),
    .A2(_19532_),
    .B1(_19534_),
    .C1(_19537_),
    .X(_19538_));
 sky130_fd_sc_hd__buf_1 _25783_ (.A(_19375_),
    .X(_19539_));
 sky130_fd_sc_hd__a21o_4 _25784_ (.A1(_19530_),
    .A2(_19538_),
    .B1(_19539_),
    .X(_19540_));
 sky130_fd_sc_hd__buf_1 _25785_ (.A(_19212_),
    .X(_19541_));
 sky130_fd_sc_hd__buf_1 _25786_ (.A(_19541_),
    .X(_19542_));
 sky130_fd_sc_hd__and2_4 _25787_ (.A(_19218_),
    .B(\cpuregs[0][3] ),
    .X(_19543_));
 sky130_fd_sc_hd__a211o_4 _25788_ (.A1(\cpuregs[1][3] ),
    .A2(_19387_),
    .B1(_19542_),
    .C1(_19543_),
    .X(_19544_));
 sky130_fd_sc_hd__buf_1 _25789_ (.A(_19525_),
    .X(_19545_));
 sky130_vsdinv _25790_ (.A(\cpuregs[2][3] ),
    .Y(_19546_));
 sky130_fd_sc_hd__buf_1 _25791_ (.A(_19322_),
    .X(_19547_));
 sky130_fd_sc_hd__nor2_4 _25792_ (.A(_19546_),
    .B(_19547_),
    .Y(_19548_));
 sky130_fd_sc_hd__a211o_4 _25793_ (.A1(\cpuregs[3][3] ),
    .A2(_19545_),
    .B1(_19390_),
    .C1(_19548_),
    .X(_19549_));
 sky130_fd_sc_hd__a21o_4 _25794_ (.A1(_19544_),
    .A2(_19549_),
    .B1(_19241_),
    .X(_19550_));
 sky130_fd_sc_hd__nand3_4 _25795_ (.A(_19540_),
    .B(_19550_),
    .C(_19358_),
    .Y(_19551_));
 sky130_fd_sc_hd__buf_1 _25796_ (.A(_19383_),
    .X(_19552_));
 sky130_fd_sc_hd__and2_4 _25797_ (.A(_19219_),
    .B(\cpuregs[16][3] ),
    .X(_19553_));
 sky130_fd_sc_hd__a211o_4 _25798_ (.A1(\cpuregs[17][3] ),
    .A2(_19401_),
    .B1(_19402_),
    .C1(_19553_),
    .X(_19554_));
 sky130_fd_sc_hd__buf_1 _25799_ (.A(_19308_),
    .X(_19555_));
 sky130_fd_sc_hd__buf_1 _25800_ (.A(_19555_),
    .X(_19556_));
 sky130_fd_sc_hd__buf_1 _25801_ (.A(_19556_),
    .X(_19557_));
 sky130_fd_sc_hd__buf_1 _25802_ (.A(_19557_),
    .X(_19558_));
 sky130_vsdinv _25803_ (.A(\cpuregs[18][3] ),
    .Y(_19559_));
 sky130_fd_sc_hd__nor2_4 _25804_ (.A(_19559_),
    .B(_19406_),
    .Y(_19560_));
 sky130_fd_sc_hd__a211o_4 _25805_ (.A1(\cpuregs[19][3] ),
    .A2(_19558_),
    .B1(_19391_),
    .C1(_19560_),
    .X(_19561_));
 sky130_fd_sc_hd__a21oi_4 _25806_ (.A1(_19554_),
    .A2(_19561_),
    .B1(_19279_),
    .Y(_19562_));
 sky130_fd_sc_hd__a2111o_4 _25807_ (.A1(_19523_),
    .A2(_19551_),
    .B1(_19479_),
    .C1(_19552_),
    .D1(_19562_),
    .X(_19563_));
 sky130_vsdinv _25808_ (.A(_18918_),
    .Y(_19564_));
 sky130_fd_sc_hd__nand4_4 _25809_ (.A(_19564_),
    .B(_18914_),
    .C(_18915_),
    .D(_18916_),
    .Y(_19565_));
 sky130_vsdinv _25810_ (.A(_19565_),
    .Y(_19566_));
 sky130_fd_sc_hd__nor2_4 _25811_ (.A(_18918_),
    .B(_19422_),
    .Y(_19567_));
 sky130_fd_sc_hd__a21oi_4 _25812_ (.A1(_19567_),
    .A2(_18915_),
    .B1(_18917_),
    .Y(_19568_));
 sky130_fd_sc_hd__o21ai_4 _25813_ (.A1(_19566_),
    .A2(_19568_),
    .B1(_19492_),
    .Y(_19569_));
 sky130_fd_sc_hd__a21oi_4 _25814_ (.A1(_19563_),
    .A2(_19569_),
    .B1(_19496_),
    .Y(_00651_));
 sky130_fd_sc_hd__buf_1 _25815_ (.A(_19285_),
    .X(_19570_));
 sky130_fd_sc_hd__buf_1 _25816_ (.A(_19570_),
    .X(_19571_));
 sky130_vsdinv _25817_ (.A(\cpuregs[14][4] ),
    .Y(_19572_));
 sky130_fd_sc_hd__buf_1 _25818_ (.A(_19308_),
    .X(_19573_));
 sky130_fd_sc_hd__buf_1 _25819_ (.A(_19573_),
    .X(_19574_));
 sky130_fd_sc_hd__nor2_4 _25820_ (.A(_19572_),
    .B(_19574_),
    .Y(_19575_));
 sky130_fd_sc_hd__a211o_4 _25821_ (.A1(\cpuregs[15][4] ),
    .A2(_19468_),
    .B1(_19571_),
    .C1(_19575_),
    .X(_19576_));
 sky130_fd_sc_hd__buf_1 _25822_ (.A(_19524_),
    .X(_19577_));
 sky130_fd_sc_hd__buf_1 _25823_ (.A(_19213_),
    .X(_19578_));
 sky130_vsdinv _25824_ (.A(\cpuregs[12][4] ),
    .Y(_19579_));
 sky130_fd_sc_hd__buf_1 _25825_ (.A(_19428_),
    .X(_19580_));
 sky130_fd_sc_hd__nor2_4 _25826_ (.A(_19579_),
    .B(_19580_),
    .Y(_19581_));
 sky130_fd_sc_hd__a211o_4 _25827_ (.A1(\cpuregs[13][4] ),
    .A2(_19577_),
    .B1(_19578_),
    .C1(_19581_),
    .X(_19582_));
 sky130_fd_sc_hd__buf_1 _25828_ (.A(_19250_),
    .X(_19583_));
 sky130_fd_sc_hd__buf_1 _25829_ (.A(_19583_),
    .X(_19584_));
 sky130_fd_sc_hd__a21o_4 _25830_ (.A1(_19576_),
    .A2(_19582_),
    .B1(_19584_),
    .X(_19585_));
 sky130_fd_sc_hd__buf_1 _25831_ (.A(_19367_),
    .X(_19586_));
 sky130_fd_sc_hd__buf_1 _25832_ (.A(_19211_),
    .X(_19587_));
 sky130_fd_sc_hd__buf_1 _25833_ (.A(_19587_),
    .X(_19588_));
 sky130_vsdinv _25834_ (.A(\cpuregs[8][4] ),
    .Y(_19589_));
 sky130_fd_sc_hd__buf_1 _25835_ (.A(_19291_),
    .X(_19590_));
 sky130_fd_sc_hd__nor2_4 _25836_ (.A(_19589_),
    .B(_19590_),
    .Y(_19591_));
 sky130_fd_sc_hd__a211o_4 _25837_ (.A1(\cpuregs[9][4] ),
    .A2(_19586_),
    .B1(_19588_),
    .C1(_19591_),
    .X(_19592_));
 sky130_fd_sc_hd__buf_1 _25838_ (.A(_19385_),
    .X(_19593_));
 sky130_fd_sc_hd__buf_1 _25839_ (.A(_19455_),
    .X(_19594_));
 sky130_vsdinv _25840_ (.A(\cpuregs[10][4] ),
    .Y(_19595_));
 sky130_fd_sc_hd__buf_1 _25841_ (.A(_19301_),
    .X(_19596_));
 sky130_fd_sc_hd__nor2_4 _25842_ (.A(_19595_),
    .B(_19596_),
    .Y(_19597_));
 sky130_fd_sc_hd__a211o_4 _25843_ (.A1(\cpuregs[11][4] ),
    .A2(_19593_),
    .B1(_19594_),
    .C1(_19597_),
    .X(_19598_));
 sky130_fd_sc_hd__buf_1 _25844_ (.A(_19472_),
    .X(_19599_));
 sky130_fd_sc_hd__a21o_4 _25845_ (.A1(_19592_),
    .A2(_19598_),
    .B1(_19599_),
    .X(_19600_));
 sky130_fd_sc_hd__buf_1 _25846_ (.A(_19275_),
    .X(_19601_));
 sky130_fd_sc_hd__nand3_4 _25847_ (.A(_19585_),
    .B(_19600_),
    .C(_19601_),
    .Y(_19602_));
 sky130_fd_sc_hd__buf_1 _25848_ (.A(_19329_),
    .X(_19603_));
 sky130_fd_sc_hd__and2_4 _25849_ (.A(_19602_),
    .B(_19603_),
    .X(_19604_));
 sky130_fd_sc_hd__buf_1 _25850_ (.A(_19334_),
    .X(_19605_));
 sky130_fd_sc_hd__buf_1 _25851_ (.A(_19370_),
    .X(_19606_));
 sky130_fd_sc_hd__and2_4 _25852_ (.A(_19338_),
    .B(\cpuregs[0][4] ),
    .X(_19607_));
 sky130_fd_sc_hd__a211o_4 _25853_ (.A1(\cpuregs[1][4] ),
    .A2(_19605_),
    .B1(_19606_),
    .C1(_19607_),
    .X(_19608_));
 sky130_fd_sc_hd__buf_1 _25854_ (.A(_19385_),
    .X(_19609_));
 sky130_fd_sc_hd__buf_1 _25855_ (.A(_19609_),
    .X(_19610_));
 sky130_vsdinv _25856_ (.A(\cpuregs[2][4] ),
    .Y(_19611_));
 sky130_fd_sc_hd__buf_1 _25857_ (.A(_19349_),
    .X(_19612_));
 sky130_fd_sc_hd__nor2_4 _25858_ (.A(_19611_),
    .B(_19612_),
    .Y(_19613_));
 sky130_fd_sc_hd__a211o_4 _25859_ (.A1(\cpuregs[3][4] ),
    .A2(_19610_),
    .B1(_19346_),
    .C1(_19613_),
    .X(_19614_));
 sky130_fd_sc_hd__a21o_4 _25860_ (.A1(_19608_),
    .A2(_19614_),
    .B1(_19355_),
    .X(_19615_));
 sky130_fd_sc_hd__buf_1 _25861_ (.A(_19357_),
    .X(_19616_));
 sky130_vsdinv _25862_ (.A(\cpuregs[6][4] ),
    .Y(_19617_));
 sky130_fd_sc_hd__nor2_4 _25863_ (.A(_19617_),
    .B(_19536_),
    .Y(_19618_));
 sky130_fd_sc_hd__a211o_4 _25864_ (.A1(\cpuregs[7][4] ),
    .A2(_19532_),
    .B1(_19534_),
    .C1(_19618_),
    .X(_19619_));
 sky130_fd_sc_hd__buf_1 _25865_ (.A(_19394_),
    .X(_19620_));
 sky130_fd_sc_hd__buf_1 _25866_ (.A(_19541_),
    .X(_19621_));
 sky130_vsdinv _25867_ (.A(\cpuregs[4][4] ),
    .Y(_19622_));
 sky130_fd_sc_hd__buf_1 _25868_ (.A(_19314_),
    .X(_19623_));
 sky130_fd_sc_hd__buf_1 _25869_ (.A(_19623_),
    .X(_19624_));
 sky130_fd_sc_hd__nor2_4 _25870_ (.A(_19622_),
    .B(_19624_),
    .Y(_19625_));
 sky130_fd_sc_hd__a211o_4 _25871_ (.A1(\cpuregs[5][4] ),
    .A2(_19620_),
    .B1(_19621_),
    .C1(_19625_),
    .X(_19626_));
 sky130_fd_sc_hd__buf_1 _25872_ (.A(_19375_),
    .X(_19627_));
 sky130_fd_sc_hd__a21o_4 _25873_ (.A1(_19619_),
    .A2(_19626_),
    .B1(_19627_),
    .X(_19628_));
 sky130_fd_sc_hd__nand3_4 _25874_ (.A(_19615_),
    .B(_19616_),
    .C(_19628_),
    .Y(_19629_));
 sky130_fd_sc_hd__buf_1 _25875_ (.A(_19480_),
    .X(_19630_));
 sky130_fd_sc_hd__buf_1 _25876_ (.A(_19630_),
    .X(_19631_));
 sky130_fd_sc_hd__buf_1 _25877_ (.A(_19631_),
    .X(_19632_));
 sky130_fd_sc_hd__buf_1 _25878_ (.A(_19389_),
    .X(_19633_));
 sky130_fd_sc_hd__buf_1 _25879_ (.A(_19633_),
    .X(_19634_));
 sky130_vsdinv _25880_ (.A(\cpuregs[18][4] ),
    .Y(_19635_));
 sky130_fd_sc_hd__buf_1 _25881_ (.A(_19369_),
    .X(_19636_));
 sky130_fd_sc_hd__nor2_4 _25882_ (.A(_19635_),
    .B(_19636_),
    .Y(_19637_));
 sky130_fd_sc_hd__a211o_4 _25883_ (.A1(\cpuregs[19][4] ),
    .A2(_19632_),
    .B1(_19634_),
    .C1(_19637_),
    .X(_19638_));
 sky130_fd_sc_hd__buf_1 _25884_ (.A(_19334_),
    .X(_19639_));
 sky130_fd_sc_hd__buf_1 _25885_ (.A(_19639_),
    .X(_19640_));
 sky130_fd_sc_hd__buf_1 _25886_ (.A(_19527_),
    .X(_19641_));
 sky130_vsdinv _25887_ (.A(\cpuregs[16][4] ),
    .Y(_19642_));
 sky130_fd_sc_hd__buf_1 _25888_ (.A(_19386_),
    .X(_19643_));
 sky130_fd_sc_hd__buf_1 _25889_ (.A(_19643_),
    .X(_19644_));
 sky130_fd_sc_hd__nor2_4 _25890_ (.A(_19642_),
    .B(_19644_),
    .Y(_19645_));
 sky130_fd_sc_hd__a211o_4 _25891_ (.A1(\cpuregs[17][4] ),
    .A2(_19640_),
    .B1(_19641_),
    .C1(_19645_),
    .X(_19646_));
 sky130_fd_sc_hd__buf_1 _25892_ (.A(_19224_),
    .X(_19647_));
 sky130_fd_sc_hd__a21oi_4 _25893_ (.A1(_19638_),
    .A2(_19646_),
    .B1(_19647_),
    .Y(_19648_));
 sky130_fd_sc_hd__a2111o_4 _25894_ (.A1(_19604_),
    .A2(_19629_),
    .B1(_19479_),
    .C1(_19552_),
    .D1(_19648_),
    .X(_19649_));
 sky130_vsdinv _25895_ (.A(\timer[4] ),
    .Y(_19650_));
 sky130_fd_sc_hd__xor2_4 _25896_ (.A(_19650_),
    .B(_19565_),
    .X(_19651_));
 sky130_fd_sc_hd__nand2_4 _25897_ (.A(_19421_),
    .B(_19651_),
    .Y(_19652_));
 sky130_fd_sc_hd__a21oi_4 _25898_ (.A1(_19649_),
    .A2(_19652_),
    .B1(_19496_),
    .Y(_00652_));
 sky130_fd_sc_hd__buf_1 _25899_ (.A(_19196_),
    .X(_19653_));
 sky130_vsdinv _25900_ (.A(\cpuregs[14][5] ),
    .Y(_19654_));
 sky130_fd_sc_hd__buf_1 _25901_ (.A(_19296_),
    .X(_19655_));
 sky130_fd_sc_hd__nor2_4 _25902_ (.A(_19654_),
    .B(_19655_),
    .Y(_19656_));
 sky130_fd_sc_hd__a211o_4 _25903_ (.A1(\cpuregs[15][5] ),
    .A2(_19653_),
    .B1(_19571_),
    .C1(_19656_),
    .X(_19657_));
 sky130_vsdinv _25904_ (.A(\cpuregs[12][5] ),
    .Y(_19658_));
 sky130_fd_sc_hd__buf_1 _25905_ (.A(_19428_),
    .X(_19659_));
 sky130_fd_sc_hd__nor2_4 _25906_ (.A(_19658_),
    .B(_19659_),
    .Y(_19660_));
 sky130_fd_sc_hd__a211o_4 _25907_ (.A1(\cpuregs[13][5] ),
    .A2(_19577_),
    .B1(_19578_),
    .C1(_19660_),
    .X(_19661_));
 sky130_fd_sc_hd__a21o_4 _25908_ (.A1(_19657_),
    .A2(_19661_),
    .B1(_19584_),
    .X(_19662_));
 sky130_vsdinv _25909_ (.A(\cpuregs[8][5] ),
    .Y(_19663_));
 sky130_fd_sc_hd__nor2_4 _25910_ (.A(_19663_),
    .B(_19590_),
    .Y(_19664_));
 sky130_fd_sc_hd__a211o_4 _25911_ (.A1(\cpuregs[9][5] ),
    .A2(_19586_),
    .B1(_19588_),
    .C1(_19664_),
    .X(_19665_));
 sky130_vsdinv _25912_ (.A(\cpuregs[10][5] ),
    .Y(_19666_));
 sky130_fd_sc_hd__nor2_4 _25913_ (.A(_19666_),
    .B(_19596_),
    .Y(_19667_));
 sky130_fd_sc_hd__a211o_4 _25914_ (.A1(\cpuregs[11][5] ),
    .A2(_19197_),
    .B1(_19594_),
    .C1(_19667_),
    .X(_19668_));
 sky130_fd_sc_hd__a21o_4 _25915_ (.A1(_19665_),
    .A2(_19668_),
    .B1(_19599_),
    .X(_19669_));
 sky130_fd_sc_hd__nand3_4 _25916_ (.A(_19662_),
    .B(_19669_),
    .C(_19601_),
    .Y(_19670_));
 sky130_fd_sc_hd__and2_4 _25917_ (.A(_19670_),
    .B(_19603_),
    .X(_19671_));
 sky130_fd_sc_hd__and2_4 _25918_ (.A(_19338_),
    .B(\cpuregs[0][5] ),
    .X(_19672_));
 sky130_fd_sc_hd__a211o_4 _25919_ (.A1(\cpuregs[1][5] ),
    .A2(_19605_),
    .B1(_19606_),
    .C1(_19672_),
    .X(_19673_));
 sky130_vsdinv _25920_ (.A(\cpuregs[2][5] ),
    .Y(_19674_));
 sky130_fd_sc_hd__nor2_4 _25921_ (.A(_19674_),
    .B(_19612_),
    .Y(_19675_));
 sky130_fd_sc_hd__a211o_4 _25922_ (.A1(\cpuregs[3][5] ),
    .A2(_19610_),
    .B1(_19346_),
    .C1(_19675_),
    .X(_19676_));
 sky130_fd_sc_hd__buf_1 _25923_ (.A(_19518_),
    .X(_19677_));
 sky130_fd_sc_hd__a21o_4 _25924_ (.A1(_19673_),
    .A2(_19676_),
    .B1(_19677_),
    .X(_19678_));
 sky130_vsdinv _25925_ (.A(\cpuregs[6][5] ),
    .Y(_19679_));
 sky130_fd_sc_hd__nor2_4 _25926_ (.A(_19679_),
    .B(_19536_),
    .Y(_19680_));
 sky130_fd_sc_hd__a211o_4 _25927_ (.A1(\cpuregs[7][5] ),
    .A2(_19557_),
    .B1(_19534_),
    .C1(_19680_),
    .X(_19681_));
 sky130_vsdinv _25928_ (.A(\cpuregs[4][5] ),
    .Y(_19682_));
 sky130_fd_sc_hd__nor2_4 _25929_ (.A(_19682_),
    .B(_19624_),
    .Y(_19683_));
 sky130_fd_sc_hd__a211o_4 _25930_ (.A1(\cpuregs[5][5] ),
    .A2(_19620_),
    .B1(_19621_),
    .C1(_19683_),
    .X(_19684_));
 sky130_fd_sc_hd__a21o_4 _25931_ (.A1(_19681_),
    .A2(_19684_),
    .B1(_19376_),
    .X(_19685_));
 sky130_fd_sc_hd__nand3_4 _25932_ (.A(_19678_),
    .B(_19616_),
    .C(_19685_),
    .Y(_19686_));
 sky130_vsdinv _25933_ (.A(\cpuregs[18][5] ),
    .Y(_19687_));
 sky130_fd_sc_hd__nor2_4 _25934_ (.A(_19687_),
    .B(_19636_),
    .Y(_19688_));
 sky130_fd_sc_hd__a211o_4 _25935_ (.A1(\cpuregs[19][5] ),
    .A2(_19632_),
    .B1(_19634_),
    .C1(_19688_),
    .X(_19689_));
 sky130_vsdinv _25936_ (.A(\cpuregs[16][5] ),
    .Y(_19690_));
 sky130_fd_sc_hd__nor2_4 _25937_ (.A(_19690_),
    .B(_19644_),
    .Y(_19691_));
 sky130_fd_sc_hd__a211o_4 _25938_ (.A1(\cpuregs[17][5] ),
    .A2(_19640_),
    .B1(_19641_),
    .C1(_19691_),
    .X(_19692_));
 sky130_fd_sc_hd__a21oi_4 _25939_ (.A1(_19689_),
    .A2(_19692_),
    .B1(_19647_),
    .Y(_19693_));
 sky130_fd_sc_hd__a2111o_4 _25940_ (.A1(_19671_),
    .A2(_19686_),
    .B1(_19479_),
    .C1(_19552_),
    .D1(_19693_),
    .X(_19694_));
 sky130_fd_sc_hd__and4_4 _25941_ (.A(_18911_),
    .B(_19567_),
    .C(_18915_),
    .D(_18917_),
    .X(_19695_));
 sky130_fd_sc_hd__buf_1 _25942_ (.A(_19695_),
    .X(_19696_));
 sky130_fd_sc_hd__o21a_4 _25943_ (.A1(\timer[4] ),
    .A2(_19565_),
    .B1(\timer[5] ),
    .X(_19697_));
 sky130_fd_sc_hd__o21ai_4 _25944_ (.A1(_19696_),
    .A2(_19697_),
    .B1(_19492_),
    .Y(_19698_));
 sky130_fd_sc_hd__a21oi_4 _25945_ (.A1(_19694_),
    .A2(_19698_),
    .B1(_19496_),
    .Y(_00653_));
 sky130_vsdinv _25946_ (.A(\cpuregs[14][6] ),
    .Y(_19699_));
 sky130_fd_sc_hd__nor2_4 _25947_ (.A(_19699_),
    .B(_19655_),
    .Y(_19700_));
 sky130_fd_sc_hd__a211o_4 _25948_ (.A1(\cpuregs[15][6] ),
    .A2(_19653_),
    .B1(_19571_),
    .C1(_19700_),
    .X(_19701_));
 sky130_fd_sc_hd__buf_1 _25949_ (.A(_19213_),
    .X(_19702_));
 sky130_vsdinv _25950_ (.A(\cpuregs[12][6] ),
    .Y(_19703_));
 sky130_fd_sc_hd__nor2_4 _25951_ (.A(_19703_),
    .B(_19659_),
    .Y(_19704_));
 sky130_fd_sc_hd__a211o_4 _25952_ (.A1(\cpuregs[13][6] ),
    .A2(_19577_),
    .B1(_19702_),
    .C1(_19704_),
    .X(_19705_));
 sky130_fd_sc_hd__buf_1 _25953_ (.A(_19583_),
    .X(_19706_));
 sky130_fd_sc_hd__a21o_4 _25954_ (.A1(_19701_),
    .A2(_19705_),
    .B1(_19706_),
    .X(_19707_));
 sky130_vsdinv _25955_ (.A(\cpuregs[8][6] ),
    .Y(_19708_));
 sky130_fd_sc_hd__nor2_4 _25956_ (.A(_19708_),
    .B(_19590_),
    .Y(_19709_));
 sky130_fd_sc_hd__a211o_4 _25957_ (.A1(\cpuregs[9][6] ),
    .A2(_19586_),
    .B1(_19588_),
    .C1(_19709_),
    .X(_19710_));
 sky130_fd_sc_hd__buf_1 _25958_ (.A(_19286_),
    .X(_19711_));
 sky130_vsdinv _25959_ (.A(\cpuregs[10][6] ),
    .Y(_19712_));
 sky130_fd_sc_hd__nor2_4 _25960_ (.A(_19712_),
    .B(_19349_),
    .Y(_19713_));
 sky130_fd_sc_hd__a211o_4 _25961_ (.A1(\cpuregs[11][6] ),
    .A2(_19197_),
    .B1(_19711_),
    .C1(_19713_),
    .X(_19714_));
 sky130_fd_sc_hd__a21o_4 _25962_ (.A1(_19710_),
    .A2(_19714_),
    .B1(_19599_),
    .X(_19715_));
 sky130_fd_sc_hd__buf_1 _25963_ (.A(_19275_),
    .X(_19716_));
 sky130_fd_sc_hd__nand3_4 _25964_ (.A(_19707_),
    .B(_19715_),
    .C(_19716_),
    .Y(_19717_));
 sky130_fd_sc_hd__buf_1 _25965_ (.A(_19223_),
    .X(_19718_));
 sky130_fd_sc_hd__and2_4 _25966_ (.A(_19717_),
    .B(_19718_),
    .X(_19719_));
 sky130_fd_sc_hd__buf_1 _25967_ (.A(_19370_),
    .X(_19720_));
 sky130_fd_sc_hd__and2_4 _25968_ (.A(_19528_),
    .B(\cpuregs[0][6] ),
    .X(_19721_));
 sky130_fd_sc_hd__a211o_4 _25969_ (.A1(\cpuregs[1][6] ),
    .A2(_19605_),
    .B1(_19720_),
    .C1(_19721_),
    .X(_19722_));
 sky130_fd_sc_hd__buf_1 _25970_ (.A(_19533_),
    .X(_19723_));
 sky130_vsdinv _25971_ (.A(\cpuregs[2][6] ),
    .Y(_19724_));
 sky130_fd_sc_hd__nor2_4 _25972_ (.A(_19724_),
    .B(_19612_),
    .Y(_19725_));
 sky130_fd_sc_hd__a211o_4 _25973_ (.A1(\cpuregs[3][6] ),
    .A2(_19610_),
    .B1(_19723_),
    .C1(_19725_),
    .X(_19726_));
 sky130_fd_sc_hd__a21o_4 _25974_ (.A1(_19722_),
    .A2(_19726_),
    .B1(_19677_),
    .X(_19727_));
 sky130_fd_sc_hd__buf_1 _25975_ (.A(_19533_),
    .X(_19728_));
 sky130_vsdinv _25976_ (.A(\cpuregs[6][6] ),
    .Y(_19729_));
 sky130_fd_sc_hd__buf_1 _25977_ (.A(_19393_),
    .X(_19730_));
 sky130_fd_sc_hd__buf_1 _25978_ (.A(_19730_),
    .X(_19731_));
 sky130_fd_sc_hd__nor2_4 _25979_ (.A(_19729_),
    .B(_19731_),
    .Y(_19732_));
 sky130_fd_sc_hd__a211o_4 _25980_ (.A1(\cpuregs[7][6] ),
    .A2(_19557_),
    .B1(_19728_),
    .C1(_19732_),
    .X(_19733_));
 sky130_vsdinv _25981_ (.A(\cpuregs[4][6] ),
    .Y(_19734_));
 sky130_fd_sc_hd__nor2_4 _25982_ (.A(_19734_),
    .B(_19624_),
    .Y(_19735_));
 sky130_fd_sc_hd__a211o_4 _25983_ (.A1(\cpuregs[5][6] ),
    .A2(_19400_),
    .B1(_19371_),
    .C1(_19735_),
    .X(_19736_));
 sky130_fd_sc_hd__a21o_4 _25984_ (.A1(_19733_),
    .A2(_19736_),
    .B1(_19376_),
    .X(_19737_));
 sky130_fd_sc_hd__nand3_4 _25985_ (.A(_19727_),
    .B(_19358_),
    .C(_19737_),
    .Y(_19738_));
 sky130_fd_sc_hd__buf_1 _25986_ (.A(_19165_),
    .X(_19739_));
 sky130_fd_sc_hd__buf_1 _25987_ (.A(_19284_),
    .X(_19740_));
 sky130_fd_sc_hd__buf_1 _25988_ (.A(_19740_),
    .X(_19741_));
 sky130_vsdinv _25989_ (.A(\cpuregs[18][6] ),
    .Y(_19742_));
 sky130_fd_sc_hd__buf_1 _25990_ (.A(_19369_),
    .X(_19743_));
 sky130_fd_sc_hd__nor2_4 _25991_ (.A(_19742_),
    .B(_19743_),
    .Y(_19744_));
 sky130_fd_sc_hd__a211o_4 _25992_ (.A1(\cpuregs[19][6] ),
    .A2(_19741_),
    .B1(_19634_),
    .C1(_19744_),
    .X(_19745_));
 sky130_vsdinv _25993_ (.A(\cpuregs[16][6] ),
    .Y(_19746_));
 sky130_fd_sc_hd__nor2_4 _25994_ (.A(_19746_),
    .B(_19644_),
    .Y(_19747_));
 sky130_fd_sc_hd__a211o_4 _25995_ (.A1(\cpuregs[17][6] ),
    .A2(_19640_),
    .B1(_19641_),
    .C1(_19747_),
    .X(_19748_));
 sky130_fd_sc_hd__a21oi_4 _25996_ (.A1(_19745_),
    .A2(_19748_),
    .B1(_19647_),
    .Y(_19749_));
 sky130_fd_sc_hd__a2111o_4 _25997_ (.A1(_19719_),
    .A2(_19738_),
    .B1(_19739_),
    .C1(_19552_),
    .D1(_19749_),
    .X(_19750_));
 sky130_fd_sc_hd__xor2_4 _25998_ (.A(\timer[6] ),
    .B(_19696_),
    .X(_19751_));
 sky130_fd_sc_hd__nand2_4 _25999_ (.A(_19421_),
    .B(_19751_),
    .Y(_19752_));
 sky130_fd_sc_hd__buf_1 _26000_ (.A(_19495_),
    .X(_19753_));
 sky130_fd_sc_hd__a21oi_4 _26001_ (.A1(_19750_),
    .A2(_19752_),
    .B1(_19753_),
    .Y(_00654_));
 sky130_vsdinv _26002_ (.A(\cpuregs[14][7] ),
    .Y(_19754_));
 sky130_fd_sc_hd__nor2_4 _26003_ (.A(_19754_),
    .B(_19655_),
    .Y(_19755_));
 sky130_fd_sc_hd__a211o_4 _26004_ (.A1(\cpuregs[15][7] ),
    .A2(_19653_),
    .B1(_19201_),
    .C1(_19755_),
    .X(_19756_));
 sky130_vsdinv _26005_ (.A(\cpuregs[12][7] ),
    .Y(_19757_));
 sky130_fd_sc_hd__nor2_4 _26006_ (.A(_19757_),
    .B(_19659_),
    .Y(_19758_));
 sky130_fd_sc_hd__a211o_4 _26007_ (.A1(\cpuregs[13][7] ),
    .A2(_19577_),
    .B1(_19702_),
    .C1(_19758_),
    .X(_19759_));
 sky130_fd_sc_hd__a21o_4 _26008_ (.A1(_19756_),
    .A2(_19759_),
    .B1(_19706_),
    .X(_19760_));
 sky130_fd_sc_hd__buf_1 _26009_ (.A(_19318_),
    .X(_19761_));
 sky130_vsdinv _26010_ (.A(\cpuregs[8][7] ),
    .Y(_19762_));
 sky130_fd_sc_hd__nor2_4 _26011_ (.A(_19762_),
    .B(_19590_),
    .Y(_19763_));
 sky130_fd_sc_hd__a211o_4 _26012_ (.A1(\cpuregs[9][7] ),
    .A2(_19761_),
    .B1(_19588_),
    .C1(_19763_),
    .X(_19764_));
 sky130_vsdinv _26013_ (.A(\cpuregs[10][7] ),
    .Y(_19765_));
 sky130_fd_sc_hd__nor2_4 _26014_ (.A(_19765_),
    .B(_19349_),
    .Y(_19766_));
 sky130_fd_sc_hd__a211o_4 _26015_ (.A1(\cpuregs[11][7] ),
    .A2(_19197_),
    .B1(_19711_),
    .C1(_19766_),
    .X(_19767_));
 sky130_fd_sc_hd__a21o_4 _26016_ (.A1(_19764_),
    .A2(_19767_),
    .B1(_19599_),
    .X(_19768_));
 sky130_fd_sc_hd__nand3_4 _26017_ (.A(_19760_),
    .B(_19768_),
    .C(_19716_),
    .Y(_19769_));
 sky130_fd_sc_hd__and2_4 _26018_ (.A(_19769_),
    .B(_19718_),
    .X(_19770_));
 sky130_fd_sc_hd__and2_4 _26019_ (.A(_19528_),
    .B(\cpuregs[0][7] ),
    .X(_19771_));
 sky130_fd_sc_hd__a211o_4 _26020_ (.A1(\cpuregs[1][7] ),
    .A2(_19605_),
    .B1(_19720_),
    .C1(_19771_),
    .X(_19772_));
 sky130_fd_sc_hd__buf_1 _26021_ (.A(_19507_),
    .X(_19773_));
 sky130_vsdinv _26022_ (.A(\cpuregs[2][7] ),
    .Y(_19774_));
 sky130_fd_sc_hd__nor2_4 _26023_ (.A(_19774_),
    .B(_19612_),
    .Y(_19775_));
 sky130_fd_sc_hd__a211o_4 _26024_ (.A1(\cpuregs[3][7] ),
    .A2(_19773_),
    .B1(_19723_),
    .C1(_19775_),
    .X(_19776_));
 sky130_fd_sc_hd__a21o_4 _26025_ (.A1(_19772_),
    .A2(_19776_),
    .B1(_19677_),
    .X(_19777_));
 sky130_vsdinv _26026_ (.A(\cpuregs[6][7] ),
    .Y(_19778_));
 sky130_fd_sc_hd__nor2_4 _26027_ (.A(_19778_),
    .B(_19731_),
    .Y(_19779_));
 sky130_fd_sc_hd__a211o_4 _26028_ (.A1(\cpuregs[7][7] ),
    .A2(_19557_),
    .B1(_19728_),
    .C1(_19779_),
    .X(_19780_));
 sky130_vsdinv _26029_ (.A(\cpuregs[4][7] ),
    .Y(_19781_));
 sky130_fd_sc_hd__nor2_4 _26030_ (.A(_19781_),
    .B(_19547_),
    .Y(_19782_));
 sky130_fd_sc_hd__a211o_4 _26031_ (.A1(\cpuregs[5][7] ),
    .A2(_19400_),
    .B1(_19371_),
    .C1(_19782_),
    .X(_19783_));
 sky130_fd_sc_hd__a21o_4 _26032_ (.A1(_19780_),
    .A2(_19783_),
    .B1(_19376_),
    .X(_19784_));
 sky130_fd_sc_hd__nand3_4 _26033_ (.A(_19777_),
    .B(_19358_),
    .C(_19784_),
    .Y(_19785_));
 sky130_fd_sc_hd__buf_1 _26034_ (.A(_19383_),
    .X(_19786_));
 sky130_fd_sc_hd__buf_1 _26035_ (.A(_19320_),
    .X(_19787_));
 sky130_fd_sc_hd__buf_1 _26036_ (.A(_19787_),
    .X(_19788_));
 sky130_vsdinv _26037_ (.A(\cpuregs[18][7] ),
    .Y(_19789_));
 sky130_fd_sc_hd__nor2_4 _26038_ (.A(_19789_),
    .B(_19743_),
    .Y(_19790_));
 sky130_fd_sc_hd__a211o_4 _26039_ (.A1(\cpuregs[19][7] ),
    .A2(_19741_),
    .B1(_19788_),
    .C1(_19790_),
    .X(_19791_));
 sky130_fd_sc_hd__buf_1 _26040_ (.A(_19542_),
    .X(_19792_));
 sky130_vsdinv _26041_ (.A(\cpuregs[16][7] ),
    .Y(_19793_));
 sky130_fd_sc_hd__nor2_4 _26042_ (.A(_19793_),
    .B(_19644_),
    .Y(_19794_));
 sky130_fd_sc_hd__a211o_4 _26043_ (.A1(\cpuregs[17][7] ),
    .A2(_19640_),
    .B1(_19792_),
    .C1(_19794_),
    .X(_19795_));
 sky130_fd_sc_hd__buf_1 _26044_ (.A(_19409_),
    .X(_19796_));
 sky130_fd_sc_hd__a21oi_4 _26045_ (.A1(_19791_),
    .A2(_19795_),
    .B1(_19796_),
    .Y(_19797_));
 sky130_fd_sc_hd__a2111o_4 _26046_ (.A1(_19770_),
    .A2(_19785_),
    .B1(_19739_),
    .C1(_19786_),
    .D1(_19797_),
    .X(_19798_));
 sky130_fd_sc_hd__and4_4 _26047_ (.A(_19566_),
    .B(_19150_),
    .C(_19147_),
    .D(_18912_),
    .X(_19799_));
 sky130_fd_sc_hd__buf_1 _26048_ (.A(_19147_),
    .X(_19800_));
 sky130_fd_sc_hd__buf_1 _26049_ (.A(_19150_),
    .X(_19801_));
 sky130_fd_sc_hd__a41oi_4 _26050_ (.A1(_19800_),
    .A2(_19146_),
    .A3(_18917_),
    .A4(_18912_),
    .B1(_19801_),
    .Y(_19802_));
 sky130_fd_sc_hd__o21ai_4 _26051_ (.A1(_19799_),
    .A2(_19802_),
    .B1(_19492_),
    .Y(_19803_));
 sky130_fd_sc_hd__a21oi_4 _26052_ (.A1(_19798_),
    .A2(_19803_),
    .B1(_19753_),
    .Y(_00655_));
 sky130_fd_sc_hd__buf_1 _26053_ (.A(_19309_),
    .X(_19804_));
 sky130_fd_sc_hd__buf_1 _26054_ (.A(_19570_),
    .X(_19805_));
 sky130_vsdinv _26055_ (.A(\cpuregs[14][8] ),
    .Y(_19806_));
 sky130_fd_sc_hd__buf_1 _26056_ (.A(_19428_),
    .X(_19807_));
 sky130_fd_sc_hd__nor2_4 _26057_ (.A(_19806_),
    .B(_19807_),
    .Y(_19808_));
 sky130_fd_sc_hd__a211o_4 _26058_ (.A1(\cpuregs[15][8] ),
    .A2(_19804_),
    .B1(_19805_),
    .C1(_19808_),
    .X(_19809_));
 sky130_fd_sc_hd__buf_1 _26059_ (.A(_19587_),
    .X(_19810_));
 sky130_vsdinv _26060_ (.A(\cpuregs[12][8] ),
    .Y(_19811_));
 sky130_fd_sc_hd__buf_1 _26061_ (.A(_19291_),
    .X(_19812_));
 sky130_fd_sc_hd__nor2_4 _26062_ (.A(_19811_),
    .B(_19812_),
    .Y(_19813_));
 sky130_fd_sc_hd__a211o_4 _26063_ (.A1(\cpuregs[13][8] ),
    .A2(_19761_),
    .B1(_19810_),
    .C1(_19813_),
    .X(_19814_));
 sky130_fd_sc_hd__buf_1 _26064_ (.A(_19305_),
    .X(_19815_));
 sky130_fd_sc_hd__a21o_4 _26065_ (.A1(_19809_),
    .A2(_19814_),
    .B1(_19815_),
    .X(_19816_));
 sky130_fd_sc_hd__buf_1 _26066_ (.A(_19573_),
    .X(_19817_));
 sky130_vsdinv _26067_ (.A(\cpuregs[8][8] ),
    .Y(_19818_));
 sky130_fd_sc_hd__buf_1 _26068_ (.A(_19348_),
    .X(_19819_));
 sky130_fd_sc_hd__nor2_4 _26069_ (.A(_19818_),
    .B(_19819_),
    .Y(_19820_));
 sky130_fd_sc_hd__a211o_4 _26070_ (.A1(\cpuregs[9][8] ),
    .A2(_19817_),
    .B1(_19508_),
    .C1(_19820_),
    .X(_19821_));
 sky130_fd_sc_hd__buf_1 _26071_ (.A(_19333_),
    .X(_19822_));
 sky130_vsdinv _26072_ (.A(\cpuregs[10][8] ),
    .Y(_19823_));
 sky130_fd_sc_hd__nor2_4 _26073_ (.A(_19823_),
    .B(_19515_),
    .Y(_19824_));
 sky130_fd_sc_hd__a211o_4 _26074_ (.A1(\cpuregs[11][8] ),
    .A2(_19822_),
    .B1(_19513_),
    .C1(_19824_),
    .X(_19825_));
 sky130_fd_sc_hd__buf_1 _26075_ (.A(_19353_),
    .X(_19826_));
 sky130_fd_sc_hd__a21o_4 _26076_ (.A1(_19821_),
    .A2(_19825_),
    .B1(_19826_),
    .X(_19827_));
 sky130_fd_sc_hd__nand3_4 _26077_ (.A(_19816_),
    .B(_19827_),
    .C(_19520_),
    .Y(_19828_));
 sky130_fd_sc_hd__and2_4 _26078_ (.A(_19828_),
    .B(_19522_),
    .X(_19829_));
 sky130_fd_sc_hd__buf_1 _26079_ (.A(_19311_),
    .X(_19830_));
 sky130_fd_sc_hd__buf_1 _26080_ (.A(_19830_),
    .X(_19831_));
 sky130_fd_sc_hd__and2_4 _26081_ (.A(_19528_),
    .B(\cpuregs[0][8] ),
    .X(_19832_));
 sky130_fd_sc_hd__a211o_4 _26082_ (.A1(\cpuregs[1][8] ),
    .A2(_19343_),
    .B1(_19831_),
    .C1(_19832_),
    .X(_19833_));
 sky130_vsdinv _26083_ (.A(\cpuregs[2][8] ),
    .Y(_19834_));
 sky130_fd_sc_hd__nor2_4 _26084_ (.A(_19834_),
    .B(_19731_),
    .Y(_19835_));
 sky130_fd_sc_hd__a211o_4 _26085_ (.A1(\cpuregs[3][8] ),
    .A2(_19387_),
    .B1(_19728_),
    .C1(_19835_),
    .X(_19836_));
 sky130_fd_sc_hd__a21o_4 _26086_ (.A1(_19833_),
    .A2(_19836_),
    .B1(_19677_),
    .X(_19837_));
 sky130_fd_sc_hd__buf_1 _26087_ (.A(_19357_),
    .X(_19838_));
 sky130_fd_sc_hd__buf_1 _26088_ (.A(_19359_),
    .X(_19839_));
 sky130_vsdinv _26089_ (.A(\cpuregs[6][8] ),
    .Y(_19840_));
 sky130_fd_sc_hd__buf_1 _26090_ (.A(_19623_),
    .X(_19841_));
 sky130_fd_sc_hd__nor2_4 _26091_ (.A(_19840_),
    .B(_19841_),
    .Y(_19842_));
 sky130_fd_sc_hd__a211o_4 _26092_ (.A1(\cpuregs[7][8] ),
    .A2(_19839_),
    .B1(_19361_),
    .C1(_19842_),
    .X(_19843_));
 sky130_fd_sc_hd__buf_1 _26093_ (.A(_19291_),
    .X(_19844_));
 sky130_fd_sc_hd__buf_1 _26094_ (.A(_19844_),
    .X(_19845_));
 sky130_fd_sc_hd__buf_1 _26095_ (.A(_19541_),
    .X(_19846_));
 sky130_vsdinv _26096_ (.A(\cpuregs[4][8] ),
    .Y(_19847_));
 sky130_fd_sc_hd__nor2_4 _26097_ (.A(_19847_),
    .B(_19229_),
    .Y(_19848_));
 sky130_fd_sc_hd__a211o_4 _26098_ (.A1(\cpuregs[5][8] ),
    .A2(_19845_),
    .B1(_19846_),
    .C1(_19848_),
    .X(_19849_));
 sky130_fd_sc_hd__buf_1 _26099_ (.A(_19250_),
    .X(_19850_));
 sky130_fd_sc_hd__buf_1 _26100_ (.A(_19850_),
    .X(_19851_));
 sky130_fd_sc_hd__a21o_4 _26101_ (.A1(_19843_),
    .A2(_19849_),
    .B1(_19851_),
    .X(_19852_));
 sky130_fd_sc_hd__nand3_4 _26102_ (.A(_19837_),
    .B(_19838_),
    .C(_19852_),
    .Y(_19853_));
 sky130_fd_sc_hd__buf_1 _26103_ (.A(_19639_),
    .X(_19854_));
 sky130_vsdinv _26104_ (.A(\cpuregs[18][8] ),
    .Y(_19855_));
 sky130_fd_sc_hd__buf_1 _26105_ (.A(_19643_),
    .X(_19856_));
 sky130_fd_sc_hd__nor2_4 _26106_ (.A(_19855_),
    .B(_19856_),
    .Y(_19857_));
 sky130_fd_sc_hd__a211o_4 _26107_ (.A1(\cpuregs[19][8] ),
    .A2(_19854_),
    .B1(_19788_),
    .C1(_19857_),
    .X(_19858_));
 sky130_vsdinv _26108_ (.A(\cpuregs[16][8] ),
    .Y(_19859_));
 sky130_fd_sc_hd__nor2_4 _26109_ (.A(_19859_),
    .B(_19396_),
    .Y(_19860_));
 sky130_fd_sc_hd__a211o_4 _26110_ (.A1(\cpuregs[17][8] ),
    .A2(_19388_),
    .B1(_19792_),
    .C1(_19860_),
    .X(_19861_));
 sky130_fd_sc_hd__a21oi_4 _26111_ (.A1(_19858_),
    .A2(_19861_),
    .B1(_19796_),
    .Y(_19862_));
 sky130_fd_sc_hd__a2111o_4 _26112_ (.A1(_19829_),
    .A2(_19853_),
    .B1(_19739_),
    .C1(_19786_),
    .D1(_19862_),
    .X(_19863_));
 sky130_fd_sc_hd__and4_4 _26113_ (.A(_19696_),
    .B(_19149_),
    .C(_19150_),
    .D(_19800_),
    .X(_19864_));
 sky130_fd_sc_hd__buf_1 _26114_ (.A(_19149_),
    .X(_19865_));
 sky130_fd_sc_hd__a41oi_4 _26115_ (.A1(_19801_),
    .A2(_19566_),
    .A3(_19800_),
    .A4(_18912_),
    .B1(_19865_),
    .Y(_19866_));
 sky130_fd_sc_hd__buf_1 _26116_ (.A(_19419_),
    .X(_19867_));
 sky130_fd_sc_hd__o21ai_4 _26117_ (.A1(_19864_),
    .A2(_19866_),
    .B1(_19867_),
    .Y(_19868_));
 sky130_fd_sc_hd__a21oi_4 _26118_ (.A1(_19863_),
    .A2(_19868_),
    .B1(_19753_),
    .Y(_00656_));
 sky130_vsdinv _26119_ (.A(\cpuregs[14][9] ),
    .Y(_19869_));
 sky130_fd_sc_hd__nor2_4 _26120_ (.A(_19869_),
    .B(_19807_),
    .Y(_19870_));
 sky130_fd_sc_hd__a211o_4 _26121_ (.A1(\cpuregs[15][9] ),
    .A2(_19804_),
    .B1(_19805_),
    .C1(_19870_),
    .X(_19871_));
 sky130_vsdinv _26122_ (.A(\cpuregs[12][9] ),
    .Y(_19872_));
 sky130_fd_sc_hd__nor2_4 _26123_ (.A(_19872_),
    .B(_19812_),
    .Y(_19873_));
 sky130_fd_sc_hd__a211o_4 _26124_ (.A1(\cpuregs[13][9] ),
    .A2(_19761_),
    .B1(_19810_),
    .C1(_19873_),
    .X(_19874_));
 sky130_fd_sc_hd__a21o_4 _26125_ (.A1(_19871_),
    .A2(_19874_),
    .B1(_19815_),
    .X(_19875_));
 sky130_fd_sc_hd__buf_1 _26126_ (.A(_19298_),
    .X(_19876_));
 sky130_vsdinv _26127_ (.A(\cpuregs[8][9] ),
    .Y(_19877_));
 sky130_fd_sc_hd__buf_1 _26128_ (.A(_19301_),
    .X(_19878_));
 sky130_fd_sc_hd__nor2_4 _26129_ (.A(_19877_),
    .B(_19878_),
    .Y(_19879_));
 sky130_fd_sc_hd__a211o_4 _26130_ (.A1(\cpuregs[9][9] ),
    .A2(_19817_),
    .B1(_19876_),
    .C1(_19879_),
    .X(_19880_));
 sky130_vsdinv _26131_ (.A(\cpuregs[10][9] ),
    .Y(_19881_));
 sky130_fd_sc_hd__buf_1 _26132_ (.A(_19393_),
    .X(_19882_));
 sky130_fd_sc_hd__nor2_4 _26133_ (.A(_19881_),
    .B(_19882_),
    .Y(_19883_));
 sky130_fd_sc_hd__a211o_4 _26134_ (.A1(\cpuregs[11][9] ),
    .A2(_19822_),
    .B1(_19513_),
    .C1(_19883_),
    .X(_19884_));
 sky130_fd_sc_hd__a21o_4 _26135_ (.A1(_19880_),
    .A2(_19884_),
    .B1(_19826_),
    .X(_19885_));
 sky130_fd_sc_hd__nand3_4 _26136_ (.A(_19875_),
    .B(_19885_),
    .C(_19520_),
    .Y(_19886_));
 sky130_fd_sc_hd__buf_1 _26137_ (.A(_19223_),
    .X(_19887_));
 sky130_fd_sc_hd__and2_4 _26138_ (.A(_19886_),
    .B(_19887_),
    .X(_19888_));
 sky130_fd_sc_hd__buf_1 _26139_ (.A(_19217_),
    .X(_19889_));
 sky130_fd_sc_hd__and2_4 _26140_ (.A(_19889_),
    .B(\cpuregs[0][9] ),
    .X(_19890_));
 sky130_fd_sc_hd__a211o_4 _26141_ (.A1(\cpuregs[1][9] ),
    .A2(_19343_),
    .B1(_19831_),
    .C1(_19890_),
    .X(_19891_));
 sky130_fd_sc_hd__buf_1 _26142_ (.A(_19555_),
    .X(_19892_));
 sky130_fd_sc_hd__buf_1 _26143_ (.A(_19892_),
    .X(_19893_));
 sky130_vsdinv _26144_ (.A(\cpuregs[2][9] ),
    .Y(_19894_));
 sky130_fd_sc_hd__nor2_4 _26145_ (.A(_19894_),
    .B(_19731_),
    .Y(_19895_));
 sky130_fd_sc_hd__a211o_4 _26146_ (.A1(\cpuregs[3][9] ),
    .A2(_19893_),
    .B1(_19728_),
    .C1(_19895_),
    .X(_19896_));
 sky130_fd_sc_hd__buf_1 _26147_ (.A(_19826_),
    .X(_19897_));
 sky130_fd_sc_hd__a21o_4 _26148_ (.A1(_19891_),
    .A2(_19896_),
    .B1(_19897_),
    .X(_19898_));
 sky130_fd_sc_hd__buf_1 _26149_ (.A(_19394_),
    .X(_19899_));
 sky130_vsdinv _26150_ (.A(\cpuregs[6][9] ),
    .Y(_19900_));
 sky130_fd_sc_hd__nor2_4 _26151_ (.A(_19900_),
    .B(_19841_),
    .Y(_19901_));
 sky130_fd_sc_hd__a211o_4 _26152_ (.A1(\cpuregs[7][9] ),
    .A2(_19899_),
    .B1(_19361_),
    .C1(_19901_),
    .X(_19902_));
 sky130_vsdinv _26153_ (.A(\cpuregs[4][9] ),
    .Y(_19903_));
 sky130_fd_sc_hd__nor2_4 _26154_ (.A(_19903_),
    .B(_19229_),
    .Y(_19904_));
 sky130_fd_sc_hd__a211o_4 _26155_ (.A1(\cpuregs[5][9] ),
    .A2(_19845_),
    .B1(_19846_),
    .C1(_19904_),
    .X(_19905_));
 sky130_fd_sc_hd__a21o_4 _26156_ (.A1(_19902_),
    .A2(_19905_),
    .B1(_19851_),
    .X(_19906_));
 sky130_fd_sc_hd__nand3_4 _26157_ (.A(_19898_),
    .B(_19838_),
    .C(_19906_),
    .Y(_19907_));
 sky130_fd_sc_hd__buf_1 _26158_ (.A(_19787_),
    .X(_19908_));
 sky130_vsdinv _26159_ (.A(\cpuregs[18][9] ),
    .Y(_19909_));
 sky130_fd_sc_hd__nor2_4 _26160_ (.A(_19909_),
    .B(_19856_),
    .Y(_19910_));
 sky130_fd_sc_hd__a211o_4 _26161_ (.A1(\cpuregs[19][9] ),
    .A2(_19854_),
    .B1(_19908_),
    .C1(_19910_),
    .X(_19911_));
 sky130_fd_sc_hd__buf_1 _26162_ (.A(_19387_),
    .X(_19912_));
 sky130_fd_sc_hd__buf_1 _26163_ (.A(_19542_),
    .X(_19913_));
 sky130_vsdinv _26164_ (.A(\cpuregs[16][9] ),
    .Y(_19914_));
 sky130_fd_sc_hd__buf_1 _26165_ (.A(_19395_),
    .X(_19915_));
 sky130_fd_sc_hd__nor2_4 _26166_ (.A(_19914_),
    .B(_19915_),
    .Y(_19916_));
 sky130_fd_sc_hd__a211o_4 _26167_ (.A1(\cpuregs[17][9] ),
    .A2(_19912_),
    .B1(_19913_),
    .C1(_19916_),
    .X(_19917_));
 sky130_fd_sc_hd__buf_1 _26168_ (.A(_19409_),
    .X(_19918_));
 sky130_fd_sc_hd__a21oi_4 _26169_ (.A1(_19911_),
    .A2(_19917_),
    .B1(_19918_),
    .Y(_19919_));
 sky130_fd_sc_hd__a2111o_4 _26170_ (.A1(_19888_),
    .A2(_19907_),
    .B1(_19739_),
    .C1(_19786_),
    .D1(_19919_),
    .X(_19920_));
 sky130_vsdinv _26171_ (.A(\timer[9] ),
    .Y(_19921_));
 sky130_fd_sc_hd__a41oi_4 _26172_ (.A1(_19865_),
    .A2(_19696_),
    .A3(_19801_),
    .A4(_19800_),
    .B1(_19921_),
    .Y(_19922_));
 sky130_fd_sc_hd__and4_4 _26173_ (.A(_19148_),
    .B(_19921_),
    .C(_19865_),
    .D(_19801_),
    .X(_19923_));
 sky130_fd_sc_hd__o21ai_4 _26174_ (.A1(_19922_),
    .A2(_19923_),
    .B1(_19867_),
    .Y(_19924_));
 sky130_fd_sc_hd__a21oi_4 _26175_ (.A1(_19920_),
    .A2(_19924_),
    .B1(_19753_),
    .Y(_00657_));
 sky130_fd_sc_hd__buf_1 _26176_ (.A(_19415_),
    .X(_19925_));
 sky130_fd_sc_hd__buf_1 _26177_ (.A(_19157_),
    .X(_19926_));
 sky130_vsdinv _26178_ (.A(_19152_),
    .Y(_19927_));
 sky130_fd_sc_hd__a41oi_4 _26179_ (.A1(_19925_),
    .A2(_19416_),
    .A3(_19417_),
    .A4(_19926_),
    .B1(_19927_),
    .Y(_19928_));
 sky130_vsdinv _26180_ (.A(_19928_),
    .Y(_19929_));
 sky130_vsdinv _26181_ (.A(_19923_),
    .Y(_19930_));
 sky130_fd_sc_hd__buf_1 _26182_ (.A(_19418_),
    .X(_19931_));
 sky130_fd_sc_hd__buf_1 _26183_ (.A(_19931_),
    .X(_19932_));
 sky130_fd_sc_hd__a21oi_4 _26184_ (.A1(_19930_),
    .A2(\timer[10] ),
    .B1(_19932_),
    .Y(_19933_));
 sky130_fd_sc_hd__and2_4 _26185_ (.A(_19217_),
    .B(\cpuregs[0][10] ),
    .X(_19934_));
 sky130_fd_sc_hd__a211o_4 _26186_ (.A1(\cpuregs[1][10] ),
    .A2(_19297_),
    .B1(_19312_),
    .C1(_19934_),
    .X(_19935_));
 sky130_fd_sc_hd__buf_1 _26187_ (.A(_19367_),
    .X(_19936_));
 sky130_vsdinv _26188_ (.A(\cpuregs[2][10] ),
    .Y(_19937_));
 sky130_fd_sc_hd__nor2_4 _26189_ (.A(_19937_),
    .B(_19315_),
    .Y(_19938_));
 sky130_fd_sc_hd__a211o_4 _26190_ (.A1(\cpuregs[3][10] ),
    .A2(_19936_),
    .B1(_19389_),
    .C1(_19938_),
    .X(_19939_));
 sky130_fd_sc_hd__a21o_4 _26191_ (.A1(_19935_),
    .A2(_19939_),
    .B1(_19240_),
    .X(_19940_));
 sky130_vsdinv _26192_ (.A(\cpuregs[6][10] ),
    .Y(_19941_));
 sky130_fd_sc_hd__nor2_4 _26193_ (.A(_19941_),
    .B(_19228_),
    .Y(_19942_));
 sky130_fd_sc_hd__a211o_4 _26194_ (.A1(\cpuregs[7][10] ),
    .A2(_19342_),
    .B1(_19345_),
    .C1(_19942_),
    .X(_19943_));
 sky130_fd_sc_hd__buf_1 _26195_ (.A(_19311_),
    .X(_19944_));
 sky130_vsdinv _26196_ (.A(\cpuregs[4][10] ),
    .Y(_19945_));
 sky130_fd_sc_hd__nor2_4 _26197_ (.A(_19945_),
    .B(_19172_),
    .Y(_19946_));
 sky130_fd_sc_hd__a211o_4 _26198_ (.A1(\cpuregs[5][10] ),
    .A2(_19556_),
    .B1(_19944_),
    .C1(_19946_),
    .X(_19947_));
 sky130_fd_sc_hd__a21o_4 _26199_ (.A1(_19943_),
    .A2(_19947_),
    .B1(_19251_),
    .X(_19948_));
 sky130_fd_sc_hd__nand3_4 _26200_ (.A(_19940_),
    .B(_19254_),
    .C(_19948_),
    .Y(_19949_));
 sky130_vsdinv _26201_ (.A(\cpuregs[14][10] ),
    .Y(_19950_));
 sky130_fd_sc_hd__nor2_4 _26202_ (.A(_19950_),
    .B(_19322_),
    .Y(_19951_));
 sky130_fd_sc_hd__a211o_4 _26203_ (.A1(\cpuregs[15][10] ),
    .A2(_19368_),
    .B1(_19320_),
    .C1(_19951_),
    .X(_19952_));
 sky130_vsdinv _26204_ (.A(\cpuregs[12][10] ),
    .Y(_19953_));
 sky130_fd_sc_hd__nor2_4 _26205_ (.A(_19953_),
    .B(_19257_),
    .Y(_19954_));
 sky130_fd_sc_hd__a211o_4 _26206_ (.A1(\cpuregs[13][10] ),
    .A2(_19574_),
    .B1(_19830_),
    .C1(_19954_),
    .X(_19955_));
 sky130_fd_sc_hd__a21o_4 _26207_ (.A1(_19952_),
    .A2(_19955_),
    .B1(_19850_),
    .X(_19956_));
 sky130_vsdinv _26208_ (.A(\cpuregs[8][10] ),
    .Y(_19957_));
 sky130_fd_sc_hd__nor2_4 _26209_ (.A(_19957_),
    .B(_19172_),
    .Y(_19958_));
 sky130_fd_sc_hd__a211o_4 _26210_ (.A1(\cpuregs[9][10] ),
    .A2(_19892_),
    .B1(_19944_),
    .C1(_19958_),
    .X(_19959_));
 sky130_vsdinv _26211_ (.A(\cpuregs[10][10] ),
    .Y(_19960_));
 sky130_fd_sc_hd__nor2_4 _26212_ (.A(_19960_),
    .B(_19234_),
    .Y(_19961_));
 sky130_fd_sc_hd__a211o_4 _26213_ (.A1(\cpuregs[11][10] ),
    .A2(_19399_),
    .B1(_19230_),
    .C1(_19961_),
    .X(_19962_));
 sky130_fd_sc_hd__a21o_4 _26214_ (.A1(_19959_),
    .A2(_19962_),
    .B1(_19263_),
    .X(_19963_));
 sky130_fd_sc_hd__nand3_4 _26215_ (.A(_19956_),
    .B(_19963_),
    .C(_19327_),
    .Y(_19964_));
 sky130_fd_sc_hd__nand3_4 _26216_ (.A(_19949_),
    .B(_19522_),
    .C(_19964_),
    .Y(_19965_));
 sky130_vsdinv _26217_ (.A(\cpuregs[18][10] ),
    .Y(_19966_));
 sky130_fd_sc_hd__nor2_4 _26218_ (.A(_19966_),
    .B(_19547_),
    .Y(_19967_));
 sky130_fd_sc_hd__a211o_4 _26219_ (.A1(\cpuregs[19][10] ),
    .A2(_19369_),
    .B1(_19231_),
    .C1(_19967_),
    .X(_19968_));
 sky130_fd_sc_hd__buf_1 _26220_ (.A(_19531_),
    .X(_19969_));
 sky130_vsdinv _26221_ (.A(\cpuregs[16][10] ),
    .Y(_19970_));
 sky130_fd_sc_hd__nor2_4 _26222_ (.A(_19970_),
    .B(_19258_),
    .Y(_19971_));
 sky130_fd_sc_hd__a211o_4 _26223_ (.A1(\cpuregs[17][10] ),
    .A2(_19969_),
    .B1(_19237_),
    .C1(_19971_),
    .X(_19972_));
 sky130_fd_sc_hd__a21oi_4 _26224_ (.A1(_19968_),
    .A2(_19972_),
    .B1(_19278_),
    .Y(_19973_));
 sky130_fd_sc_hd__nor2_4 _26225_ (.A(_19381_),
    .B(_19973_),
    .Y(_19974_));
 sky130_fd_sc_hd__nand2_4 _26226_ (.A(_19965_),
    .B(_19974_),
    .Y(_19975_));
 sky130_fd_sc_hd__buf_1 _26227_ (.A(_19418_),
    .X(_19976_));
 sky130_fd_sc_hd__buf_1 _26228_ (.A(_18478_),
    .X(_19977_));
 sky130_fd_sc_hd__a21o_4 _26229_ (.A1(_19975_),
    .A2(_19976_),
    .B1(_19977_),
    .X(_19978_));
 sky130_fd_sc_hd__a21oi_4 _26230_ (.A1(_19929_),
    .A2(_19933_),
    .B1(_19978_),
    .Y(_00627_));
 sky130_fd_sc_hd__buf_1 _26231_ (.A(_19153_),
    .X(_19979_));
 sky130_fd_sc_hd__nand2_4 _26232_ (.A(_19928_),
    .B(_19979_),
    .Y(_19980_));
 sky130_vsdinv _26233_ (.A(_19980_),
    .Y(_19981_));
 sky130_fd_sc_hd__o21ai_4 _26234_ (.A1(_19979_),
    .A2(_19152_),
    .B1(_19380_),
    .Y(_19982_));
 sky130_fd_sc_hd__buf_1 _26235_ (.A(_19511_),
    .X(_19983_));
 sky130_vsdinv _26236_ (.A(\cpuregs[14][11] ),
    .Y(_19984_));
 sky130_fd_sc_hd__buf_1 _26237_ (.A(_19555_),
    .X(_19985_));
 sky130_fd_sc_hd__nor2_4 _26238_ (.A(_19984_),
    .B(_19985_),
    .Y(_19986_));
 sky130_fd_sc_hd__a211o_4 _26239_ (.A1(\cpuregs[15][11] ),
    .A2(_19983_),
    .B1(_19201_),
    .C1(_19986_),
    .X(_19987_));
 sky130_fd_sc_hd__buf_1 _26240_ (.A(_19524_),
    .X(_19988_));
 sky130_vsdinv _26241_ (.A(\cpuregs[12][11] ),
    .Y(_19989_));
 sky130_fd_sc_hd__buf_1 _26242_ (.A(_19341_),
    .X(_19990_));
 sky130_fd_sc_hd__nor2_4 _26243_ (.A(_19989_),
    .B(_19990_),
    .Y(_19991_));
 sky130_fd_sc_hd__a211o_4 _26244_ (.A1(\cpuregs[13][11] ),
    .A2(_19988_),
    .B1(_19702_),
    .C1(_19991_),
    .X(_19992_));
 sky130_fd_sc_hd__a21o_4 _26245_ (.A1(_19987_),
    .A2(_19992_),
    .B1(_19706_),
    .X(_19993_));
 sky130_fd_sc_hd__buf_1 _26246_ (.A(_19298_),
    .X(_19994_));
 sky130_vsdinv _26247_ (.A(\cpuregs[8][11] ),
    .Y(_19995_));
 sky130_fd_sc_hd__nor2_4 _26248_ (.A(_19995_),
    .B(_19844_),
    .Y(_19996_));
 sky130_fd_sc_hd__a211o_4 _26249_ (.A1(\cpuregs[9][11] ),
    .A2(_19284_),
    .B1(_19994_),
    .C1(_19996_),
    .X(_19997_));
 sky130_vsdinv _26250_ (.A(\cpuregs[10][11] ),
    .Y(_19998_));
 sky130_fd_sc_hd__nor2_4 _26251_ (.A(_19998_),
    .B(_19302_),
    .Y(_19999_));
 sky130_fd_sc_hd__a211o_4 _26252_ (.A1(\cpuregs[11][11] ),
    .A2(_19297_),
    .B1(_19711_),
    .C1(_19999_),
    .X(_20000_));
 sky130_fd_sc_hd__buf_1 _26253_ (.A(_19472_),
    .X(_20001_));
 sky130_fd_sc_hd__a21o_4 _26254_ (.A1(_19997_),
    .A2(_20000_),
    .B1(_20001_),
    .X(_20002_));
 sky130_fd_sc_hd__nand3_4 _26255_ (.A(_19993_),
    .B(_20002_),
    .C(_19716_),
    .Y(_20003_));
 sky130_fd_sc_hd__and2_4 _26256_ (.A(_20003_),
    .B(_19718_),
    .X(_20004_));
 sky130_fd_sc_hd__buf_1 _26257_ (.A(_19936_),
    .X(_20005_));
 sky130_fd_sc_hd__buf_1 _26258_ (.A(_19312_),
    .X(_20006_));
 sky130_fd_sc_hd__buf_1 _26259_ (.A(_19337_),
    .X(_20007_));
 sky130_fd_sc_hd__and2_4 _26260_ (.A(_20007_),
    .B(\cpuregs[0][11] ),
    .X(_20008_));
 sky130_fd_sc_hd__a211o_4 _26261_ (.A1(\cpuregs[1][11] ),
    .A2(_20005_),
    .B1(_20006_),
    .C1(_20008_),
    .X(_20009_));
 sky130_fd_sc_hd__buf_1 _26262_ (.A(_19345_),
    .X(_20010_));
 sky130_vsdinv _26263_ (.A(\cpuregs[2][11] ),
    .Y(_20011_));
 sky130_fd_sc_hd__buf_1 _26264_ (.A(_19819_),
    .X(_20012_));
 sky130_fd_sc_hd__nor2_4 _26265_ (.A(_20011_),
    .B(_20012_),
    .Y(_20013_));
 sky130_fd_sc_hd__a211o_4 _26266_ (.A1(\cpuregs[3][11] ),
    .A2(_19526_),
    .B1(_20010_),
    .C1(_20013_),
    .X(_20014_));
 sky130_fd_sc_hd__buf_1 _26267_ (.A(_19353_),
    .X(_20015_));
 sky130_fd_sc_hd__buf_1 _26268_ (.A(_20015_),
    .X(_20016_));
 sky130_fd_sc_hd__a21o_4 _26269_ (.A1(_20009_),
    .A2(_20014_),
    .B1(_20016_),
    .X(_20017_));
 sky130_fd_sc_hd__buf_1 _26270_ (.A(_19476_),
    .X(_20018_));
 sky130_vsdinv _26271_ (.A(\cpuregs[6][11] ),
    .Y(_20019_));
 sky130_fd_sc_hd__nor2_4 _26272_ (.A(_20019_),
    .B(_19440_),
    .Y(_20020_));
 sky130_fd_sc_hd__a211o_4 _26273_ (.A1(\cpuregs[7][11] ),
    .A2(_19773_),
    .B1(_19723_),
    .C1(_20020_),
    .X(_20021_));
 sky130_fd_sc_hd__buf_1 _26274_ (.A(_19359_),
    .X(_20022_));
 sky130_vsdinv _26275_ (.A(\cpuregs[4][11] ),
    .Y(_20023_));
 sky130_fd_sc_hd__nor2_4 _26276_ (.A(_20023_),
    .B(_19363_),
    .Y(_20024_));
 sky130_fd_sc_hd__a211o_4 _26277_ (.A1(\cpuregs[5][11] ),
    .A2(_20022_),
    .B1(_19542_),
    .C1(_20024_),
    .X(_20025_));
 sky130_fd_sc_hd__buf_1 _26278_ (.A(_19375_),
    .X(_20026_));
 sky130_fd_sc_hd__a21o_4 _26279_ (.A1(_20021_),
    .A2(_20025_),
    .B1(_20026_),
    .X(_20027_));
 sky130_fd_sc_hd__nand3_4 _26280_ (.A(_20017_),
    .B(_20018_),
    .C(_20027_),
    .Y(_20028_));
 sky130_fd_sc_hd__buf_1 _26281_ (.A(_19192_),
    .X(_20029_));
 sky130_fd_sc_hd__buf_1 _26282_ (.A(_20029_),
    .X(_20030_));
 sky130_fd_sc_hd__buf_1 _26283_ (.A(_20030_),
    .X(_20031_));
 sky130_fd_sc_hd__buf_1 _26284_ (.A(_19936_),
    .X(_20032_));
 sky130_fd_sc_hd__buf_1 _26285_ (.A(_20032_),
    .X(_20033_));
 sky130_fd_sc_hd__buf_1 _26286_ (.A(_19200_),
    .X(_20034_));
 sky130_fd_sc_hd__buf_1 _26287_ (.A(_20034_),
    .X(_20035_));
 sky130_fd_sc_hd__buf_1 _26288_ (.A(_20035_),
    .X(_20036_));
 sky130_vsdinv _26289_ (.A(\cpuregs[18][11] ),
    .Y(_20037_));
 sky130_fd_sc_hd__buf_1 _26290_ (.A(_19545_),
    .X(_20038_));
 sky130_fd_sc_hd__nor2_4 _26291_ (.A(_20037_),
    .B(_20038_),
    .Y(_20039_));
 sky130_fd_sc_hd__a211o_4 _26292_ (.A1(\cpuregs[19][11] ),
    .A2(_20033_),
    .B1(_20036_),
    .C1(_20039_),
    .X(_20040_));
 sky130_fd_sc_hd__buf_1 _26293_ (.A(_19526_),
    .X(_20041_));
 sky130_fd_sc_hd__buf_1 _26294_ (.A(_19527_),
    .X(_20042_));
 sky130_vsdinv _26295_ (.A(\cpuregs[16][11] ),
    .Y(_20043_));
 sky130_fd_sc_hd__buf_1 _26296_ (.A(_19655_),
    .X(_20044_));
 sky130_fd_sc_hd__buf_1 _26297_ (.A(_20044_),
    .X(_20045_));
 sky130_fd_sc_hd__nor2_4 _26298_ (.A(_20043_),
    .B(_20045_),
    .Y(_20046_));
 sky130_fd_sc_hd__a211o_4 _26299_ (.A1(\cpuregs[17][11] ),
    .A2(_20041_),
    .B1(_20042_),
    .C1(_20046_),
    .X(_20047_));
 sky130_fd_sc_hd__buf_1 _26300_ (.A(_19224_),
    .X(_20048_));
 sky130_fd_sc_hd__a21oi_4 _26301_ (.A1(_20040_),
    .A2(_20047_),
    .B1(_20048_),
    .Y(_20049_));
 sky130_fd_sc_hd__a211o_4 _26302_ (.A1(_20004_),
    .A2(_20028_),
    .B1(_20031_),
    .C1(_20049_),
    .X(_20050_));
 sky130_fd_sc_hd__buf_1 _26303_ (.A(_19931_),
    .X(_20051_));
 sky130_fd_sc_hd__a21oi_4 _26304_ (.A1(_20050_),
    .A2(_20051_),
    .B1(_18229_),
    .Y(_20052_));
 sky130_fd_sc_hd__o21a_4 _26305_ (.A1(_19981_),
    .A2(_19982_),
    .B1(_20052_),
    .X(_00628_));
 sky130_fd_sc_hd__nor4_4 _26306_ (.A(\timer[11] ),
    .B(\timer[12] ),
    .C(_19927_),
    .D(_19161_),
    .Y(_20053_));
 sky130_fd_sc_hd__buf_1 _26307_ (.A(_19155_),
    .X(_20054_));
 sky130_fd_sc_hd__and4_4 _26308_ (.A(_19799_),
    .B(_19865_),
    .C(_19153_),
    .D(_18910_),
    .X(_20055_));
 sky130_fd_sc_hd__o21ai_4 _26309_ (.A1(_20054_),
    .A2(_20055_),
    .B1(_19380_),
    .Y(_20056_));
 sky130_fd_sc_hd__buf_1 _26310_ (.A(_19480_),
    .X(_20057_));
 sky130_fd_sc_hd__buf_1 _26311_ (.A(_19455_),
    .X(_20058_));
 sky130_vsdinv _26312_ (.A(\cpuregs[14][12] ),
    .Y(_20059_));
 sky130_fd_sc_hd__nor2_4 _26313_ (.A(_20059_),
    .B(_19310_),
    .Y(_20060_));
 sky130_fd_sc_hd__a211o_4 _26314_ (.A1(\cpuregs[15][12] ),
    .A2(_20057_),
    .B1(_20058_),
    .C1(_20060_),
    .X(_20061_));
 sky130_vsdinv _26315_ (.A(\cpuregs[12][12] ),
    .Y(_20062_));
 sky130_fd_sc_hd__nor2_4 _26316_ (.A(_20062_),
    .B(_19319_),
    .Y(_20063_));
 sky130_fd_sc_hd__a211o_4 _26317_ (.A1(\cpuregs[13][12] ),
    .A2(_19445_),
    .B1(_19271_),
    .C1(_20063_),
    .X(_20064_));
 sky130_fd_sc_hd__buf_1 _26318_ (.A(_19583_),
    .X(_20065_));
 sky130_fd_sc_hd__a21o_4 _26319_ (.A1(_20061_),
    .A2(_20064_),
    .B1(_20065_),
    .X(_20066_));
 sky130_fd_sc_hd__buf_1 _26320_ (.A(_19511_),
    .X(_20067_));
 sky130_fd_sc_hd__buf_1 _26321_ (.A(_19213_),
    .X(_20068_));
 sky130_vsdinv _26322_ (.A(\cpuregs[8][12] ),
    .Y(_20069_));
 sky130_fd_sc_hd__nor2_4 _26323_ (.A(_20069_),
    .B(_19386_),
    .Y(_20070_));
 sky130_fd_sc_hd__a211o_4 _26324_ (.A1(\cpuregs[9][12] ),
    .A2(_20067_),
    .B1(_20068_),
    .C1(_20070_),
    .X(_20071_));
 sky130_vsdinv _26325_ (.A(\cpuregs[10][12] ),
    .Y(_20072_));
 sky130_fd_sc_hd__nor2_4 _26326_ (.A(_20072_),
    .B(_19359_),
    .Y(_20073_));
 sky130_fd_sc_hd__a211o_4 _26327_ (.A1(\cpuregs[11][12] ),
    .A2(_19630_),
    .B1(_19456_),
    .C1(_20073_),
    .X(_20074_));
 sky130_fd_sc_hd__a21o_4 _26328_ (.A1(_20071_),
    .A2(_20074_),
    .B1(_19473_),
    .X(_20075_));
 sky130_fd_sc_hd__buf_1 _26329_ (.A(_19275_),
    .X(_20076_));
 sky130_fd_sc_hd__nand3_4 _26330_ (.A(_20066_),
    .B(_20075_),
    .C(_20076_),
    .Y(_20077_));
 sky130_fd_sc_hd__buf_1 _26331_ (.A(_19329_),
    .X(_20078_));
 sky130_fd_sc_hd__and2_4 _26332_ (.A(_20077_),
    .B(_20078_),
    .X(_20079_));
 sky130_fd_sc_hd__buf_1 _26333_ (.A(_19268_),
    .X(_20080_));
 sky130_fd_sc_hd__buf_1 _26334_ (.A(_20080_),
    .X(_20081_));
 sky130_fd_sc_hd__buf_1 _26335_ (.A(_19270_),
    .X(_20082_));
 sky130_fd_sc_hd__buf_1 _26336_ (.A(_20082_),
    .X(_20083_));
 sky130_fd_sc_hd__buf_1 _26337_ (.A(_19498_),
    .X(_20084_));
 sky130_fd_sc_hd__and2_4 _26338_ (.A(_20084_),
    .B(\cpuregs[0][12] ),
    .X(_20085_));
 sky130_fd_sc_hd__a211o_4 _26339_ (.A1(\cpuregs[1][12] ),
    .A2(_20081_),
    .B1(_20083_),
    .C1(_20085_),
    .X(_20086_));
 sky130_fd_sc_hd__buf_1 _26340_ (.A(_19594_),
    .X(_20087_));
 sky130_vsdinv _26341_ (.A(\cpuregs[2][12] ),
    .Y(_20088_));
 sky130_fd_sc_hd__buf_1 _26342_ (.A(_19319_),
    .X(_20089_));
 sky130_fd_sc_hd__nor2_4 _26343_ (.A(_20088_),
    .B(_20089_),
    .Y(_20090_));
 sky130_fd_sc_hd__a211o_4 _26344_ (.A1(\cpuregs[3][12] ),
    .A2(_19459_),
    .B1(_20087_),
    .C1(_20090_),
    .X(_20091_));
 sky130_fd_sc_hd__a21o_4 _26345_ (.A1(_20086_),
    .A2(_20091_),
    .B1(_19474_),
    .X(_20092_));
 sky130_fd_sc_hd__buf_1 _26346_ (.A(_19822_),
    .X(_20093_));
 sky130_vsdinv _26347_ (.A(\cpuregs[6][12] ),
    .Y(_20094_));
 sky130_fd_sc_hd__nor2_4 _26348_ (.A(_20094_),
    .B(_19430_),
    .Y(_20095_));
 sky130_fd_sc_hd__a211o_4 _26349_ (.A1(\cpuregs[7][12] ),
    .A2(_20093_),
    .B1(_20035_),
    .C1(_20095_),
    .X(_20096_));
 sky130_vsdinv _26350_ (.A(\cpuregs[4][12] ),
    .Y(_20097_));
 sky130_fd_sc_hd__nor2_4 _26351_ (.A(_20097_),
    .B(_19434_),
    .Y(_20098_));
 sky130_fd_sc_hd__a211o_4 _26352_ (.A1(\cpuregs[5][12] ),
    .A2(_19335_),
    .B1(_19606_),
    .C1(_20098_),
    .X(_20099_));
 sky130_fd_sc_hd__a21o_4 _26353_ (.A1(_20096_),
    .A2(_20099_),
    .B1(_19463_),
    .X(_20100_));
 sky130_fd_sc_hd__nand3_4 _26354_ (.A(_20092_),
    .B(_19477_),
    .C(_20100_),
    .Y(_20101_));
 sky130_fd_sc_hd__buf_1 _26355_ (.A(_19192_),
    .X(_20102_));
 sky130_fd_sc_hd__buf_1 _26356_ (.A(_20102_),
    .X(_20103_));
 sky130_vsdinv _26357_ (.A(\cpuregs[18][12] ),
    .Y(_20104_));
 sky130_fd_sc_hd__nor2_4 _26358_ (.A(_20104_),
    .B(_19558_),
    .Y(_20105_));
 sky130_fd_sc_hd__a211o_4 _26359_ (.A1(\cpuregs[19][12] ),
    .A2(_19199_),
    .B1(_20036_),
    .C1(_20105_),
    .X(_20106_));
 sky130_vsdinv _26360_ (.A(\cpuregs[16][12] ),
    .Y(_20107_));
 sky130_fd_sc_hd__nor2_4 _26361_ (.A(_20107_),
    .B(_19743_),
    .Y(_20108_));
 sky130_fd_sc_hd__a211o_4 _26362_ (.A1(\cpuregs[17][12] ),
    .A2(_19741_),
    .B1(_20042_),
    .C1(_20108_),
    .X(_20109_));
 sky130_fd_sc_hd__a21oi_4 _26363_ (.A1(_20106_),
    .A2(_20109_),
    .B1(_20048_),
    .Y(_20110_));
 sky130_fd_sc_hd__a211o_4 _26364_ (.A1(_20079_),
    .A2(_20101_),
    .B1(_20103_),
    .C1(_20110_),
    .X(_20111_));
 sky130_fd_sc_hd__a21oi_4 _26365_ (.A1(_20111_),
    .A2(_20051_),
    .B1(_18229_),
    .Y(_20112_));
 sky130_fd_sc_hd__o21a_4 _26366_ (.A1(_20053_),
    .A2(_20056_),
    .B1(_20112_),
    .X(_00629_));
 sky130_fd_sc_hd__nand4_4 _26367_ (.A(_19979_),
    .B(_19152_),
    .C(_18908_),
    .D(_20054_),
    .Y(_20113_));
 sky130_fd_sc_hd__o21a_4 _26368_ (.A1(_18908_),
    .A2(_20053_),
    .B1(_20113_),
    .X(_20114_));
 sky130_fd_sc_hd__buf_1 _26369_ (.A(_19570_),
    .X(_20115_));
 sky130_vsdinv _26370_ (.A(\cpuregs[14][13] ),
    .Y(_20116_));
 sky130_fd_sc_hd__nor2_4 _26371_ (.A(_20116_),
    .B(_19985_),
    .Y(_20117_));
 sky130_fd_sc_hd__a211o_4 _26372_ (.A1(\cpuregs[15][13] ),
    .A2(_19983_),
    .B1(_20115_),
    .C1(_20117_),
    .X(_20118_));
 sky130_fd_sc_hd__buf_1 _26373_ (.A(_19587_),
    .X(_20119_));
 sky130_vsdinv _26374_ (.A(\cpuregs[12][13] ),
    .Y(_20120_));
 sky130_fd_sc_hd__nor2_4 _26375_ (.A(_20120_),
    .B(_19990_),
    .Y(_20121_));
 sky130_fd_sc_hd__a211o_4 _26376_ (.A1(\cpuregs[13][13] ),
    .A2(_19988_),
    .B1(_20119_),
    .C1(_20121_),
    .X(_20122_));
 sky130_fd_sc_hd__buf_1 _26377_ (.A(_19583_),
    .X(_20123_));
 sky130_fd_sc_hd__a21o_4 _26378_ (.A1(_20118_),
    .A2(_20122_),
    .B1(_20123_),
    .X(_20124_));
 sky130_vsdinv _26379_ (.A(\cpuregs[8][13] ),
    .Y(_20125_));
 sky130_fd_sc_hd__nor2_4 _26380_ (.A(_20125_),
    .B(_19844_),
    .Y(_20126_));
 sky130_fd_sc_hd__a211o_4 _26381_ (.A1(\cpuregs[9][13] ),
    .A2(_19284_),
    .B1(_19994_),
    .C1(_20126_),
    .X(_20127_));
 sky130_fd_sc_hd__buf_1 _26382_ (.A(_19296_),
    .X(_20128_));
 sky130_vsdinv _26383_ (.A(\cpuregs[10][13] ),
    .Y(_20129_));
 sky130_fd_sc_hd__nor2_4 _26384_ (.A(_20129_),
    .B(_19302_),
    .Y(_20130_));
 sky130_fd_sc_hd__a211o_4 _26385_ (.A1(\cpuregs[11][13] ),
    .A2(_20128_),
    .B1(_19711_),
    .C1(_20130_),
    .X(_20131_));
 sky130_fd_sc_hd__a21o_4 _26386_ (.A1(_20127_),
    .A2(_20131_),
    .B1(_20001_),
    .X(_20132_));
 sky130_fd_sc_hd__nand3_4 _26387_ (.A(_20124_),
    .B(_20132_),
    .C(_19716_),
    .Y(_20133_));
 sky130_fd_sc_hd__and2_4 _26388_ (.A(_20133_),
    .B(_19718_),
    .X(_20134_));
 sky130_fd_sc_hd__and2_4 _26389_ (.A(_20007_),
    .B(\cpuregs[0][13] ),
    .X(_20135_));
 sky130_fd_sc_hd__a211o_4 _26390_ (.A1(\cpuregs[1][13] ),
    .A2(_20005_),
    .B1(_20006_),
    .C1(_20135_),
    .X(_20136_));
 sky130_fd_sc_hd__buf_1 _26391_ (.A(_19573_),
    .X(_20137_));
 sky130_fd_sc_hd__buf_1 _26392_ (.A(_20137_),
    .X(_20138_));
 sky130_vsdinv _26393_ (.A(\cpuregs[2][13] ),
    .Y(_20139_));
 sky130_fd_sc_hd__nor2_4 _26394_ (.A(_20139_),
    .B(_20012_),
    .Y(_20140_));
 sky130_fd_sc_hd__a211o_4 _26395_ (.A1(\cpuregs[3][13] ),
    .A2(_20138_),
    .B1(_20010_),
    .C1(_20140_),
    .X(_20141_));
 sky130_fd_sc_hd__buf_1 _26396_ (.A(_19354_),
    .X(_20142_));
 sky130_fd_sc_hd__a21o_4 _26397_ (.A1(_20136_),
    .A2(_20141_),
    .B1(_20142_),
    .X(_20143_));
 sky130_fd_sc_hd__buf_1 _26398_ (.A(_19357_),
    .X(_20144_));
 sky130_vsdinv _26399_ (.A(\cpuregs[6][13] ),
    .Y(_20145_));
 sky130_fd_sc_hd__nor2_4 _26400_ (.A(_20145_),
    .B(_19440_),
    .Y(_20146_));
 sky130_fd_sc_hd__a211o_4 _26401_ (.A1(\cpuregs[7][13] ),
    .A2(_19773_),
    .B1(_19723_),
    .C1(_20146_),
    .X(_20147_));
 sky130_fd_sc_hd__buf_1 _26402_ (.A(_19541_),
    .X(_20148_));
 sky130_vsdinv _26403_ (.A(\cpuregs[4][13] ),
    .Y(_20149_));
 sky130_fd_sc_hd__buf_1 _26404_ (.A(_19623_),
    .X(_20150_));
 sky130_fd_sc_hd__nor2_4 _26405_ (.A(_20149_),
    .B(_20150_),
    .Y(_20151_));
 sky130_fd_sc_hd__a211o_4 _26406_ (.A1(\cpuregs[5][13] ),
    .A2(_20022_),
    .B1(_20148_),
    .C1(_20151_),
    .X(_20152_));
 sky130_fd_sc_hd__a21o_4 _26407_ (.A1(_20147_),
    .A2(_20152_),
    .B1(_20026_),
    .X(_20153_));
 sky130_fd_sc_hd__nand3_4 _26408_ (.A(_20143_),
    .B(_20144_),
    .C(_20153_),
    .Y(_20154_));
 sky130_fd_sc_hd__buf_1 _26409_ (.A(_19192_),
    .X(_20155_));
 sky130_fd_sc_hd__buf_1 _26410_ (.A(_20155_),
    .X(_20156_));
 sky130_fd_sc_hd__buf_1 _26411_ (.A(_20156_),
    .X(_20157_));
 sky130_fd_sc_hd__buf_1 _26412_ (.A(_19633_),
    .X(_20158_));
 sky130_vsdinv _26413_ (.A(\cpuregs[18][13] ),
    .Y(_20159_));
 sky130_fd_sc_hd__nor2_4 _26414_ (.A(_20159_),
    .B(_20038_),
    .Y(_20160_));
 sky130_fd_sc_hd__a211o_4 _26415_ (.A1(\cpuregs[19][13] ),
    .A2(_20033_),
    .B1(_20158_),
    .C1(_20160_),
    .X(_20161_));
 sky130_fd_sc_hd__buf_1 _26416_ (.A(_19526_),
    .X(_20162_));
 sky130_fd_sc_hd__buf_1 _26417_ (.A(_19527_),
    .X(_20163_));
 sky130_vsdinv _26418_ (.A(\cpuregs[16][13] ),
    .Y(_20164_));
 sky130_fd_sc_hd__buf_1 _26419_ (.A(_20044_),
    .X(_20165_));
 sky130_fd_sc_hd__nor2_4 _26420_ (.A(_20164_),
    .B(_20165_),
    .Y(_20166_));
 sky130_fd_sc_hd__a211o_4 _26421_ (.A1(\cpuregs[17][13] ),
    .A2(_20162_),
    .B1(_20163_),
    .C1(_20166_),
    .X(_20167_));
 sky130_fd_sc_hd__buf_1 _26422_ (.A(_19224_),
    .X(_20168_));
 sky130_fd_sc_hd__a21oi_4 _26423_ (.A1(_20161_),
    .A2(_20167_),
    .B1(_20168_),
    .Y(_20169_));
 sky130_fd_sc_hd__a211o_4 _26424_ (.A1(_20134_),
    .A2(_20154_),
    .B1(_20157_),
    .C1(_20169_),
    .X(_20170_));
 sky130_fd_sc_hd__a21oi_4 _26425_ (.A1(_20170_),
    .A2(_20051_),
    .B1(_18229_),
    .Y(_20171_));
 sky130_fd_sc_hd__o21a_4 _26426_ (.A1(_19932_),
    .A2(_20114_),
    .B1(_20171_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_1 _26427_ (.A(_19417_),
    .X(_20172_));
 sky130_fd_sc_hd__buf_1 _26428_ (.A(_19416_),
    .X(_20173_));
 sky130_fd_sc_hd__buf_1 _26429_ (.A(\timer[15] ),
    .X(_20174_));
 sky130_vsdinv _26430_ (.A(_19157_),
    .Y(_20175_));
 sky130_fd_sc_hd__and4_4 _26431_ (.A(_20055_),
    .B(_19154_),
    .C(_20054_),
    .D(_19159_),
    .X(_20176_));
 sky130_fd_sc_hd__buf_1 _26432_ (.A(_20176_),
    .X(_20177_));
 sky130_fd_sc_hd__o21ai_4 _26433_ (.A1(_20174_),
    .A2(_20175_),
    .B1(_20177_),
    .Y(_20178_));
 sky130_fd_sc_hd__o21ai_4 _26434_ (.A1(_20172_),
    .A2(_20173_),
    .B1(_20178_),
    .Y(_20179_));
 sky130_vsdinv _26435_ (.A(\cpuregs[14][14] ),
    .Y(_20180_));
 sky130_fd_sc_hd__buf_1 _26436_ (.A(_19555_),
    .X(_20181_));
 sky130_fd_sc_hd__nor2_4 _26437_ (.A(_20180_),
    .B(_20181_),
    .Y(_20182_));
 sky130_fd_sc_hd__a211o_4 _26438_ (.A1(\cpuregs[15][14] ),
    .A2(_19983_),
    .B1(_20115_),
    .C1(_20182_),
    .X(_20183_));
 sky130_vsdinv _26439_ (.A(\cpuregs[12][14] ),
    .Y(_20184_));
 sky130_fd_sc_hd__nor2_4 _26440_ (.A(_20184_),
    .B(_19990_),
    .Y(_20185_));
 sky130_fd_sc_hd__a211o_4 _26441_ (.A1(\cpuregs[13][14] ),
    .A2(_19988_),
    .B1(_20119_),
    .C1(_20185_),
    .X(_20186_));
 sky130_fd_sc_hd__a21o_4 _26442_ (.A1(_20183_),
    .A2(_20186_),
    .B1(_20123_),
    .X(_20187_));
 sky130_fd_sc_hd__buf_1 _26443_ (.A(_19318_),
    .X(_20188_));
 sky130_vsdinv _26444_ (.A(\cpuregs[8][14] ),
    .Y(_20189_));
 sky130_fd_sc_hd__nor2_4 _26445_ (.A(_20189_),
    .B(_19844_),
    .Y(_20190_));
 sky130_fd_sc_hd__a211o_4 _26446_ (.A1(\cpuregs[9][14] ),
    .A2(_20188_),
    .B1(_19994_),
    .C1(_20190_),
    .X(_20191_));
 sky130_fd_sc_hd__buf_1 _26447_ (.A(_19286_),
    .X(_20192_));
 sky130_vsdinv _26448_ (.A(\cpuregs[10][14] ),
    .Y(_20193_));
 sky130_fd_sc_hd__buf_1 _26449_ (.A(_19301_),
    .X(_20194_));
 sky130_fd_sc_hd__nor2_4 _26450_ (.A(_20193_),
    .B(_20194_),
    .Y(_20195_));
 sky130_fd_sc_hd__a211o_4 _26451_ (.A1(\cpuregs[11][14] ),
    .A2(_20128_),
    .B1(_20192_),
    .C1(_20195_),
    .X(_20196_));
 sky130_fd_sc_hd__a21o_4 _26452_ (.A1(_20191_),
    .A2(_20196_),
    .B1(_20001_),
    .X(_20197_));
 sky130_fd_sc_hd__buf_1 _26453_ (.A(_19326_),
    .X(_20198_));
 sky130_fd_sc_hd__nand3_4 _26454_ (.A(_20187_),
    .B(_20197_),
    .C(_20198_),
    .Y(_20199_));
 sky130_fd_sc_hd__buf_1 _26455_ (.A(_19223_),
    .X(_20200_));
 sky130_fd_sc_hd__and2_4 _26456_ (.A(_20199_),
    .B(_20200_),
    .X(_20201_));
 sky130_fd_sc_hd__buf_1 _26457_ (.A(_19337_),
    .X(_20202_));
 sky130_fd_sc_hd__and2_4 _26458_ (.A(_20202_),
    .B(\cpuregs[0][14] ),
    .X(_20203_));
 sky130_fd_sc_hd__a211o_4 _26459_ (.A1(\cpuregs[1][14] ),
    .A2(_20005_),
    .B1(_20006_),
    .C1(_20203_),
    .X(_20204_));
 sky130_vsdinv _26460_ (.A(\cpuregs[2][14] ),
    .Y(_20205_));
 sky130_fd_sc_hd__nor2_4 _26461_ (.A(_20205_),
    .B(_20012_),
    .Y(_20206_));
 sky130_fd_sc_hd__a211o_4 _26462_ (.A1(\cpuregs[3][14] ),
    .A2(_20138_),
    .B1(_20010_),
    .C1(_20206_),
    .X(_20207_));
 sky130_fd_sc_hd__a21o_4 _26463_ (.A1(_20204_),
    .A2(_20207_),
    .B1(_20142_),
    .X(_20208_));
 sky130_fd_sc_hd__buf_1 _26464_ (.A(_19531_),
    .X(_20209_));
 sky130_fd_sc_hd__buf_1 _26465_ (.A(_19533_),
    .X(_20210_));
 sky130_vsdinv _26466_ (.A(\cpuregs[6][14] ),
    .Y(_20211_));
 sky130_fd_sc_hd__nor2_4 _26467_ (.A(_20211_),
    .B(_19440_),
    .Y(_20212_));
 sky130_fd_sc_hd__a211o_4 _26468_ (.A1(\cpuregs[7][14] ),
    .A2(_20209_),
    .B1(_20210_),
    .C1(_20212_),
    .X(_20213_));
 sky130_vsdinv _26469_ (.A(\cpuregs[4][14] ),
    .Y(_20214_));
 sky130_fd_sc_hd__nor2_4 _26470_ (.A(_20214_),
    .B(_20150_),
    .Y(_20215_));
 sky130_fd_sc_hd__a211o_4 _26471_ (.A1(\cpuregs[5][14] ),
    .A2(_20022_),
    .B1(_20148_),
    .C1(_20215_),
    .X(_20216_));
 sky130_fd_sc_hd__a21o_4 _26472_ (.A1(_20213_),
    .A2(_20216_),
    .B1(_20026_),
    .X(_20217_));
 sky130_fd_sc_hd__nand3_4 _26473_ (.A(_20208_),
    .B(_20144_),
    .C(_20217_),
    .Y(_20218_));
 sky130_vsdinv _26474_ (.A(\cpuregs[18][14] ),
    .Y(_20219_));
 sky130_fd_sc_hd__nor2_4 _26475_ (.A(_20219_),
    .B(_20038_),
    .Y(_20220_));
 sky130_fd_sc_hd__a211o_4 _26476_ (.A1(\cpuregs[19][14] ),
    .A2(_20033_),
    .B1(_20158_),
    .C1(_20220_),
    .X(_20221_));
 sky130_vsdinv _26477_ (.A(\cpuregs[16][14] ),
    .Y(_20222_));
 sky130_fd_sc_hd__nor2_4 _26478_ (.A(_20222_),
    .B(_20165_),
    .Y(_20223_));
 sky130_fd_sc_hd__a211o_4 _26479_ (.A1(\cpuregs[17][14] ),
    .A2(_20162_),
    .B1(_20163_),
    .C1(_20223_),
    .X(_20224_));
 sky130_fd_sc_hd__a21oi_4 _26480_ (.A1(_20221_),
    .A2(_20224_),
    .B1(_20168_),
    .Y(_20225_));
 sky130_fd_sc_hd__a211o_4 _26481_ (.A1(_20201_),
    .A2(_20218_),
    .B1(_20030_),
    .C1(_20225_),
    .X(_20226_));
 sky130_fd_sc_hd__o21ai_4 _26482_ (.A1(_18512_),
    .A2(_20226_),
    .B1(_19097_),
    .Y(_20227_));
 sky130_fd_sc_hd__a21o_4 _26483_ (.A1(_18512_),
    .A2(_20179_),
    .B1(_20227_),
    .X(_20228_));
 sky130_vsdinv _26484_ (.A(_20173_),
    .Y(_20229_));
 sky130_fd_sc_hd__buf_1 _26485_ (.A(_18797_),
    .X(_20230_));
 sky130_fd_sc_hd__buf_1 _26486_ (.A(_20230_),
    .X(_20231_));
 sky130_fd_sc_hd__buf_1 _26487_ (.A(_20231_),
    .X(_20232_));
 sky130_fd_sc_hd__buf_1 _26488_ (.A(_20176_),
    .X(_20233_));
 sky130_fd_sc_hd__o21a_4 _26489_ (.A1(_20174_),
    .A2(_20175_),
    .B1(_20233_),
    .X(_20234_));
 sky130_fd_sc_hd__a211o_4 _26490_ (.A1(\timer[14] ),
    .A2(_20229_),
    .B1(_20232_),
    .C1(_20234_),
    .X(_20235_));
 sky130_fd_sc_hd__and3_4 _26491_ (.A(_20228_),
    .B(_19034_),
    .C(_20235_),
    .X(_00631_));
 sky130_vsdinv _26492_ (.A(\cpuregs[14][15] ),
    .Y(_20236_));
 sky130_fd_sc_hd__nor2_4 _26493_ (.A(_20236_),
    .B(_20181_),
    .Y(_20237_));
 sky130_fd_sc_hd__a211o_4 _26494_ (.A1(\cpuregs[15][15] ),
    .A2(_19983_),
    .B1(_20115_),
    .C1(_20237_),
    .X(_20238_));
 sky130_vsdinv _26495_ (.A(\cpuregs[12][15] ),
    .Y(_20239_));
 sky130_fd_sc_hd__nor2_4 _26496_ (.A(_20239_),
    .B(_19503_),
    .Y(_20240_));
 sky130_fd_sc_hd__a211o_4 _26497_ (.A1(\cpuregs[13][15] ),
    .A2(_20080_),
    .B1(_20119_),
    .C1(_20240_),
    .X(_20241_));
 sky130_fd_sc_hd__a21o_4 _26498_ (.A1(_20238_),
    .A2(_20241_),
    .B1(_20123_),
    .X(_20242_));
 sky130_vsdinv _26499_ (.A(\cpuregs[8][15] ),
    .Y(_20243_));
 sky130_fd_sc_hd__nor2_4 _26500_ (.A(_20243_),
    .B(_19404_),
    .Y(_20244_));
 sky130_fd_sc_hd__a211o_4 _26501_ (.A1(\cpuregs[9][15] ),
    .A2(_20188_),
    .B1(_19994_),
    .C1(_20244_),
    .X(_20245_));
 sky130_vsdinv _26502_ (.A(\cpuregs[10][15] ),
    .Y(_20246_));
 sky130_fd_sc_hd__nor2_4 _26503_ (.A(_20246_),
    .B(_20194_),
    .Y(_20247_));
 sky130_fd_sc_hd__a211o_4 _26504_ (.A1(\cpuregs[11][15] ),
    .A2(_20128_),
    .B1(_20192_),
    .C1(_20247_),
    .X(_20248_));
 sky130_fd_sc_hd__a21o_4 _26505_ (.A1(_20245_),
    .A2(_20248_),
    .B1(_20001_),
    .X(_20249_));
 sky130_fd_sc_hd__nand3_4 _26506_ (.A(_20242_),
    .B(_20249_),
    .C(_20198_),
    .Y(_20250_));
 sky130_fd_sc_hd__and2_4 _26507_ (.A(_20250_),
    .B(_20200_),
    .X(_20251_));
 sky130_fd_sc_hd__and2_4 _26508_ (.A(_20202_),
    .B(\cpuregs[0][15] ),
    .X(_20252_));
 sky130_fd_sc_hd__a211o_4 _26509_ (.A1(\cpuregs[1][15] ),
    .A2(_19631_),
    .B1(_19336_),
    .C1(_20252_),
    .X(_20253_));
 sky130_vsdinv _26510_ (.A(\cpuregs[2][15] ),
    .Y(_20254_));
 sky130_fd_sc_hd__nor2_4 _26511_ (.A(_20254_),
    .B(_20012_),
    .Y(_20255_));
 sky130_fd_sc_hd__a211o_4 _26512_ (.A1(\cpuregs[3][15] ),
    .A2(_20138_),
    .B1(_20010_),
    .C1(_20255_),
    .X(_20256_));
 sky130_fd_sc_hd__a21o_4 _26513_ (.A1(_20253_),
    .A2(_20256_),
    .B1(_20142_),
    .X(_20257_));
 sky130_vsdinv _26514_ (.A(\cpuregs[6][15] ),
    .Y(_20258_));
 sky130_fd_sc_hd__buf_1 _26515_ (.A(_19515_),
    .X(_20259_));
 sky130_fd_sc_hd__nor2_4 _26516_ (.A(_20258_),
    .B(_20259_),
    .Y(_20260_));
 sky130_fd_sc_hd__a211o_4 _26517_ (.A1(\cpuregs[7][15] ),
    .A2(_20209_),
    .B1(_20210_),
    .C1(_20260_),
    .X(_20261_));
 sky130_vsdinv _26518_ (.A(\cpuregs[4][15] ),
    .Y(_20262_));
 sky130_fd_sc_hd__nor2_4 _26519_ (.A(_20262_),
    .B(_20150_),
    .Y(_20263_));
 sky130_fd_sc_hd__a211o_4 _26520_ (.A1(\cpuregs[5][15] ),
    .A2(_20022_),
    .B1(_20148_),
    .C1(_20263_),
    .X(_20264_));
 sky130_fd_sc_hd__a21o_4 _26521_ (.A1(_20261_),
    .A2(_20264_),
    .B1(_20026_),
    .X(_20265_));
 sky130_fd_sc_hd__nand3_4 _26522_ (.A(_20257_),
    .B(_20144_),
    .C(_20265_),
    .Y(_20266_));
 sky130_fd_sc_hd__buf_1 _26523_ (.A(_19193_),
    .X(_20267_));
 sky130_vsdinv _26524_ (.A(\cpuregs[18][15] ),
    .Y(_20268_));
 sky130_fd_sc_hd__nor2_4 _26525_ (.A(_20268_),
    .B(_20038_),
    .Y(_20269_));
 sky130_fd_sc_hd__a211o_4 _26526_ (.A1(\cpuregs[19][15] ),
    .A2(_20033_),
    .B1(_20158_),
    .C1(_20269_),
    .X(_20270_));
 sky130_vsdinv _26527_ (.A(\cpuregs[16][15] ),
    .Y(_20271_));
 sky130_fd_sc_hd__nor2_4 _26528_ (.A(_20271_),
    .B(_20165_),
    .Y(_20272_));
 sky130_fd_sc_hd__a211o_4 _26529_ (.A1(\cpuregs[17][15] ),
    .A2(_20162_),
    .B1(_20163_),
    .C1(_20272_),
    .X(_20273_));
 sky130_fd_sc_hd__a21oi_4 _26530_ (.A1(_20270_),
    .A2(_20273_),
    .B1(_20168_),
    .Y(_20274_));
 sky130_fd_sc_hd__a211o_4 _26531_ (.A1(_20251_),
    .A2(_20266_),
    .B1(_20267_),
    .C1(_20274_),
    .X(_20275_));
 sky130_fd_sc_hd__nand2_4 _26532_ (.A(_20275_),
    .B(_19976_),
    .Y(_20276_));
 sky130_vsdinv _26533_ (.A(_20233_),
    .Y(_20277_));
 sky130_fd_sc_hd__and3_4 _26534_ (.A(_20177_),
    .B(_19415_),
    .C(_20175_),
    .X(_20278_));
 sky130_fd_sc_hd__a211o_4 _26535_ (.A1(_20174_),
    .A2(_20277_),
    .B1(_19931_),
    .C1(_20278_),
    .X(_20279_));
 sky130_fd_sc_hd__nand3_4 _26536_ (.A(_20276_),
    .B(_20279_),
    .C(_18843_),
    .Y(_20280_));
 sky130_vsdinv _26537_ (.A(_20280_),
    .Y(_00632_));
 sky130_vsdinv _26538_ (.A(\cpuregs[14][16] ),
    .Y(_20281_));
 sky130_fd_sc_hd__nor2_4 _26539_ (.A(_20281_),
    .B(_19807_),
    .Y(_20282_));
 sky130_fd_sc_hd__a211o_4 _26540_ (.A1(\cpuregs[15][16] ),
    .A2(_19804_),
    .B1(_19805_),
    .C1(_20282_),
    .X(_20283_));
 sky130_vsdinv _26541_ (.A(\cpuregs[12][16] ),
    .Y(_20284_));
 sky130_fd_sc_hd__nor2_4 _26542_ (.A(_20284_),
    .B(_19812_),
    .Y(_20285_));
 sky130_fd_sc_hd__a211o_4 _26543_ (.A1(\cpuregs[13][16] ),
    .A2(_19761_),
    .B1(_19810_),
    .C1(_20285_),
    .X(_20286_));
 sky130_fd_sc_hd__a21o_4 _26544_ (.A1(_20283_),
    .A2(_20286_),
    .B1(_19815_),
    .X(_20287_));
 sky130_vsdinv _26545_ (.A(\cpuregs[8][16] ),
    .Y(_20288_));
 sky130_fd_sc_hd__nor2_4 _26546_ (.A(_20288_),
    .B(_19878_),
    .Y(_20289_));
 sky130_fd_sc_hd__a211o_4 _26547_ (.A1(\cpuregs[9][16] ),
    .A2(_19817_),
    .B1(_19876_),
    .C1(_20289_),
    .X(_20290_));
 sky130_fd_sc_hd__buf_1 _26548_ (.A(_19333_),
    .X(_20291_));
 sky130_vsdinv _26549_ (.A(\cpuregs[10][16] ),
    .Y(_20292_));
 sky130_fd_sc_hd__nor2_4 _26550_ (.A(_20292_),
    .B(_19882_),
    .Y(_20293_));
 sky130_fd_sc_hd__a211o_4 _26551_ (.A1(\cpuregs[11][16] ),
    .A2(_20291_),
    .B1(_19513_),
    .C1(_20293_),
    .X(_20294_));
 sky130_fd_sc_hd__a21o_4 _26552_ (.A1(_20290_),
    .A2(_20294_),
    .B1(_19826_),
    .X(_20295_));
 sky130_fd_sc_hd__nand3_4 _26553_ (.A(_20287_),
    .B(_20295_),
    .C(_19520_),
    .Y(_20296_));
 sky130_fd_sc_hd__and2_4 _26554_ (.A(_20296_),
    .B(_19887_),
    .X(_20297_));
 sky130_fd_sc_hd__buf_1 _26555_ (.A(_19342_),
    .X(_20298_));
 sky130_fd_sc_hd__and2_4 _26556_ (.A(_19889_),
    .B(\cpuregs[0][16] ),
    .X(_20299_));
 sky130_fd_sc_hd__a211o_4 _26557_ (.A1(\cpuregs[1][16] ),
    .A2(_20298_),
    .B1(_19831_),
    .C1(_20299_),
    .X(_20300_));
 sky130_fd_sc_hd__buf_1 _26558_ (.A(_19183_),
    .X(_20301_));
 sky130_vsdinv _26559_ (.A(\cpuregs[2][16] ),
    .Y(_20302_));
 sky130_fd_sc_hd__buf_1 _26560_ (.A(_19730_),
    .X(_20303_));
 sky130_fd_sc_hd__nor2_4 _26561_ (.A(_20302_),
    .B(_20303_),
    .Y(_20304_));
 sky130_fd_sc_hd__a211o_4 _26562_ (.A1(\cpuregs[3][16] ),
    .A2(_19893_),
    .B1(_20301_),
    .C1(_20304_),
    .X(_20305_));
 sky130_fd_sc_hd__a21o_4 _26563_ (.A1(_20300_),
    .A2(_20305_),
    .B1(_19897_),
    .X(_20306_));
 sky130_fd_sc_hd__buf_1 _26564_ (.A(_19183_),
    .X(_20307_));
 sky130_vsdinv _26565_ (.A(\cpuregs[6][16] ),
    .Y(_20308_));
 sky130_fd_sc_hd__buf_1 _26566_ (.A(_19623_),
    .X(_20309_));
 sky130_fd_sc_hd__nor2_4 _26567_ (.A(_20308_),
    .B(_20309_),
    .Y(_20310_));
 sky130_fd_sc_hd__a211o_4 _26568_ (.A1(\cpuregs[7][16] ),
    .A2(_19899_),
    .B1(_20307_),
    .C1(_20310_),
    .X(_20311_));
 sky130_vsdinv _26569_ (.A(\cpuregs[4][16] ),
    .Y(_20312_));
 sky130_fd_sc_hd__buf_1 _26570_ (.A(_19228_),
    .X(_20313_));
 sky130_fd_sc_hd__nor2_4 _26571_ (.A(_20312_),
    .B(_20313_),
    .Y(_20314_));
 sky130_fd_sc_hd__a211o_4 _26572_ (.A1(\cpuregs[5][16] ),
    .A2(_19845_),
    .B1(_19846_),
    .C1(_20314_),
    .X(_20315_));
 sky130_fd_sc_hd__a21o_4 _26573_ (.A1(_20311_),
    .A2(_20315_),
    .B1(_19851_),
    .X(_20316_));
 sky130_fd_sc_hd__nand3_4 _26574_ (.A(_20306_),
    .B(_19838_),
    .C(_20316_),
    .Y(_20317_));
 sky130_fd_sc_hd__buf_1 _26575_ (.A(_19164_),
    .X(_20318_));
 sky130_vsdinv _26576_ (.A(\cpuregs[18][16] ),
    .Y(_20319_));
 sky130_fd_sc_hd__nor2_4 _26577_ (.A(_20319_),
    .B(_19856_),
    .Y(_20320_));
 sky130_fd_sc_hd__a211o_4 _26578_ (.A1(\cpuregs[19][16] ),
    .A2(_19854_),
    .B1(_19908_),
    .C1(_20320_),
    .X(_20321_));
 sky130_vsdinv _26579_ (.A(\cpuregs[16][16] ),
    .Y(_20322_));
 sky130_fd_sc_hd__nor2_4 _26580_ (.A(_20322_),
    .B(_19915_),
    .Y(_20323_));
 sky130_fd_sc_hd__a211o_4 _26581_ (.A1(\cpuregs[17][16] ),
    .A2(_19912_),
    .B1(_19913_),
    .C1(_20323_),
    .X(_20324_));
 sky130_fd_sc_hd__a21oi_4 _26582_ (.A1(_20321_),
    .A2(_20324_),
    .B1(_19918_),
    .Y(_20325_));
 sky130_fd_sc_hd__a2111o_4 _26583_ (.A1(_20297_),
    .A2(_20317_),
    .B1(_20318_),
    .C1(_19786_),
    .D1(_20325_),
    .X(_20326_));
 sky130_fd_sc_hd__and4_4 _26584_ (.A(_19864_),
    .B(_19979_),
    .C(_20054_),
    .D(_18910_),
    .X(_20327_));
 sky130_fd_sc_hd__buf_1 _26585_ (.A(\timer[16] ),
    .X(_20328_));
 sky130_fd_sc_hd__a41o_4 _26586_ (.A1(_20327_),
    .A2(_19154_),
    .A3(_19925_),
    .A4(_20172_),
    .B1(_20328_),
    .X(_20329_));
 sky130_fd_sc_hd__buf_1 _26587_ (.A(_19925_),
    .X(_20330_));
 sky130_fd_sc_hd__nand4_4 _26588_ (.A(_20330_),
    .B(_20173_),
    .C(_20172_),
    .D(_20328_),
    .Y(_20331_));
 sky130_fd_sc_hd__nand3_4 _26589_ (.A(_19421_),
    .B(_20329_),
    .C(_20331_),
    .Y(_20332_));
 sky130_fd_sc_hd__buf_1 _26590_ (.A(_19495_),
    .X(_20333_));
 sky130_fd_sc_hd__a21oi_4 _26591_ (.A1(_20326_),
    .A2(_20332_),
    .B1(_20333_),
    .Y(_00633_));
 sky130_fd_sc_hd__buf_1 _26592_ (.A(_19268_),
    .X(_20334_));
 sky130_vsdinv _26593_ (.A(\cpuregs[14][17] ),
    .Y(_20335_));
 sky130_fd_sc_hd__nor2_4 _26594_ (.A(_20335_),
    .B(_19936_),
    .Y(_20336_));
 sky130_fd_sc_hd__a211o_4 _26595_ (.A1(\cpuregs[15][17] ),
    .A2(_20334_),
    .B1(_20058_),
    .C1(_20336_),
    .X(_20337_));
 sky130_fd_sc_hd__buf_1 _26596_ (.A(_19270_),
    .X(_20338_));
 sky130_vsdinv _26597_ (.A(\cpuregs[12][17] ),
    .Y(_20339_));
 sky130_fd_sc_hd__nor2_4 _26598_ (.A(_20339_),
    .B(_20137_),
    .Y(_20340_));
 sky130_fd_sc_hd__a211o_4 _26599_ (.A1(\cpuregs[13][17] ),
    .A2(_19445_),
    .B1(_20338_),
    .C1(_20340_),
    .X(_20341_));
 sky130_fd_sc_hd__a21o_4 _26600_ (.A1(_20337_),
    .A2(_20341_),
    .B1(_20065_),
    .X(_20342_));
 sky130_vsdinv _26601_ (.A(\cpuregs[8][17] ),
    .Y(_20343_));
 sky130_fd_sc_hd__nor2_4 _26602_ (.A(_20343_),
    .B(_19985_),
    .Y(_20344_));
 sky130_fd_sc_hd__a211o_4 _26603_ (.A1(\cpuregs[9][17] ),
    .A2(_20067_),
    .B1(_20068_),
    .C1(_20344_),
    .X(_20345_));
 sky130_vsdinv _26604_ (.A(\cpuregs[10][17] ),
    .Y(_20346_));
 sky130_fd_sc_hd__nor2_4 _26605_ (.A(_20346_),
    .B(_19394_),
    .Y(_20347_));
 sky130_fd_sc_hd__a211o_4 _26606_ (.A1(\cpuregs[11][17] ),
    .A2(_19630_),
    .B1(_19456_),
    .C1(_20347_),
    .X(_20348_));
 sky130_fd_sc_hd__a21o_4 _26607_ (.A1(_20345_),
    .A2(_20348_),
    .B1(_20015_),
    .X(_20349_));
 sky130_fd_sc_hd__nand3_4 _26608_ (.A(_20342_),
    .B(_20349_),
    .C(_20076_),
    .Y(_20350_));
 sky130_fd_sc_hd__and2_4 _26609_ (.A(_20350_),
    .B(_20078_),
    .X(_20351_));
 sky130_fd_sc_hd__and2_4 _26610_ (.A(_20084_),
    .B(\cpuregs[0][17] ),
    .X(_20352_));
 sky130_fd_sc_hd__a211o_4 _26611_ (.A1(\cpuregs[1][17] ),
    .A2(_19459_),
    .B1(_20083_),
    .C1(_20352_),
    .X(_20353_));
 sky130_vsdinv _26612_ (.A(\cpuregs[2][17] ),
    .Y(_20354_));
 sky130_fd_sc_hd__nor2_4 _26613_ (.A(_20354_),
    .B(_19969_),
    .Y(_20355_));
 sky130_fd_sc_hd__a211o_4 _26614_ (.A1(\cpuregs[3][17] ),
    .A2(_19198_),
    .B1(_19202_),
    .C1(_20355_),
    .X(_20356_));
 sky130_fd_sc_hd__a21o_4 _26615_ (.A1(_20353_),
    .A2(_20356_),
    .B1(_20016_),
    .X(_20357_));
 sky130_vsdinv _26616_ (.A(\cpuregs[6][17] ),
    .Y(_20358_));
 sky130_fd_sc_hd__nor2_4 _26617_ (.A(_20358_),
    .B(_19395_),
    .Y(_20359_));
 sky130_fd_sc_hd__a211o_4 _26618_ (.A1(\cpuregs[7][17] ),
    .A2(_20032_),
    .B1(_20035_),
    .C1(_20359_),
    .X(_20360_));
 sky130_vsdinv _26619_ (.A(\cpuregs[4][17] ),
    .Y(_20361_));
 sky130_fd_sc_hd__nor2_4 _26620_ (.A(_20361_),
    .B(_19405_),
    .Y(_20362_));
 sky130_fd_sc_hd__a211o_4 _26621_ (.A1(\cpuregs[5][17] ),
    .A2(_19740_),
    .B1(_19720_),
    .C1(_20362_),
    .X(_20363_));
 sky130_fd_sc_hd__a21o_4 _26622_ (.A1(_20360_),
    .A2(_20363_),
    .B1(_19539_),
    .X(_20364_));
 sky130_fd_sc_hd__nand3_4 _26623_ (.A(_20357_),
    .B(_20018_),
    .C(_20364_),
    .Y(_20365_));
 sky130_vsdinv _26624_ (.A(\cpuregs[18][17] ),
    .Y(_20366_));
 sky130_fd_sc_hd__buf_1 _26625_ (.A(_19360_),
    .X(_20367_));
 sky130_fd_sc_hd__nor2_4 _26626_ (.A(_20366_),
    .B(_20367_),
    .Y(_20368_));
 sky130_fd_sc_hd__a211o_4 _26627_ (.A1(\cpuregs[19][17] ),
    .A2(_19210_),
    .B1(_20036_),
    .C1(_20368_),
    .X(_20369_));
 sky130_vsdinv _26628_ (.A(\cpuregs[16][17] ),
    .Y(_20370_));
 sky130_fd_sc_hd__nor2_4 _26629_ (.A(_20370_),
    .B(_19743_),
    .Y(_20371_));
 sky130_fd_sc_hd__a211o_4 _26630_ (.A1(\cpuregs[17][17] ),
    .A2(_19741_),
    .B1(_20042_),
    .C1(_20371_),
    .X(_20372_));
 sky130_fd_sc_hd__a21oi_4 _26631_ (.A1(_20369_),
    .A2(_20372_),
    .B1(_20048_),
    .Y(_20373_));
 sky130_fd_sc_hd__a211o_4 _26632_ (.A1(_20351_),
    .A2(_20365_),
    .B1(_20031_),
    .C1(_20373_),
    .X(_20374_));
 sky130_fd_sc_hd__nand2_4 _26633_ (.A(_20374_),
    .B(_20051_),
    .Y(_20375_));
 sky130_vsdinv _26634_ (.A(_20328_),
    .Y(_20376_));
 sky130_fd_sc_hd__buf_1 _26635_ (.A(_20376_),
    .X(_20377_));
 sky130_fd_sc_hd__and4_4 _26636_ (.A(_20327_),
    .B(_19154_),
    .C(_19414_),
    .D(_19159_),
    .X(_20378_));
 sky130_fd_sc_hd__buf_1 _26637_ (.A(_20378_),
    .X(_20379_));
 sky130_fd_sc_hd__o21ai_4 _26638_ (.A1(_20377_),
    .A2(_19926_),
    .B1(_20379_),
    .Y(_20380_));
 sky130_fd_sc_hd__buf_1 _26639_ (.A(_19418_),
    .X(_20381_));
 sky130_vsdinv _26640_ (.A(\timer[17] ),
    .Y(_20382_));
 sky130_fd_sc_hd__buf_1 _26641_ (.A(_20382_),
    .X(_20383_));
 sky130_fd_sc_hd__nand4_4 _26642_ (.A(_19415_),
    .B(_20177_),
    .C(_20383_),
    .D(_20377_),
    .Y(_20384_));
 sky130_fd_sc_hd__nor2_4 _26643_ (.A(_19926_),
    .B(_20384_),
    .Y(_20385_));
 sky130_fd_sc_hd__a211o_4 _26644_ (.A1(\timer[17] ),
    .A2(_20380_),
    .B1(_20381_),
    .C1(_20385_),
    .X(_20386_));
 sky130_fd_sc_hd__and3_4 _26645_ (.A(_20375_),
    .B(_19034_),
    .C(_20386_),
    .X(_00634_));
 sky130_fd_sc_hd__buf_1 _26646_ (.A(\timer[18] ),
    .X(_20387_));
 sky130_fd_sc_hd__buf_1 _26647_ (.A(_20378_),
    .X(_20388_));
 sky130_fd_sc_hd__nand4_4 _26648_ (.A(_20383_),
    .B(_20388_),
    .C(_20377_),
    .D(_20387_),
    .Y(_20389_));
 sky130_fd_sc_hd__o21a_4 _26649_ (.A1(_20387_),
    .A2(_20385_),
    .B1(_20389_),
    .X(_20390_));
 sky130_vsdinv _26650_ (.A(\cpuregs[14][18] ),
    .Y(_20391_));
 sky130_fd_sc_hd__nor2_4 _26651_ (.A(_20391_),
    .B(_20181_),
    .Y(_20392_));
 sky130_fd_sc_hd__a211o_4 _26652_ (.A1(\cpuregs[15][18] ),
    .A2(_19497_),
    .B1(_20115_),
    .C1(_20392_),
    .X(_20393_));
 sky130_vsdinv _26653_ (.A(\cpuregs[12][18] ),
    .Y(_20394_));
 sky130_fd_sc_hd__nor2_4 _26654_ (.A(_20394_),
    .B(_19503_),
    .Y(_20395_));
 sky130_fd_sc_hd__a211o_4 _26655_ (.A1(\cpuregs[13][18] ),
    .A2(_20080_),
    .B1(_20119_),
    .C1(_20395_),
    .X(_20396_));
 sky130_fd_sc_hd__a21o_4 _26656_ (.A1(_20393_),
    .A2(_20396_),
    .B1(_20123_),
    .X(_20397_));
 sky130_vsdinv _26657_ (.A(\cpuregs[8][18] ),
    .Y(_20398_));
 sky130_fd_sc_hd__nor2_4 _26658_ (.A(_20398_),
    .B(_19404_),
    .Y(_20399_));
 sky130_fd_sc_hd__a211o_4 _26659_ (.A1(\cpuregs[9][18] ),
    .A2(_20188_),
    .B1(_19508_),
    .C1(_20399_),
    .X(_20400_));
 sky130_vsdinv _26660_ (.A(\cpuregs[10][18] ),
    .Y(_20401_));
 sky130_fd_sc_hd__nor2_4 _26661_ (.A(_20401_),
    .B(_20194_),
    .Y(_20402_));
 sky130_fd_sc_hd__a211o_4 _26662_ (.A1(\cpuregs[11][18] ),
    .A2(_20128_),
    .B1(_20192_),
    .C1(_20402_),
    .X(_20403_));
 sky130_fd_sc_hd__a21o_4 _26663_ (.A1(_20400_),
    .A2(_20403_),
    .B1(_19518_),
    .X(_20404_));
 sky130_fd_sc_hd__nand3_4 _26664_ (.A(_20397_),
    .B(_20404_),
    .C(_20198_),
    .Y(_20405_));
 sky130_fd_sc_hd__and2_4 _26665_ (.A(_20405_),
    .B(_20200_),
    .X(_20406_));
 sky130_fd_sc_hd__and2_4 _26666_ (.A(_20202_),
    .B(\cpuregs[0][18] ),
    .X(_20407_));
 sky130_fd_sc_hd__a211o_4 _26667_ (.A1(\cpuregs[1][18] ),
    .A2(_19631_),
    .B1(_19336_),
    .C1(_20407_),
    .X(_20408_));
 sky130_vsdinv _26668_ (.A(\cpuregs[2][18] ),
    .Y(_20409_));
 sky130_fd_sc_hd__nor2_4 _26669_ (.A(_20409_),
    .B(_19350_),
    .Y(_20410_));
 sky130_fd_sc_hd__a211o_4 _26670_ (.A1(\cpuregs[3][18] ),
    .A2(_20138_),
    .B1(_19787_),
    .C1(_20410_),
    .X(_20411_));
 sky130_fd_sc_hd__a21o_4 _26671_ (.A1(_20408_),
    .A2(_20411_),
    .B1(_20142_),
    .X(_20412_));
 sky130_vsdinv _26672_ (.A(\cpuregs[6][18] ),
    .Y(_20413_));
 sky130_fd_sc_hd__nor2_4 _26673_ (.A(_20413_),
    .B(_20259_),
    .Y(_20414_));
 sky130_fd_sc_hd__a211o_4 _26674_ (.A1(\cpuregs[7][18] ),
    .A2(_20209_),
    .B1(_20210_),
    .C1(_20414_),
    .X(_20415_));
 sky130_vsdinv _26675_ (.A(\cpuregs[4][18] ),
    .Y(_20416_));
 sky130_fd_sc_hd__nor2_4 _26676_ (.A(_20416_),
    .B(_20150_),
    .Y(_20417_));
 sky130_fd_sc_hd__a211o_4 _26677_ (.A1(\cpuregs[5][18] ),
    .A2(_19839_),
    .B1(_20148_),
    .C1(_20417_),
    .X(_20418_));
 sky130_fd_sc_hd__a21o_4 _26678_ (.A1(_20415_),
    .A2(_20418_),
    .B1(_19627_),
    .X(_20419_));
 sky130_fd_sc_hd__nand3_4 _26679_ (.A(_20412_),
    .B(_20144_),
    .C(_20419_),
    .Y(_20420_));
 sky130_vsdinv _26680_ (.A(\cpuregs[18][18] ),
    .Y(_20421_));
 sky130_fd_sc_hd__nor2_4 _26681_ (.A(_20421_),
    .B(_19636_),
    .Y(_20422_));
 sky130_fd_sc_hd__a211o_4 _26682_ (.A1(\cpuregs[19][18] ),
    .A2(_19632_),
    .B1(_20158_),
    .C1(_20422_),
    .X(_20423_));
 sky130_vsdinv _26683_ (.A(\cpuregs[16][18] ),
    .Y(_20424_));
 sky130_fd_sc_hd__nor2_4 _26684_ (.A(_20424_),
    .B(_20165_),
    .Y(_20425_));
 sky130_fd_sc_hd__a211o_4 _26685_ (.A1(\cpuregs[17][18] ),
    .A2(_20162_),
    .B1(_20163_),
    .C1(_20425_),
    .X(_20426_));
 sky130_fd_sc_hd__a21oi_4 _26686_ (.A1(_20423_),
    .A2(_20426_),
    .B1(_20168_),
    .Y(_20427_));
 sky130_fd_sc_hd__a211o_4 _26687_ (.A1(_20406_),
    .A2(_20420_),
    .B1(_20157_),
    .C1(_20427_),
    .X(_20428_));
 sky130_fd_sc_hd__buf_1 _26688_ (.A(_19931_),
    .X(_20429_));
 sky130_fd_sc_hd__buf_1 _26689_ (.A(_18228_),
    .X(_20430_));
 sky130_fd_sc_hd__a21oi_4 _26690_ (.A1(_20428_),
    .A2(_20429_),
    .B1(_20430_),
    .Y(_20431_));
 sky130_fd_sc_hd__o21a_4 _26691_ (.A1(_19932_),
    .A2(_20390_),
    .B1(_20431_),
    .X(_00635_));
 sky130_fd_sc_hd__and4_4 _26692_ (.A(_20176_),
    .B(_19414_),
    .C(_20382_),
    .D(_20376_),
    .X(_20432_));
 sky130_fd_sc_hd__buf_1 _26693_ (.A(_20432_),
    .X(_20433_));
 sky130_fd_sc_hd__nor2_4 _26694_ (.A(\timer[19] ),
    .B(_20387_),
    .Y(_20434_));
 sky130_fd_sc_hd__buf_1 _26695_ (.A(_20434_),
    .X(_20435_));
 sky130_fd_sc_hd__and3_4 _26696_ (.A(_20433_),
    .B(_20175_),
    .C(_20435_),
    .X(_20436_));
 sky130_fd_sc_hd__o21ai_4 _26697_ (.A1(_18923_),
    .A2(_19926_),
    .B1(_20388_),
    .Y(_20437_));
 sky130_fd_sc_hd__a21o_4 _26698_ (.A1(_20437_),
    .A2(\timer[19] ),
    .B1(_20381_),
    .X(_20438_));
 sky130_vsdinv _26699_ (.A(\cpuregs[14][19] ),
    .Y(_20439_));
 sky130_fd_sc_hd__nor2_4 _26700_ (.A(_20439_),
    .B(_19512_),
    .Y(_20440_));
 sky130_fd_sc_hd__a211o_4 _26701_ (.A1(\cpuregs[15][19] ),
    .A2(_20057_),
    .B1(_19243_),
    .C1(_20440_),
    .X(_20441_));
 sky130_vsdinv _26702_ (.A(\cpuregs[12][19] ),
    .Y(_20442_));
 sky130_fd_sc_hd__nor2_4 _26703_ (.A(_20442_),
    .B(_19525_),
    .Y(_20443_));
 sky130_fd_sc_hd__a211o_4 _26704_ (.A1(\cpuregs[13][19] ),
    .A2(_20334_),
    .B1(_19271_),
    .C1(_20443_),
    .X(_20444_));
 sky130_fd_sc_hd__a21o_4 _26705_ (.A1(_20441_),
    .A2(_20444_),
    .B1(_19252_),
    .X(_20445_));
 sky130_fd_sc_hd__buf_1 _26706_ (.A(_19196_),
    .X(_20446_));
 sky130_vsdinv _26707_ (.A(\cpuregs[8][19] ),
    .Y(_20447_));
 sky130_fd_sc_hd__nor2_4 _26708_ (.A(_20447_),
    .B(_19609_),
    .Y(_20448_));
 sky130_fd_sc_hd__a211o_4 _26709_ (.A1(\cpuregs[9][19] ),
    .A2(_20446_),
    .B1(_20338_),
    .C1(_20448_),
    .X(_20449_));
 sky130_fd_sc_hd__buf_1 _26710_ (.A(_19570_),
    .X(_20450_));
 sky130_vsdinv _26711_ (.A(\cpuregs[10][19] ),
    .Y(_20451_));
 sky130_fd_sc_hd__nor2_4 _26712_ (.A(_20451_),
    .B(_19892_),
    .Y(_20452_));
 sky130_fd_sc_hd__a211o_4 _26713_ (.A1(\cpuregs[11][19] ),
    .A2(_19481_),
    .B1(_20450_),
    .C1(_20452_),
    .X(_20453_));
 sky130_fd_sc_hd__a21o_4 _26714_ (.A1(_20449_),
    .A2(_20453_),
    .B1(_19473_),
    .X(_20454_));
 sky130_fd_sc_hd__nand3_4 _26715_ (.A(_20445_),
    .B(_20454_),
    .C(_19276_),
    .Y(_20455_));
 sky130_fd_sc_hd__and2_4 _26716_ (.A(_20455_),
    .B(_19279_),
    .X(_20456_));
 sky130_fd_sc_hd__and2_4 _26717_ (.A(_20084_),
    .B(\cpuregs[0][19] ),
    .X(_20457_));
 sky130_fd_sc_hd__a211o_4 _26718_ (.A1(\cpuregs[1][19] ),
    .A2(_19482_),
    .B1(_19452_),
    .C1(_20457_),
    .X(_20458_));
 sky130_vsdinv _26719_ (.A(\cpuregs[2][19] ),
    .Y(_20459_));
 sky130_fd_sc_hd__nor2_4 _26720_ (.A(_20459_),
    .B(_19400_),
    .Y(_20460_));
 sky130_fd_sc_hd__a211o_4 _26721_ (.A1(\cpuregs[3][19] ),
    .A2(_20081_),
    .B1(_19457_),
    .C1(_20460_),
    .X(_20461_));
 sky130_fd_sc_hd__a21o_4 _26722_ (.A1(_20458_),
    .A2(_20461_),
    .B1(_19474_),
    .X(_20462_));
 sky130_vsdinv _26723_ (.A(\cpuregs[6][19] ),
    .Y(_20463_));
 sky130_fd_sc_hd__nor2_4 _26724_ (.A(_20463_),
    .B(_20044_),
    .Y(_20464_));
 sky130_fd_sc_hd__a211o_4 _26725_ (.A1(\cpuregs[7][19] ),
    .A2(_19469_),
    .B1(_20087_),
    .C1(_20464_),
    .X(_20465_));
 sky130_vsdinv _26726_ (.A(\cpuregs[4][19] ),
    .Y(_20466_));
 sky130_fd_sc_hd__nor2_4 _26727_ (.A(_20466_),
    .B(_19430_),
    .Y(_20467_));
 sky130_fd_sc_hd__a211o_4 _26728_ (.A1(\cpuregs[5][19] ),
    .A2(_20093_),
    .B1(_19215_),
    .C1(_20467_),
    .X(_20468_));
 sky130_fd_sc_hd__a21o_4 _26729_ (.A1(_20465_),
    .A2(_20468_),
    .B1(_19463_),
    .X(_20469_));
 sky130_fd_sc_hd__nand3_4 _26730_ (.A(_20462_),
    .B(_19477_),
    .C(_20469_),
    .Y(_20470_));
 sky130_vsdinv _26731_ (.A(\cpuregs[18][19] ),
    .Y(_20471_));
 sky130_fd_sc_hd__nor2_4 _26732_ (.A(_20471_),
    .B(_19558_),
    .Y(_20472_));
 sky130_fd_sc_hd__a211o_4 _26733_ (.A1(\cpuregs[19][19] ),
    .A2(_19199_),
    .B1(_19203_),
    .C1(_20472_),
    .X(_20473_));
 sky130_vsdinv _26734_ (.A(\cpuregs[16][19] ),
    .Y(_20474_));
 sky130_fd_sc_hd__nor2_4 _26735_ (.A(_20474_),
    .B(_20367_),
    .Y(_20475_));
 sky130_fd_sc_hd__a211o_4 _26736_ (.A1(\cpuregs[17][19] ),
    .A2(_19210_),
    .B1(_19216_),
    .C1(_20475_),
    .X(_20476_));
 sky130_fd_sc_hd__a21oi_4 _26737_ (.A1(_20473_),
    .A2(_20476_),
    .B1(_19225_),
    .Y(_20477_));
 sky130_fd_sc_hd__a211o_4 _26738_ (.A1(_20456_),
    .A2(_20470_),
    .B1(_20030_),
    .C1(_20477_),
    .X(_20478_));
 sky130_fd_sc_hd__a21oi_4 _26739_ (.A1(_20478_),
    .A2(_20429_),
    .B1(_20430_),
    .Y(_20479_));
 sky130_fd_sc_hd__o21a_4 _26740_ (.A1(_20436_),
    .A2(_20438_),
    .B1(_20479_),
    .X(_00636_));
 sky130_fd_sc_hd__buf_1 _26741_ (.A(_19309_),
    .X(_20480_));
 sky130_vsdinv _26742_ (.A(\cpuregs[14][20] ),
    .Y(_20481_));
 sky130_fd_sc_hd__nor2_4 _26743_ (.A(_20481_),
    .B(_19807_),
    .Y(_20482_));
 sky130_fd_sc_hd__a211o_4 _26744_ (.A1(\cpuregs[15][20] ),
    .A2(_20480_),
    .B1(_19805_),
    .C1(_20482_),
    .X(_20483_));
 sky130_fd_sc_hd__buf_1 _26745_ (.A(_19318_),
    .X(_20484_));
 sky130_vsdinv _26746_ (.A(\cpuregs[12][20] ),
    .Y(_20485_));
 sky130_fd_sc_hd__nor2_4 _26747_ (.A(_20485_),
    .B(_19812_),
    .Y(_20486_));
 sky130_fd_sc_hd__a211o_4 _26748_ (.A1(\cpuregs[13][20] ),
    .A2(_20484_),
    .B1(_19810_),
    .C1(_20486_),
    .X(_20487_));
 sky130_fd_sc_hd__a21o_4 _26749_ (.A1(_20483_),
    .A2(_20487_),
    .B1(_19815_),
    .X(_20488_));
 sky130_vsdinv _26750_ (.A(\cpuregs[8][20] ),
    .Y(_20489_));
 sky130_fd_sc_hd__nor2_4 _26751_ (.A(_20489_),
    .B(_19878_),
    .Y(_20490_));
 sky130_fd_sc_hd__a211o_4 _26752_ (.A1(\cpuregs[9][20] ),
    .A2(_19817_),
    .B1(_19876_),
    .C1(_20490_),
    .X(_20491_));
 sky130_fd_sc_hd__buf_1 _26753_ (.A(_19344_),
    .X(_20492_));
 sky130_vsdinv _26754_ (.A(\cpuregs[10][20] ),
    .Y(_20493_));
 sky130_fd_sc_hd__nor2_4 _26755_ (.A(_20493_),
    .B(_19882_),
    .Y(_20494_));
 sky130_fd_sc_hd__a211o_4 _26756_ (.A1(\cpuregs[11][20] ),
    .A2(_20291_),
    .B1(_20492_),
    .C1(_20494_),
    .X(_20495_));
 sky130_fd_sc_hd__buf_1 _26757_ (.A(_19472_),
    .X(_20496_));
 sky130_fd_sc_hd__a21o_4 _26758_ (.A1(_20491_),
    .A2(_20495_),
    .B1(_20496_),
    .X(_20497_));
 sky130_fd_sc_hd__buf_1 _26759_ (.A(_19326_),
    .X(_20498_));
 sky130_fd_sc_hd__nand3_4 _26760_ (.A(_20488_),
    .B(_20497_),
    .C(_20498_),
    .Y(_20499_));
 sky130_fd_sc_hd__and2_4 _26761_ (.A(_20499_),
    .B(_19887_),
    .X(_20500_));
 sky130_fd_sc_hd__and2_4 _26762_ (.A(_19889_),
    .B(\cpuregs[0][20] ),
    .X(_20501_));
 sky130_fd_sc_hd__a211o_4 _26763_ (.A1(\cpuregs[1][20] ),
    .A2(_20298_),
    .B1(_19831_),
    .C1(_20501_),
    .X(_20502_));
 sky130_vsdinv _26764_ (.A(\cpuregs[2][20] ),
    .Y(_20503_));
 sky130_fd_sc_hd__nor2_4 _26765_ (.A(_20503_),
    .B(_20303_),
    .Y(_20504_));
 sky130_fd_sc_hd__a211o_4 _26766_ (.A1(\cpuregs[3][20] ),
    .A2(_19893_),
    .B1(_20301_),
    .C1(_20504_),
    .X(_20505_));
 sky130_fd_sc_hd__a21o_4 _26767_ (.A1(_20502_),
    .A2(_20505_),
    .B1(_19897_),
    .X(_20506_));
 sky130_vsdinv _26768_ (.A(\cpuregs[6][20] ),
    .Y(_20507_));
 sky130_fd_sc_hd__nor2_4 _26769_ (.A(_20507_),
    .B(_20309_),
    .Y(_20508_));
 sky130_fd_sc_hd__a211o_4 _26770_ (.A1(\cpuregs[7][20] ),
    .A2(_19899_),
    .B1(_20307_),
    .C1(_20508_),
    .X(_20509_));
 sky130_vsdinv _26771_ (.A(\cpuregs[4][20] ),
    .Y(_20510_));
 sky130_fd_sc_hd__nor2_4 _26772_ (.A(_20510_),
    .B(_20313_),
    .Y(_20511_));
 sky130_fd_sc_hd__a211o_4 _26773_ (.A1(\cpuregs[5][20] ),
    .A2(_19845_),
    .B1(_19846_),
    .C1(_20511_),
    .X(_20512_));
 sky130_fd_sc_hd__a21o_4 _26774_ (.A1(_20509_),
    .A2(_20512_),
    .B1(_19851_),
    .X(_20513_));
 sky130_fd_sc_hd__nand3_4 _26775_ (.A(_20506_),
    .B(_19838_),
    .C(_20513_),
    .Y(_20514_));
 sky130_fd_sc_hd__buf_1 _26776_ (.A(_19383_),
    .X(_20515_));
 sky130_fd_sc_hd__buf_1 _26777_ (.A(_19639_),
    .X(_20516_));
 sky130_vsdinv _26778_ (.A(\cpuregs[18][20] ),
    .Y(_20517_));
 sky130_fd_sc_hd__buf_1 _26779_ (.A(_19643_),
    .X(_20518_));
 sky130_fd_sc_hd__nor2_4 _26780_ (.A(_20517_),
    .B(_20518_),
    .Y(_20519_));
 sky130_fd_sc_hd__a211o_4 _26781_ (.A1(\cpuregs[19][20] ),
    .A2(_20516_),
    .B1(_19908_),
    .C1(_20519_),
    .X(_20520_));
 sky130_vsdinv _26782_ (.A(\cpuregs[16][20] ),
    .Y(_20521_));
 sky130_fd_sc_hd__nor2_4 _26783_ (.A(_20521_),
    .B(_19915_),
    .Y(_20522_));
 sky130_fd_sc_hd__a211o_4 _26784_ (.A1(\cpuregs[17][20] ),
    .A2(_19912_),
    .B1(_19913_),
    .C1(_20522_),
    .X(_20523_));
 sky130_fd_sc_hd__a21oi_4 _26785_ (.A1(_20520_),
    .A2(_20523_),
    .B1(_19918_),
    .Y(_20524_));
 sky130_fd_sc_hd__a2111o_4 _26786_ (.A1(_20500_),
    .A2(_20514_),
    .B1(_20318_),
    .C1(_20515_),
    .D1(_20524_),
    .X(_20525_));
 sky130_vsdinv _26787_ (.A(\timer[20] ),
    .Y(_20526_));
 sky130_fd_sc_hd__a41o_4 _26788_ (.A1(_20379_),
    .A2(_20383_),
    .A3(_20377_),
    .A4(_20434_),
    .B1(_20526_),
    .X(_20527_));
 sky130_fd_sc_hd__nand3_4 _26789_ (.A(_20433_),
    .B(_20526_),
    .C(_20435_),
    .Y(_20528_));
 sky130_vsdinv _26790_ (.A(_19419_),
    .Y(_20529_));
 sky130_fd_sc_hd__a21o_4 _26791_ (.A1(_20527_),
    .A2(_20528_),
    .B1(_20529_),
    .X(_20530_));
 sky130_fd_sc_hd__a21oi_4 _26792_ (.A1(_20525_),
    .A2(_20530_),
    .B1(_20333_),
    .Y(_00638_));
 sky130_vsdinv _26793_ (.A(_19161_),
    .Y(_20531_));
 sky130_fd_sc_hd__buf_1 _26794_ (.A(_18925_),
    .X(_20532_));
 sky130_fd_sc_hd__and4_4 _26795_ (.A(_20433_),
    .B(_20531_),
    .C(_20532_),
    .D(_20435_),
    .X(_20533_));
 sky130_fd_sc_hd__a21o_4 _26796_ (.A1(_20528_),
    .A2(\timer[21] ),
    .B1(_20381_),
    .X(_20534_));
 sky130_fd_sc_hd__buf_1 _26797_ (.A(_19455_),
    .X(_20535_));
 sky130_vsdinv _26798_ (.A(\cpuregs[14][21] ),
    .Y(_20536_));
 sky130_fd_sc_hd__nor2_4 _26799_ (.A(_20536_),
    .B(_19334_),
    .Y(_20537_));
 sky130_fd_sc_hd__a211o_4 _26800_ (.A1(\cpuregs[15][21] ),
    .A2(_20334_),
    .B1(_20535_),
    .C1(_20537_),
    .X(_20538_));
 sky130_vsdinv _26801_ (.A(\cpuregs[12][21] ),
    .Y(_20539_));
 sky130_fd_sc_hd__nor2_4 _26802_ (.A(_20539_),
    .B(_20137_),
    .Y(_20540_));
 sky130_fd_sc_hd__a211o_4 _26803_ (.A1(\cpuregs[13][21] ),
    .A2(_20446_),
    .B1(_20338_),
    .C1(_20540_),
    .X(_20541_));
 sky130_fd_sc_hd__a21o_4 _26804_ (.A1(_20538_),
    .A2(_20541_),
    .B1(_20065_),
    .X(_20542_));
 sky130_vsdinv _26805_ (.A(\cpuregs[8][21] ),
    .Y(_20543_));
 sky130_fd_sc_hd__nor2_4 _26806_ (.A(_20543_),
    .B(_19985_),
    .Y(_20544_));
 sky130_fd_sc_hd__a211o_4 _26807_ (.A1(\cpuregs[9][21] ),
    .A2(_20067_),
    .B1(_19214_),
    .C1(_20544_),
    .X(_20545_));
 sky130_vsdinv _26808_ (.A(\cpuregs[10][21] ),
    .Y(_20546_));
 sky130_fd_sc_hd__nor2_4 _26809_ (.A(_20546_),
    .B(_19990_),
    .Y(_20547_));
 sky130_fd_sc_hd__a211o_4 _26810_ (.A1(\cpuregs[11][21] ),
    .A2(_19988_),
    .B1(_19456_),
    .C1(_20547_),
    .X(_20548_));
 sky130_fd_sc_hd__a21o_4 _26811_ (.A1(_20545_),
    .A2(_20548_),
    .B1(_20015_),
    .X(_20549_));
 sky130_fd_sc_hd__nand3_4 _26812_ (.A(_20542_),
    .B(_20549_),
    .C(_20076_),
    .Y(_20550_));
 sky130_fd_sc_hd__and2_4 _26813_ (.A(_20550_),
    .B(_20078_),
    .X(_20551_));
 sky130_fd_sc_hd__and2_4 _26814_ (.A(_20007_),
    .B(\cpuregs[0][21] ),
    .X(_20552_));
 sky130_fd_sc_hd__a211o_4 _26815_ (.A1(\cpuregs[1][21] ),
    .A2(_19459_),
    .B1(_20083_),
    .C1(_20552_),
    .X(_20553_));
 sky130_vsdinv _26816_ (.A(\cpuregs[2][21] ),
    .Y(_20554_));
 sky130_fd_sc_hd__nor2_4 _26817_ (.A(_20554_),
    .B(_19969_),
    .Y(_20555_));
 sky130_fd_sc_hd__a211o_4 _26818_ (.A1(\cpuregs[3][21] ),
    .A2(_19198_),
    .B1(_19202_),
    .C1(_20555_),
    .X(_20556_));
 sky130_fd_sc_hd__a21o_4 _26819_ (.A1(_20553_),
    .A2(_20556_),
    .B1(_20016_),
    .X(_20557_));
 sky130_vsdinv _26820_ (.A(\cpuregs[6][21] ),
    .Y(_20558_));
 sky130_fd_sc_hd__nor2_4 _26821_ (.A(_20558_),
    .B(_19395_),
    .Y(_20559_));
 sky130_fd_sc_hd__a211o_4 _26822_ (.A1(\cpuregs[7][21] ),
    .A2(_20032_),
    .B1(_20035_),
    .C1(_20559_),
    .X(_20560_));
 sky130_vsdinv _26823_ (.A(\cpuregs[4][21] ),
    .Y(_20561_));
 sky130_fd_sc_hd__nor2_4 _26824_ (.A(_20561_),
    .B(_19405_),
    .Y(_20562_));
 sky130_fd_sc_hd__a211o_4 _26825_ (.A1(\cpuregs[5][21] ),
    .A2(_19740_),
    .B1(_19720_),
    .C1(_20562_),
    .X(_20563_));
 sky130_fd_sc_hd__a21o_4 _26826_ (.A1(_20560_),
    .A2(_20563_),
    .B1(_19539_),
    .X(_20564_));
 sky130_fd_sc_hd__nand3_4 _26827_ (.A(_20557_),
    .B(_20018_),
    .C(_20564_),
    .Y(_20565_));
 sky130_vsdinv _26828_ (.A(\cpuregs[18][21] ),
    .Y(_20566_));
 sky130_fd_sc_hd__nor2_4 _26829_ (.A(_20566_),
    .B(_20367_),
    .Y(_20567_));
 sky130_fd_sc_hd__a211o_4 _26830_ (.A1(\cpuregs[19][21] ),
    .A2(_19210_),
    .B1(_20036_),
    .C1(_20567_),
    .X(_20568_));
 sky130_vsdinv _26831_ (.A(\cpuregs[16][21] ),
    .Y(_20569_));
 sky130_fd_sc_hd__nor2_4 _26832_ (.A(_20569_),
    .B(_20045_),
    .Y(_20570_));
 sky130_fd_sc_hd__a211o_4 _26833_ (.A1(\cpuregs[17][21] ),
    .A2(_20041_),
    .B1(_20042_),
    .C1(_20570_),
    .X(_20571_));
 sky130_fd_sc_hd__a21oi_4 _26834_ (.A1(_20568_),
    .A2(_20571_),
    .B1(_20048_),
    .Y(_20572_));
 sky130_fd_sc_hd__a211o_4 _26835_ (.A1(_20551_),
    .A2(_20565_),
    .B1(_20031_),
    .C1(_20572_),
    .X(_20573_));
 sky130_fd_sc_hd__a21oi_4 _26836_ (.A1(_20573_),
    .A2(_20429_),
    .B1(_20430_),
    .Y(_20574_));
 sky130_fd_sc_hd__o21a_4 _26837_ (.A1(_20533_),
    .A2(_20534_),
    .B1(_20574_),
    .X(_00639_));
 sky130_fd_sc_hd__buf_1 _26838_ (.A(\timer[22] ),
    .X(_20575_));
 sky130_fd_sc_hd__nand4_4 _26839_ (.A(_20575_),
    .B(_20433_),
    .C(_20532_),
    .D(_20435_),
    .Y(_20576_));
 sky130_fd_sc_hd__o21ai_4 _26840_ (.A1(_20575_),
    .A2(_20533_),
    .B1(_20576_),
    .Y(_20577_));
 sky130_fd_sc_hd__and2_4 _26841_ (.A(_19337_),
    .B(\cpuregs[0][22] ),
    .X(_20578_));
 sky130_fd_sc_hd__a211o_4 _26842_ (.A1(\cpuregs[1][22] ),
    .A2(_19297_),
    .B1(_19299_),
    .C1(_20578_),
    .X(_20579_));
 sky130_vsdinv _26843_ (.A(\cpuregs[2][22] ),
    .Y(_20580_));
 sky130_fd_sc_hd__nor2_4 _26844_ (.A(_20580_),
    .B(_19315_),
    .Y(_20581_));
 sky130_fd_sc_hd__a211o_4 _26845_ (.A1(\cpuregs[3][22] ),
    .A2(_19310_),
    .B1(_19389_),
    .C1(_20581_),
    .X(_20582_));
 sky130_fd_sc_hd__a21o_4 _26846_ (.A1(_20579_),
    .A2(_20582_),
    .B1(_19240_),
    .X(_20583_));
 sky130_vsdinv _26847_ (.A(\cpuregs[6][22] ),
    .Y(_20584_));
 sky130_fd_sc_hd__nor2_4 _26848_ (.A(_20584_),
    .B(_19228_),
    .Y(_20585_));
 sky130_fd_sc_hd__a211o_4 _26849_ (.A1(\cpuregs[7][22] ),
    .A2(_19342_),
    .B1(_19345_),
    .C1(_20585_),
    .X(_20586_));
 sky130_vsdinv _26850_ (.A(\cpuregs[4][22] ),
    .Y(_20587_));
 sky130_fd_sc_hd__nor2_4 _26851_ (.A(_20587_),
    .B(_19257_),
    .Y(_20588_));
 sky130_fd_sc_hd__a211o_4 _26852_ (.A1(\cpuregs[5][22] ),
    .A2(_19556_),
    .B1(_19944_),
    .C1(_20588_),
    .X(_20589_));
 sky130_fd_sc_hd__a21o_4 _26853_ (.A1(_20586_),
    .A2(_20589_),
    .B1(_19850_),
    .X(_20590_));
 sky130_fd_sc_hd__nand3_4 _26854_ (.A(_20583_),
    .B(_19254_),
    .C(_20590_),
    .Y(_20591_));
 sky130_vsdinv _26855_ (.A(\cpuregs[14][22] ),
    .Y(_20592_));
 sky130_fd_sc_hd__nor2_4 _26856_ (.A(_20592_),
    .B(_19322_),
    .Y(_20593_));
 sky130_fd_sc_hd__a211o_4 _26857_ (.A1(\cpuregs[15][22] ),
    .A2(_19368_),
    .B1(_19320_),
    .C1(_20593_),
    .X(_20594_));
 sky130_vsdinv _26858_ (.A(\cpuregs[12][22] ),
    .Y(_20595_));
 sky130_fd_sc_hd__nor2_4 _26859_ (.A(_20595_),
    .B(_19257_),
    .Y(_20596_));
 sky130_fd_sc_hd__a211o_4 _26860_ (.A1(\cpuregs[13][22] ),
    .A2(_19574_),
    .B1(_19830_),
    .C1(_20596_),
    .X(_20597_));
 sky130_fd_sc_hd__a21o_4 _26861_ (.A1(_20594_),
    .A2(_20597_),
    .B1(_19850_),
    .X(_20598_));
 sky130_vsdinv _26862_ (.A(\cpuregs[8][22] ),
    .Y(_20599_));
 sky130_fd_sc_hd__nor2_4 _26863_ (.A(_20599_),
    .B(_19172_),
    .Y(_20600_));
 sky130_fd_sc_hd__a211o_4 _26864_ (.A1(\cpuregs[9][22] ),
    .A2(_19556_),
    .B1(_19944_),
    .C1(_20600_),
    .X(_20601_));
 sky130_vsdinv _26865_ (.A(\cpuregs[10][22] ),
    .Y(_20602_));
 sky130_fd_sc_hd__nor2_4 _26866_ (.A(_20602_),
    .B(_19234_),
    .Y(_20603_));
 sky130_fd_sc_hd__a211o_4 _26867_ (.A1(\cpuregs[11][22] ),
    .A2(_19399_),
    .B1(_19230_),
    .C1(_20603_),
    .X(_20604_));
 sky130_fd_sc_hd__a21o_4 _26868_ (.A1(_20601_),
    .A2(_20604_),
    .B1(_19263_),
    .X(_20605_));
 sky130_fd_sc_hd__nand3_4 _26869_ (.A(_20598_),
    .B(_20605_),
    .C(_19327_),
    .Y(_20606_));
 sky130_fd_sc_hd__nand3_4 _26870_ (.A(_20591_),
    .B(_19522_),
    .C(_20606_),
    .Y(_20607_));
 sky130_vsdinv _26871_ (.A(\cpuregs[18][22] ),
    .Y(_20608_));
 sky130_fd_sc_hd__nor2_4 _26872_ (.A(_20608_),
    .B(_19547_),
    .Y(_20609_));
 sky130_fd_sc_hd__a211o_4 _26873_ (.A1(\cpuregs[19][22] ),
    .A2(_19545_),
    .B1(_19390_),
    .C1(_20609_),
    .X(_20610_));
 sky130_fd_sc_hd__buf_1 _26874_ (.A(_19236_),
    .X(_20611_));
 sky130_vsdinv _26875_ (.A(\cpuregs[16][22] ),
    .Y(_20612_));
 sky130_fd_sc_hd__nor2_4 _26876_ (.A(_20612_),
    .B(_19258_),
    .Y(_20613_));
 sky130_fd_sc_hd__a211o_4 _26877_ (.A1(\cpuregs[17][22] ),
    .A2(_19969_),
    .B1(_20611_),
    .C1(_20613_),
    .X(_20614_));
 sky130_fd_sc_hd__a21oi_4 _26878_ (.A1(_20610_),
    .A2(_20614_),
    .B1(_19278_),
    .Y(_20615_));
 sky130_fd_sc_hd__nor2_4 _26879_ (.A(_19381_),
    .B(_20615_),
    .Y(_20616_));
 sky130_fd_sc_hd__nand2_4 _26880_ (.A(_20607_),
    .B(_20616_),
    .Y(_20617_));
 sky130_fd_sc_hd__a21o_4 _26881_ (.A1(_20617_),
    .A2(_19976_),
    .B1(_19977_),
    .X(_20618_));
 sky130_fd_sc_hd__a21oi_4 _26882_ (.A1(_20577_),
    .A2(_19166_),
    .B1(_20618_),
    .Y(_00640_));
 sky130_vsdinv _26883_ (.A(\cpuregs[14][23] ),
    .Y(_20619_));
 sky130_fd_sc_hd__nor2_4 _26884_ (.A(_20619_),
    .B(_19512_),
    .Y(_20620_));
 sky130_fd_sc_hd__a211o_4 _26885_ (.A1(\cpuregs[15][23] ),
    .A2(_20057_),
    .B1(_20058_),
    .C1(_20620_),
    .X(_20621_));
 sky130_vsdinv _26886_ (.A(\cpuregs[12][23] ),
    .Y(_20622_));
 sky130_fd_sc_hd__nor2_4 _26887_ (.A(_20622_),
    .B(_19525_),
    .Y(_20623_));
 sky130_fd_sc_hd__a211o_4 _26888_ (.A1(\cpuregs[13][23] ),
    .A2(_19269_),
    .B1(_19271_),
    .C1(_20623_),
    .X(_20624_));
 sky130_fd_sc_hd__a21o_4 _26889_ (.A1(_20621_),
    .A2(_20624_),
    .B1(_19252_),
    .X(_20625_));
 sky130_vsdinv _26890_ (.A(\cpuregs[8][23] ),
    .Y(_20626_));
 sky130_fd_sc_hd__nor2_4 _26891_ (.A(_20626_),
    .B(_19609_),
    .Y(_20627_));
 sky130_fd_sc_hd__a211o_4 _26892_ (.A1(\cpuregs[9][23] ),
    .A2(_20446_),
    .B1(_20338_),
    .C1(_20627_),
    .X(_20628_));
 sky130_vsdinv _26893_ (.A(\cpuregs[10][23] ),
    .Y(_20629_));
 sky130_fd_sc_hd__nor2_4 _26894_ (.A(_20629_),
    .B(_19429_),
    .Y(_20630_));
 sky130_fd_sc_hd__a211o_4 _26895_ (.A1(\cpuregs[11][23] ),
    .A2(_19481_),
    .B1(_20450_),
    .C1(_20630_),
    .X(_20631_));
 sky130_fd_sc_hd__a21o_4 _26896_ (.A1(_20628_),
    .A2(_20631_),
    .B1(_19473_),
    .X(_20632_));
 sky130_fd_sc_hd__nand3_4 _26897_ (.A(_20625_),
    .B(_20632_),
    .C(_19276_),
    .Y(_20633_));
 sky130_fd_sc_hd__and2_4 _26898_ (.A(_20633_),
    .B(_20078_),
    .X(_20634_));
 sky130_fd_sc_hd__and2_4 _26899_ (.A(_20084_),
    .B(\cpuregs[0][23] ),
    .X(_20635_));
 sky130_fd_sc_hd__a211o_4 _26900_ (.A1(\cpuregs[1][23] ),
    .A2(_20081_),
    .B1(_20083_),
    .C1(_20635_),
    .X(_20636_));
 sky130_vsdinv _26901_ (.A(\cpuregs[2][23] ),
    .Y(_20637_));
 sky130_fd_sc_hd__nor2_4 _26902_ (.A(_20637_),
    .B(_19545_),
    .Y(_20638_));
 sky130_fd_sc_hd__a211o_4 _26903_ (.A1(\cpuregs[3][23] ),
    .A2(_20081_),
    .B1(_20087_),
    .C1(_20638_),
    .X(_20639_));
 sky130_fd_sc_hd__a21o_4 _26904_ (.A1(_20636_),
    .A2(_20639_),
    .B1(_19474_),
    .X(_20640_));
 sky130_vsdinv _26905_ (.A(\cpuregs[6][23] ),
    .Y(_20641_));
 sky130_fd_sc_hd__nor2_4 _26906_ (.A(_20641_),
    .B(_20044_),
    .Y(_20642_));
 sky130_fd_sc_hd__a211o_4 _26907_ (.A1(\cpuregs[7][23] ),
    .A2(_19469_),
    .B1(_20087_),
    .C1(_20642_),
    .X(_20643_));
 sky130_vsdinv _26908_ (.A(\cpuregs[4][23] ),
    .Y(_20644_));
 sky130_fd_sc_hd__nor2_4 _26909_ (.A(_20644_),
    .B(_19430_),
    .Y(_20645_));
 sky130_fd_sc_hd__a211o_4 _26910_ (.A1(\cpuregs[5][23] ),
    .A2(_20093_),
    .B1(_19215_),
    .C1(_20645_),
    .X(_20646_));
 sky130_fd_sc_hd__a21o_4 _26911_ (.A1(_20643_),
    .A2(_20646_),
    .B1(_19463_),
    .X(_20647_));
 sky130_fd_sc_hd__nand3_4 _26912_ (.A(_20640_),
    .B(_19477_),
    .C(_20647_),
    .Y(_20648_));
 sky130_fd_sc_hd__buf_1 _26913_ (.A(_20155_),
    .X(_20649_));
 sky130_vsdinv _26914_ (.A(\cpuregs[18][23] ),
    .Y(_20650_));
 sky130_fd_sc_hd__nor2_4 _26915_ (.A(_20650_),
    .B(_19558_),
    .Y(_20651_));
 sky130_fd_sc_hd__a211o_4 _26916_ (.A1(\cpuregs[19][23] ),
    .A2(_19483_),
    .B1(_19203_),
    .C1(_20651_),
    .X(_20652_));
 sky130_vsdinv _26917_ (.A(\cpuregs[16][23] ),
    .Y(_20653_));
 sky130_fd_sc_hd__nor2_4 _26918_ (.A(_20653_),
    .B(_20367_),
    .Y(_20654_));
 sky130_fd_sc_hd__a211o_4 _26919_ (.A1(\cpuregs[17][23] ),
    .A2(_19199_),
    .B1(_19216_),
    .C1(_20654_),
    .X(_20655_));
 sky130_fd_sc_hd__a21oi_4 _26920_ (.A1(_20652_),
    .A2(_20655_),
    .B1(_19225_),
    .Y(_20656_));
 sky130_fd_sc_hd__a211o_4 _26921_ (.A1(_20634_),
    .A2(_20648_),
    .B1(_20649_),
    .C1(_20656_),
    .X(_20657_));
 sky130_fd_sc_hd__and4_4 _26922_ (.A(_20378_),
    .B(_20383_),
    .C(_20376_),
    .D(_20434_),
    .X(_20658_));
 sky130_vsdinv _26923_ (.A(_20575_),
    .Y(_20659_));
 sky130_fd_sc_hd__and4_4 _26924_ (.A(_20658_),
    .B(\timer[23] ),
    .C(_20659_),
    .D(_20532_),
    .X(_20660_));
 sky130_fd_sc_hd__and4_4 _26925_ (.A(_20432_),
    .B(_20659_),
    .C(_20532_),
    .D(_20434_),
    .X(_20661_));
 sky130_fd_sc_hd__o21ai_4 _26926_ (.A1(\timer[23] ),
    .A2(_20661_),
    .B1(_19420_),
    .Y(_20662_));
 sky130_fd_sc_hd__o22a_4 _26927_ (.A1(_19380_),
    .A2(_20657_),
    .B1(_20660_),
    .B2(_20662_),
    .X(_20663_));
 sky130_fd_sc_hd__nor2_4 _26928_ (.A(_19427_),
    .B(_20663_),
    .Y(_00641_));
 sky130_vsdinv _26929_ (.A(\cpuregs[14][24] ),
    .Y(_20664_));
 sky130_fd_sc_hd__nor2_4 _26930_ (.A(_20664_),
    .B(_19511_),
    .Y(_20665_));
 sky130_fd_sc_hd__a211o_4 _26931_ (.A1(\cpuregs[15][24] ),
    .A2(_19444_),
    .B1(_19230_),
    .C1(_20665_),
    .X(_20666_));
 sky130_vsdinv _26932_ (.A(\cpuregs[12][24] ),
    .Y(_20667_));
 sky130_fd_sc_hd__nor2_4 _26933_ (.A(_20667_),
    .B(_19524_),
    .Y(_20668_));
 sky130_fd_sc_hd__a211o_4 _26934_ (.A1(\cpuregs[13][24] ),
    .A2(_19444_),
    .B1(_19236_),
    .C1(_20668_),
    .X(_20669_));
 sky130_fd_sc_hd__a21o_4 _26935_ (.A1(_20666_),
    .A2(_20669_),
    .B1(_19251_),
    .X(_20670_));
 sky130_vsdinv _26936_ (.A(\cpuregs[8][24] ),
    .Y(_20671_));
 sky130_fd_sc_hd__nor2_4 _26937_ (.A(_20671_),
    .B(_19573_),
    .Y(_20672_));
 sky130_fd_sc_hd__a211o_4 _26938_ (.A1(\cpuregs[9][24] ),
    .A2(_19444_),
    .B1(_19270_),
    .C1(_20672_),
    .X(_20673_));
 sky130_vsdinv _26939_ (.A(\cpuregs[10][24] ),
    .Y(_20674_));
 sky130_fd_sc_hd__nor2_4 _26940_ (.A(_20674_),
    .B(_19296_),
    .Y(_20675_));
 sky130_fd_sc_hd__a211o_4 _26941_ (.A1(\cpuregs[11][24] ),
    .A2(_19480_),
    .B1(_19200_),
    .C1(_20675_),
    .X(_20676_));
 sky130_fd_sc_hd__a21o_4 _26942_ (.A1(_20673_),
    .A2(_20676_),
    .B1(_19263_),
    .X(_20677_));
 sky130_fd_sc_hd__nand3_4 _26943_ (.A(_20670_),
    .B(_20677_),
    .C(_19327_),
    .Y(_20678_));
 sky130_fd_sc_hd__and2_4 _26944_ (.A(_20678_),
    .B(_19278_),
    .X(_20679_));
 sky130_fd_sc_hd__buf_1 _26945_ (.A(_20679_),
    .X(_20680_));
 sky130_fd_sc_hd__and2_4 _26946_ (.A(_19205_),
    .B(\cpuregs[0][24] ),
    .X(_20681_));
 sky130_fd_sc_hd__a211o_4 _26947_ (.A1(\cpuregs[1][24] ),
    .A2(_19235_),
    .B1(_19247_),
    .C1(_20681_),
    .X(_20682_));
 sky130_vsdinv _26948_ (.A(\cpuregs[2][24] ),
    .Y(_20683_));
 sky130_fd_sc_hd__nor2_4 _26949_ (.A(_20683_),
    .B(_19822_),
    .Y(_20684_));
 sky130_fd_sc_hd__a211o_4 _26950_ (.A1(\cpuregs[3][24] ),
    .A2(_20057_),
    .B1(_20058_),
    .C1(_20684_),
    .X(_20685_));
 sky130_fd_sc_hd__a21o_4 _26951_ (.A1(_20682_),
    .A2(_20685_),
    .B1(_19264_),
    .X(_20686_));
 sky130_vsdinv _26952_ (.A(\cpuregs[6][24] ),
    .Y(_20687_));
 sky130_fd_sc_hd__nor2_4 _26953_ (.A(_20687_),
    .B(_19319_),
    .Y(_20688_));
 sky130_fd_sc_hd__a211o_4 _26954_ (.A1(\cpuregs[7][24] ),
    .A2(_19445_),
    .B1(_20535_),
    .C1(_20688_),
    .X(_20689_));
 sky130_vsdinv _26955_ (.A(\cpuregs[4][24] ),
    .Y(_20690_));
 sky130_fd_sc_hd__nor2_4 _26956_ (.A(_20690_),
    .B(_19531_),
    .Y(_20691_));
 sky130_fd_sc_hd__a211o_4 _26957_ (.A1(\cpuregs[5][24] ),
    .A2(_20067_),
    .B1(_20068_),
    .C1(_20691_),
    .X(_20692_));
 sky130_fd_sc_hd__a21o_4 _26958_ (.A1(_20689_),
    .A2(_20692_),
    .B1(_19584_),
    .X(_20693_));
 sky130_fd_sc_hd__nand3_4 _26959_ (.A(_20686_),
    .B(_19476_),
    .C(_20693_),
    .Y(_20694_));
 sky130_fd_sc_hd__buf_1 _26960_ (.A(_20694_),
    .X(_20695_));
 sky130_vsdinv _26961_ (.A(\cpuregs[18][24] ),
    .Y(_20696_));
 sky130_fd_sc_hd__nor2_4 _26962_ (.A(_20696_),
    .B(_20032_),
    .Y(_20697_));
 sky130_fd_sc_hd__a211o_4 _26963_ (.A1(\cpuregs[19][24] ),
    .A2(_19482_),
    .B1(_19457_),
    .C1(_20697_),
    .X(_20698_));
 sky130_vsdinv _26964_ (.A(\cpuregs[16][24] ),
    .Y(_20699_));
 sky130_fd_sc_hd__nor2_4 _26965_ (.A(_20699_),
    .B(_19773_),
    .Y(_20700_));
 sky130_fd_sc_hd__a211o_4 _26966_ (.A1(\cpuregs[17][24] ),
    .A2(_19482_),
    .B1(_19452_),
    .C1(_20700_),
    .X(_20701_));
 sky130_fd_sc_hd__a21oi_4 _26967_ (.A1(_20698_),
    .A2(_20701_),
    .B1(_19330_),
    .Y(_20702_));
 sky130_fd_sc_hd__buf_1 _26968_ (.A(_20702_),
    .X(_20703_));
 sky130_fd_sc_hd__a2111o_4 _26969_ (.A1(_20680_),
    .A2(_20695_),
    .B1(_20318_),
    .C1(_20515_),
    .D1(_20703_),
    .X(_20704_));
 sky130_fd_sc_hd__buf_1 _26970_ (.A(_18926_),
    .X(_20705_));
 sky130_fd_sc_hd__buf_1 _26971_ (.A(_20705_),
    .X(_20706_));
 sky130_fd_sc_hd__buf_1 _26972_ (.A(_18927_),
    .X(_20707_));
 sky130_fd_sc_hd__buf_1 _26973_ (.A(_20707_),
    .X(_20708_));
 sky130_fd_sc_hd__a41oi_4 _26974_ (.A1(_20330_),
    .A2(_20173_),
    .A3(_20172_),
    .A4(_20706_),
    .B1(_20708_),
    .Y(_20709_));
 sky130_fd_sc_hd__and4_4 _26975_ (.A(_20177_),
    .B(_19925_),
    .C(_20707_),
    .D(_20705_),
    .X(_20710_));
 sky130_fd_sc_hd__o21ai_4 _26976_ (.A1(_20709_),
    .A2(_20710_),
    .B1(_19867_),
    .Y(_20711_));
 sky130_fd_sc_hd__a21oi_4 _26977_ (.A1(_20704_),
    .A2(_20711_),
    .B1(_20333_),
    .Y(_00642_));
 sky130_vsdinv _26978_ (.A(\cpuregs[14][25] ),
    .Y(_20712_));
 sky130_fd_sc_hd__nor2_4 _26979_ (.A(_20712_),
    .B(_19368_),
    .Y(_20713_));
 sky130_fd_sc_hd__a211o_4 _26980_ (.A1(\cpuregs[15][25] ),
    .A2(_19269_),
    .B1(_20535_),
    .C1(_20713_),
    .X(_20714_));
 sky130_vsdinv _26981_ (.A(\cpuregs[12][25] ),
    .Y(_20715_));
 sky130_fd_sc_hd__nor2_4 _26982_ (.A(_20715_),
    .B(_19609_),
    .Y(_20716_));
 sky130_fd_sc_hd__a211o_4 _26983_ (.A1(\cpuregs[13][25] ),
    .A2(_19468_),
    .B1(_20068_),
    .C1(_20716_),
    .X(_20717_));
 sky130_fd_sc_hd__a21o_4 _26984_ (.A1(_20714_),
    .A2(_20717_),
    .B1(_20065_),
    .X(_20718_));
 sky130_vsdinv _26985_ (.A(\cpuregs[8][25] ),
    .Y(_20719_));
 sky130_fd_sc_hd__nor2_4 _26986_ (.A(_20719_),
    .B(_19429_),
    .Y(_20720_));
 sky130_fd_sc_hd__a211o_4 _26987_ (.A1(\cpuregs[9][25] ),
    .A2(_19481_),
    .B1(_19578_),
    .C1(_20720_),
    .X(_20721_));
 sky130_vsdinv _26988_ (.A(\cpuregs[10][25] ),
    .Y(_20722_));
 sky130_fd_sc_hd__nor2_4 _26989_ (.A(_20722_),
    .B(_19433_),
    .Y(_20723_));
 sky130_fd_sc_hd__a211o_4 _26990_ (.A1(\cpuregs[11][25] ),
    .A2(_19501_),
    .B1(_19287_),
    .C1(_20723_),
    .X(_20724_));
 sky130_fd_sc_hd__a21o_4 _26991_ (.A1(_20721_),
    .A2(_20724_),
    .B1(_20015_),
    .X(_20725_));
 sky130_fd_sc_hd__nand3_4 _26992_ (.A(_20718_),
    .B(_20725_),
    .C(_20076_),
    .Y(_20726_));
 sky130_fd_sc_hd__and2_4 _26993_ (.A(_20726_),
    .B(_19603_),
    .X(_20727_));
 sky130_fd_sc_hd__and2_4 _26994_ (.A(_20007_),
    .B(\cpuregs[0][25] ),
    .X(_20728_));
 sky130_fd_sc_hd__a211o_4 _26995_ (.A1(\cpuregs[1][25] ),
    .A2(_20093_),
    .B1(_19215_),
    .C1(_20728_),
    .X(_20729_));
 sky130_vsdinv _26996_ (.A(\cpuregs[2][25] ),
    .Y(_20730_));
 sky130_fd_sc_hd__nor2_4 _26997_ (.A(_20730_),
    .B(_19434_),
    .Y(_20731_));
 sky130_fd_sc_hd__a211o_4 _26998_ (.A1(\cpuregs[3][25] ),
    .A2(_19335_),
    .B1(_19633_),
    .C1(_20731_),
    .X(_20732_));
 sky130_fd_sc_hd__a21o_4 _26999_ (.A1(_20729_),
    .A2(_20732_),
    .B1(_20016_),
    .X(_20733_));
 sky130_vsdinv _27000_ (.A(\cpuregs[6][25] ),
    .Y(_20734_));
 sky130_fd_sc_hd__nor2_4 _27001_ (.A(_20734_),
    .B(_19405_),
    .Y(_20735_));
 sky130_fd_sc_hd__a211o_4 _27002_ (.A1(\cpuregs[7][25] ),
    .A2(_19740_),
    .B1(_19633_),
    .C1(_20735_),
    .X(_20736_));
 sky130_fd_sc_hd__buf_1 _27003_ (.A(_19830_),
    .X(_20737_));
 sky130_vsdinv _27004_ (.A(\cpuregs[4][25] ),
    .Y(_20738_));
 sky130_fd_sc_hd__nor2_4 _27005_ (.A(_20738_),
    .B(_20259_),
    .Y(_20739_));
 sky130_fd_sc_hd__a211o_4 _27006_ (.A1(\cpuregs[5][25] ),
    .A2(_19532_),
    .B1(_20737_),
    .C1(_20739_),
    .X(_20740_));
 sky130_fd_sc_hd__a21o_4 _27007_ (.A1(_20736_),
    .A2(_20740_),
    .B1(_19539_),
    .X(_20741_));
 sky130_fd_sc_hd__nand3_4 _27008_ (.A(_20733_),
    .B(_20018_),
    .C(_20741_),
    .Y(_20742_));
 sky130_vsdinv _27009_ (.A(\cpuregs[18][25] ),
    .Y(_20743_));
 sky130_fd_sc_hd__nor2_4 _27010_ (.A(_20743_),
    .B(_20045_),
    .Y(_20744_));
 sky130_fd_sc_hd__a211o_4 _27011_ (.A1(\cpuregs[19][25] ),
    .A2(_20041_),
    .B1(_19788_),
    .C1(_20744_),
    .X(_20745_));
 sky130_vsdinv _27012_ (.A(\cpuregs[16][25] ),
    .Y(_20746_));
 sky130_fd_sc_hd__nor2_4 _27013_ (.A(_20746_),
    .B(_19396_),
    .Y(_20747_));
 sky130_fd_sc_hd__a211o_4 _27014_ (.A1(\cpuregs[17][25] ),
    .A2(_19388_),
    .B1(_19792_),
    .C1(_20747_),
    .X(_20748_));
 sky130_fd_sc_hd__a21oi_4 _27015_ (.A1(_20745_),
    .A2(_20748_),
    .B1(_19796_),
    .Y(_20749_));
 sky130_fd_sc_hd__a2111o_4 _27016_ (.A1(_20727_),
    .A2(_20742_),
    .B1(_20318_),
    .C1(_20515_),
    .D1(_20749_),
    .X(_20750_));
 sky130_vsdinv _27017_ (.A(\timer[25] ),
    .Y(_20751_));
 sky130_fd_sc_hd__a41oi_4 _27018_ (.A1(_20330_),
    .A2(_20233_),
    .A3(_20708_),
    .A4(_20706_),
    .B1(_20751_),
    .Y(_20752_));
 sky130_fd_sc_hd__and4_4 _27019_ (.A(_20379_),
    .B(_20751_),
    .C(_20707_),
    .D(_20705_),
    .X(_20753_));
 sky130_fd_sc_hd__o21ai_4 _27020_ (.A1(_20752_),
    .A2(_20753_),
    .B1(_19867_),
    .Y(_20754_));
 sky130_fd_sc_hd__a21oi_4 _27021_ (.A1(_20750_),
    .A2(_20754_),
    .B1(_20333_),
    .Y(_00643_));
 sky130_vsdinv _27022_ (.A(\cpuregs[14][26] ),
    .Y(_20755_));
 sky130_fd_sc_hd__nor2_4 _27023_ (.A(_20755_),
    .B(_19580_),
    .Y(_20756_));
 sky130_fd_sc_hd__a211o_4 _27024_ (.A1(\cpuregs[15][26] ),
    .A2(_20480_),
    .B1(_20034_),
    .C1(_20756_),
    .X(_20757_));
 sky130_vsdinv _27025_ (.A(\cpuregs[12][26] ),
    .Y(_20758_));
 sky130_fd_sc_hd__nor2_4 _27026_ (.A(_20758_),
    .B(_19292_),
    .Y(_20759_));
 sky130_fd_sc_hd__a211o_4 _27027_ (.A1(\cpuregs[13][26] ),
    .A2(_20484_),
    .B1(_20082_),
    .C1(_20759_),
    .X(_20760_));
 sky130_fd_sc_hd__a21o_4 _27028_ (.A1(_20757_),
    .A2(_20760_),
    .B1(_19306_),
    .X(_20761_));
 sky130_vsdinv _27029_ (.A(\cpuregs[8][26] ),
    .Y(_20762_));
 sky130_fd_sc_hd__nor2_4 _27030_ (.A(_20762_),
    .B(_19878_),
    .Y(_20763_));
 sky130_fd_sc_hd__a211o_4 _27031_ (.A1(\cpuregs[9][26] ),
    .A2(_19593_),
    .B1(_19876_),
    .C1(_20763_),
    .X(_20764_));
 sky130_vsdinv _27032_ (.A(\cpuregs[10][26] ),
    .Y(_20765_));
 sky130_fd_sc_hd__nor2_4 _27033_ (.A(_20765_),
    .B(_19882_),
    .Y(_20766_));
 sky130_fd_sc_hd__a211o_4 _27034_ (.A1(\cpuregs[11][26] ),
    .A2(_20291_),
    .B1(_20492_),
    .C1(_20766_),
    .X(_20767_));
 sky130_fd_sc_hd__a21o_4 _27035_ (.A1(_20764_),
    .A2(_20767_),
    .B1(_20496_),
    .X(_20768_));
 sky130_fd_sc_hd__nand3_4 _27036_ (.A(_20761_),
    .B(_20768_),
    .C(_20498_),
    .Y(_20769_));
 sky130_fd_sc_hd__and2_4 _27037_ (.A(_20769_),
    .B(_19887_),
    .X(_20770_));
 sky130_fd_sc_hd__and2_4 _27038_ (.A(_19889_),
    .B(\cpuregs[0][26] ),
    .X(_20771_));
 sky130_fd_sc_hd__a211o_4 _27039_ (.A1(\cpuregs[1][26] ),
    .A2(_20298_),
    .B1(_20737_),
    .C1(_20771_),
    .X(_20772_));
 sky130_vsdinv _27040_ (.A(\cpuregs[2][26] ),
    .Y(_20773_));
 sky130_fd_sc_hd__nor2_4 _27041_ (.A(_20773_),
    .B(_20303_),
    .Y(_20774_));
 sky130_fd_sc_hd__a211o_4 _27042_ (.A1(\cpuregs[3][26] ),
    .A2(_19893_),
    .B1(_20301_),
    .C1(_20774_),
    .X(_20775_));
 sky130_fd_sc_hd__a21o_4 _27043_ (.A1(_20772_),
    .A2(_20775_),
    .B1(_19897_),
    .X(_20776_));
 sky130_vsdinv _27044_ (.A(\cpuregs[6][26] ),
    .Y(_20777_));
 sky130_fd_sc_hd__nor2_4 _27045_ (.A(_20777_),
    .B(_20309_),
    .Y(_20778_));
 sky130_fd_sc_hd__a211o_4 _27046_ (.A1(\cpuregs[7][26] ),
    .A2(_19899_),
    .B1(_20307_),
    .C1(_20778_),
    .X(_20779_));
 sky130_vsdinv _27047_ (.A(\cpuregs[4][26] ),
    .Y(_20780_));
 sky130_fd_sc_hd__nor2_4 _27048_ (.A(_20780_),
    .B(_20313_),
    .Y(_20781_));
 sky130_fd_sc_hd__a211o_4 _27049_ (.A1(\cpuregs[5][26] ),
    .A2(_20089_),
    .B1(_20611_),
    .C1(_20781_),
    .X(_20782_));
 sky130_fd_sc_hd__a21o_4 _27050_ (.A1(_20779_),
    .A2(_20782_),
    .B1(_19438_),
    .X(_20783_));
 sky130_fd_sc_hd__nand3_4 _27051_ (.A(_20776_),
    .B(_19255_),
    .C(_20783_),
    .Y(_20784_));
 sky130_fd_sc_hd__buf_1 _27052_ (.A(_19164_),
    .X(_20785_));
 sky130_vsdinv _27053_ (.A(\cpuregs[18][26] ),
    .Y(_20786_));
 sky130_fd_sc_hd__nor2_4 _27054_ (.A(_20786_),
    .B(_20518_),
    .Y(_20787_));
 sky130_fd_sc_hd__a211o_4 _27055_ (.A1(\cpuregs[19][26] ),
    .A2(_20516_),
    .B1(_19908_),
    .C1(_20787_),
    .X(_20788_));
 sky130_vsdinv _27056_ (.A(\cpuregs[16][26] ),
    .Y(_20789_));
 sky130_fd_sc_hd__nor2_4 _27057_ (.A(_20789_),
    .B(_19915_),
    .Y(_20790_));
 sky130_fd_sc_hd__a211o_4 _27058_ (.A1(\cpuregs[17][26] ),
    .A2(_19912_),
    .B1(_19913_),
    .C1(_20790_),
    .X(_20791_));
 sky130_fd_sc_hd__a21oi_4 _27059_ (.A1(_20788_),
    .A2(_20791_),
    .B1(_19918_),
    .Y(_20792_));
 sky130_fd_sc_hd__a2111o_4 _27060_ (.A1(_20770_),
    .A2(_20784_),
    .B1(_20785_),
    .C1(_20515_),
    .D1(_20792_),
    .X(_20793_));
 sky130_fd_sc_hd__nand4_4 _27061_ (.A(_20751_),
    .B(_20379_),
    .C(_20707_),
    .D(_20705_),
    .Y(_20794_));
 sky130_fd_sc_hd__nand2_4 _27062_ (.A(_20794_),
    .B(\timer[26] ),
    .Y(_20795_));
 sky130_fd_sc_hd__nand4_4 _27063_ (.A(_20708_),
    .B(_20388_),
    .C(_20706_),
    .D(_18929_),
    .Y(_20796_));
 sky130_fd_sc_hd__a21o_4 _27064_ (.A1(_20795_),
    .A2(_20796_),
    .B1(_20529_),
    .X(_20797_));
 sky130_fd_sc_hd__buf_1 _27065_ (.A(_19495_),
    .X(_20798_));
 sky130_fd_sc_hd__a21oi_4 _27066_ (.A1(_20793_),
    .A2(_20797_),
    .B1(_20798_),
    .Y(_00644_));
 sky130_fd_sc_hd__nand3_4 _27067_ (.A(_20710_),
    .B(_20531_),
    .C(_18929_),
    .Y(_20799_));
 sky130_fd_sc_hd__a21oi_4 _27068_ (.A1(_20799_),
    .A2(\timer[27] ),
    .B1(_19932_),
    .Y(_20800_));
 sky130_fd_sc_hd__and4_4 _27069_ (.A(_20388_),
    .B(_20708_),
    .C(_20706_),
    .D(_18929_),
    .X(_20801_));
 sky130_fd_sc_hd__nand3_4 _27070_ (.A(_20801_),
    .B(_18928_),
    .C(_20531_),
    .Y(_20802_));
 sky130_fd_sc_hd__and2_4 _27071_ (.A(_19498_),
    .B(\cpuregs[0][27] ),
    .X(_20803_));
 sky130_fd_sc_hd__a211o_4 _27072_ (.A1(\cpuregs[1][27] ),
    .A2(_20334_),
    .B1(_19247_),
    .C1(_20803_),
    .X(_20804_));
 sky130_vsdinv _27073_ (.A(\cpuregs[2][27] ),
    .Y(_20805_));
 sky130_fd_sc_hd__nor2_4 _27074_ (.A(_20805_),
    .B(_20137_),
    .Y(_20806_));
 sky130_fd_sc_hd__a211o_4 _27075_ (.A1(\cpuregs[3][27] ),
    .A2(_20446_),
    .B1(_20535_),
    .C1(_20806_),
    .X(_20807_));
 sky130_fd_sc_hd__a21o_4 _27076_ (.A1(_20804_),
    .A2(_20807_),
    .B1(_19264_),
    .X(_20808_));
 sky130_vsdinv _27077_ (.A(\cpuregs[6][27] ),
    .Y(_20809_));
 sky130_fd_sc_hd__nor2_4 _27078_ (.A(_20809_),
    .B(_19892_),
    .Y(_20810_));
 sky130_fd_sc_hd__a211o_4 _27079_ (.A1(\cpuregs[7][27] ),
    .A2(_19497_),
    .B1(_20450_),
    .C1(_20810_),
    .X(_20811_));
 sky130_fd_sc_hd__buf_1 _27080_ (.A(_19587_),
    .X(_20812_));
 sky130_vsdinv _27081_ (.A(\cpuregs[4][27] ),
    .Y(_20813_));
 sky130_fd_sc_hd__nor2_4 _27082_ (.A(_20813_),
    .B(_19399_),
    .Y(_20814_));
 sky130_fd_sc_hd__a211o_4 _27083_ (.A1(\cpuregs[5][27] ),
    .A2(_19501_),
    .B1(_20812_),
    .C1(_20814_),
    .X(_20815_));
 sky130_fd_sc_hd__a21o_4 _27084_ (.A1(_20811_),
    .A2(_20815_),
    .B1(_19462_),
    .X(_20816_));
 sky130_fd_sc_hd__nand3_4 _27085_ (.A(_20808_),
    .B(_19476_),
    .C(_20816_),
    .Y(_20817_));
 sky130_vsdinv _27086_ (.A(\cpuregs[14][27] ),
    .Y(_20818_));
 sky130_fd_sc_hd__nor2_4 _27087_ (.A(_20818_),
    .B(_19386_),
    .Y(_20819_));
 sky130_fd_sc_hd__a211o_4 _27088_ (.A1(\cpuregs[15][27] ),
    .A2(_19653_),
    .B1(_19201_),
    .C1(_20819_),
    .X(_20820_));
 sky130_vsdinv _27089_ (.A(\cpuregs[12][27] ),
    .Y(_20821_));
 sky130_fd_sc_hd__nor2_4 _27090_ (.A(_20821_),
    .B(_19659_),
    .Y(_20822_));
 sky130_fd_sc_hd__a211o_4 _27091_ (.A1(\cpuregs[13][27] ),
    .A2(_19630_),
    .B1(_19702_),
    .C1(_20822_),
    .X(_20823_));
 sky130_fd_sc_hd__a21o_4 _27092_ (.A1(_20820_),
    .A2(_20823_),
    .B1(_19706_),
    .X(_20824_));
 sky130_vsdinv _27093_ (.A(\cpuregs[8][27] ),
    .Y(_20825_));
 sky130_fd_sc_hd__nor2_4 _27094_ (.A(_20825_),
    .B(_19433_),
    .Y(_20826_));
 sky130_fd_sc_hd__a211o_4 _27095_ (.A1(\cpuregs[9][27] ),
    .A2(_19501_),
    .B1(_20812_),
    .C1(_20826_),
    .X(_20827_));
 sky130_vsdinv _27096_ (.A(\cpuregs[10][27] ),
    .Y(_20828_));
 sky130_fd_sc_hd__nor2_4 _27097_ (.A(_20828_),
    .B(_19819_),
    .Y(_20829_));
 sky130_fd_sc_hd__a211o_4 _27098_ (.A1(\cpuregs[11][27] ),
    .A2(_19507_),
    .B1(_19287_),
    .C1(_20829_),
    .X(_20830_));
 sky130_fd_sc_hd__a21o_4 _27099_ (.A1(_20827_),
    .A2(_20830_),
    .B1(_19354_),
    .X(_20831_));
 sky130_fd_sc_hd__nand3_4 _27100_ (.A(_20824_),
    .B(_20831_),
    .C(_19601_),
    .Y(_20832_));
 sky130_fd_sc_hd__nand3_4 _27101_ (.A(_20817_),
    .B(_19279_),
    .C(_20832_),
    .Y(_20833_));
 sky130_vsdinv _27102_ (.A(\cpuregs[18][27] ),
    .Y(_20834_));
 sky130_fd_sc_hd__nor2_4 _27103_ (.A(_20834_),
    .B(_19643_),
    .Y(_20835_));
 sky130_fd_sc_hd__a211o_4 _27104_ (.A1(\cpuregs[19][27] ),
    .A2(_19469_),
    .B1(_19202_),
    .C1(_20835_),
    .X(_20836_));
 sky130_vsdinv _27105_ (.A(\cpuregs[16][27] ),
    .Y(_20837_));
 sky130_fd_sc_hd__nor2_4 _27106_ (.A(_20837_),
    .B(_19434_),
    .Y(_20838_));
 sky130_fd_sc_hd__a211o_4 _27107_ (.A1(\cpuregs[17][27] ),
    .A2(_20005_),
    .B1(_20006_),
    .C1(_20838_),
    .X(_20839_));
 sky130_fd_sc_hd__a21oi_4 _27108_ (.A1(_20836_),
    .A2(_20839_),
    .B1(_19409_),
    .Y(_20840_));
 sky130_fd_sc_hd__nor2_4 _27109_ (.A(_19381_),
    .B(_20840_),
    .Y(_20841_));
 sky130_fd_sc_hd__nand2_4 _27110_ (.A(_20833_),
    .B(_20841_),
    .Y(_20842_));
 sky130_fd_sc_hd__a21o_4 _27111_ (.A1(_20842_),
    .A2(_19976_),
    .B1(_19977_),
    .X(_20843_));
 sky130_fd_sc_hd__a21oi_4 _27112_ (.A1(_20800_),
    .A2(_20802_),
    .B1(_20843_),
    .Y(_00645_));
 sky130_vsdinv _27113_ (.A(\cpuregs[14][28] ),
    .Y(_20844_));
 sky130_fd_sc_hd__nor2_4 _27114_ (.A(_20844_),
    .B(_19580_),
    .Y(_20845_));
 sky130_fd_sc_hd__a211o_4 _27115_ (.A1(\cpuregs[15][28] ),
    .A2(_20480_),
    .B1(_20034_),
    .C1(_20845_),
    .X(_20846_));
 sky130_vsdinv _27116_ (.A(\cpuregs[12][28] ),
    .Y(_20847_));
 sky130_fd_sc_hd__nor2_4 _27117_ (.A(_20847_),
    .B(_19292_),
    .Y(_20848_));
 sky130_fd_sc_hd__a211o_4 _27118_ (.A1(\cpuregs[13][28] ),
    .A2(_20484_),
    .B1(_20082_),
    .C1(_20848_),
    .X(_20849_));
 sky130_fd_sc_hd__a21o_4 _27119_ (.A1(_20846_),
    .A2(_20849_),
    .B1(_19306_),
    .X(_20850_));
 sky130_vsdinv _27120_ (.A(\cpuregs[8][28] ),
    .Y(_20851_));
 sky130_fd_sc_hd__nor2_4 _27121_ (.A(_20851_),
    .B(_19596_),
    .Y(_20852_));
 sky130_fd_sc_hd__a211o_4 _27122_ (.A1(\cpuregs[9][28] ),
    .A2(_19593_),
    .B1(_19299_),
    .C1(_20852_),
    .X(_20853_));
 sky130_vsdinv _27123_ (.A(\cpuregs[10][28] ),
    .Y(_20854_));
 sky130_fd_sc_hd__nor2_4 _27124_ (.A(_20854_),
    .B(_19730_),
    .Y(_20855_));
 sky130_fd_sc_hd__a211o_4 _27125_ (.A1(\cpuregs[11][28] ),
    .A2(_20291_),
    .B1(_20492_),
    .C1(_20855_),
    .X(_20856_));
 sky130_fd_sc_hd__a21o_4 _27126_ (.A1(_20853_),
    .A2(_20856_),
    .B1(_20496_),
    .X(_20857_));
 sky130_fd_sc_hd__nand3_4 _27127_ (.A(_20850_),
    .B(_20857_),
    .C(_20498_),
    .Y(_20858_));
 sky130_fd_sc_hd__and2_4 _27128_ (.A(_20858_),
    .B(_19330_),
    .X(_20859_));
 sky130_fd_sc_hd__and2_4 _27129_ (.A(_19218_),
    .B(\cpuregs[0][28] ),
    .X(_20860_));
 sky130_fd_sc_hd__a211o_4 _27130_ (.A1(\cpuregs[1][28] ),
    .A2(_20298_),
    .B1(_20737_),
    .C1(_20860_),
    .X(_20861_));
 sky130_vsdinv _27131_ (.A(\cpuregs[2][28] ),
    .Y(_20862_));
 sky130_fd_sc_hd__nor2_4 _27132_ (.A(_20862_),
    .B(_20303_),
    .Y(_20863_));
 sky130_fd_sc_hd__a211o_4 _27133_ (.A1(\cpuregs[3][28] ),
    .A2(_19360_),
    .B1(_20301_),
    .C1(_20863_),
    .X(_20864_));
 sky130_fd_sc_hd__a21o_4 _27134_ (.A1(_20861_),
    .A2(_20864_),
    .B1(_19241_),
    .X(_20865_));
 sky130_vsdinv _27135_ (.A(\cpuregs[6][28] ),
    .Y(_20866_));
 sky130_fd_sc_hd__nor2_4 _27136_ (.A(_20866_),
    .B(_20309_),
    .Y(_20867_));
 sky130_fd_sc_hd__a211o_4 _27137_ (.A1(\cpuregs[7][28] ),
    .A2(_19620_),
    .B1(_20307_),
    .C1(_20867_),
    .X(_20868_));
 sky130_vsdinv _27138_ (.A(\cpuregs[4][28] ),
    .Y(_20869_));
 sky130_fd_sc_hd__nor2_4 _27139_ (.A(_20869_),
    .B(_20313_),
    .Y(_20870_));
 sky130_fd_sc_hd__a211o_4 _27140_ (.A1(\cpuregs[5][28] ),
    .A2(_20089_),
    .B1(_20611_),
    .C1(_20870_),
    .X(_20871_));
 sky130_fd_sc_hd__a21o_4 _27141_ (.A1(_20868_),
    .A2(_20871_),
    .B1(_19438_),
    .X(_20872_));
 sky130_fd_sc_hd__nand3_4 _27142_ (.A(_20865_),
    .B(_19255_),
    .C(_20872_),
    .Y(_20873_));
 sky130_fd_sc_hd__buf_1 _27143_ (.A(_20102_),
    .X(_20874_));
 sky130_fd_sc_hd__buf_1 _27144_ (.A(_20874_),
    .X(_20875_));
 sky130_vsdinv _27145_ (.A(\cpuregs[18][28] ),
    .Y(_20876_));
 sky130_fd_sc_hd__nor2_4 _27146_ (.A(_20876_),
    .B(_20518_),
    .Y(_20877_));
 sky130_fd_sc_hd__a211o_4 _27147_ (.A1(\cpuregs[19][28] ),
    .A2(_20516_),
    .B1(_19391_),
    .C1(_20877_),
    .X(_20878_));
 sky130_vsdinv _27148_ (.A(\cpuregs[16][28] ),
    .Y(_20879_));
 sky130_fd_sc_hd__nor2_4 _27149_ (.A(_20879_),
    .B(_19406_),
    .Y(_20880_));
 sky130_fd_sc_hd__a211o_4 _27150_ (.A1(\cpuregs[17][28] ),
    .A2(_19401_),
    .B1(_19402_),
    .C1(_20880_),
    .X(_20881_));
 sky130_fd_sc_hd__a21oi_4 _27151_ (.A1(_20878_),
    .A2(_20881_),
    .B1(_19410_),
    .Y(_20882_));
 sky130_fd_sc_hd__a2111o_4 _27152_ (.A1(_20859_),
    .A2(_20873_),
    .B1(_20785_),
    .C1(_20875_),
    .D1(_20882_),
    .X(_20883_));
 sky130_fd_sc_hd__buf_1 _27153_ (.A(\timer[28] ),
    .X(_20884_));
 sky130_fd_sc_hd__nand4_4 _27154_ (.A(_19414_),
    .B(_19416_),
    .C(_19417_),
    .D(_18931_),
    .Y(_20885_));
 sky130_fd_sc_hd__nor2_4 _27155_ (.A(_20884_),
    .B(_20885_),
    .Y(_20886_));
 sky130_vsdinv _27156_ (.A(_20886_),
    .Y(_20887_));
 sky130_fd_sc_hd__nand2_4 _27157_ (.A(_20885_),
    .B(_20884_),
    .Y(_20888_));
 sky130_fd_sc_hd__a21o_4 _27158_ (.A1(_20887_),
    .A2(_20888_),
    .B1(_20529_),
    .X(_20889_));
 sky130_fd_sc_hd__a21oi_4 _27159_ (.A1(_20883_),
    .A2(_20889_),
    .B1(_20798_),
    .Y(_00646_));
 sky130_fd_sc_hd__buf_1 _27160_ (.A(\timer[29] ),
    .X(_20890_));
 sky130_fd_sc_hd__nor4_4 _27161_ (.A(_20890_),
    .B(_20884_),
    .C(_18922_),
    .D(_20885_),
    .Y(_20891_));
 sky130_fd_sc_hd__a211o_4 _27162_ (.A1(_20890_),
    .A2(_20887_),
    .B1(_20381_),
    .C1(_20891_),
    .X(_20892_));
 sky130_vsdinv _27163_ (.A(\cpuregs[14][29] ),
    .Y(_20893_));
 sky130_fd_sc_hd__nor2_4 _27164_ (.A(_20893_),
    .B(_20181_),
    .Y(_20894_));
 sky130_fd_sc_hd__a211o_4 _27165_ (.A1(\cpuregs[15][29] ),
    .A2(_19497_),
    .B1(_20450_),
    .C1(_20894_),
    .X(_20895_));
 sky130_vsdinv _27166_ (.A(\cpuregs[12][29] ),
    .Y(_20896_));
 sky130_fd_sc_hd__nor2_4 _27167_ (.A(_20896_),
    .B(_19503_),
    .Y(_20897_));
 sky130_fd_sc_hd__a211o_4 _27168_ (.A1(\cpuregs[13][29] ),
    .A2(_20080_),
    .B1(_20812_),
    .C1(_20897_),
    .X(_20898_));
 sky130_fd_sc_hd__a21o_4 _27169_ (.A1(_20895_),
    .A2(_20898_),
    .B1(_19462_),
    .X(_20899_));
 sky130_vsdinv _27170_ (.A(\cpuregs[8][29] ),
    .Y(_20900_));
 sky130_fd_sc_hd__nor2_4 _27171_ (.A(_20900_),
    .B(_19404_),
    .Y(_20901_));
 sky130_fd_sc_hd__a211o_4 _27172_ (.A1(\cpuregs[9][29] ),
    .A2(_20188_),
    .B1(_19508_),
    .C1(_20901_),
    .X(_20902_));
 sky130_vsdinv _27173_ (.A(\cpuregs[10][29] ),
    .Y(_20903_));
 sky130_fd_sc_hd__nor2_4 _27174_ (.A(_20903_),
    .B(_20194_),
    .Y(_20904_));
 sky130_fd_sc_hd__a211o_4 _27175_ (.A1(\cpuregs[11][29] ),
    .A2(_19512_),
    .B1(_20192_),
    .C1(_20904_),
    .X(_20905_));
 sky130_fd_sc_hd__a21o_4 _27176_ (.A1(_20902_),
    .A2(_20905_),
    .B1(_19518_),
    .X(_20906_));
 sky130_fd_sc_hd__nand3_4 _27177_ (.A(_20899_),
    .B(_20906_),
    .C(_20198_),
    .Y(_20907_));
 sky130_fd_sc_hd__and2_4 _27178_ (.A(_20907_),
    .B(_20200_),
    .X(_20908_));
 sky130_fd_sc_hd__and2_4 _27179_ (.A(_20202_),
    .B(\cpuregs[0][29] ),
    .X(_20909_));
 sky130_fd_sc_hd__a211o_4 _27180_ (.A1(\cpuregs[1][29] ),
    .A2(_19631_),
    .B1(_19336_),
    .C1(_20909_),
    .X(_20910_));
 sky130_vsdinv _27181_ (.A(\cpuregs[2][29] ),
    .Y(_20911_));
 sky130_fd_sc_hd__nor2_4 _27182_ (.A(_20911_),
    .B(_19350_),
    .Y(_20912_));
 sky130_fd_sc_hd__a211o_4 _27183_ (.A1(\cpuregs[3][29] ),
    .A2(_19639_),
    .B1(_19787_),
    .C1(_20912_),
    .X(_20913_));
 sky130_fd_sc_hd__a21o_4 _27184_ (.A1(_20910_),
    .A2(_20913_),
    .B1(_19355_),
    .X(_20914_));
 sky130_vsdinv _27185_ (.A(\cpuregs[6][29] ),
    .Y(_20915_));
 sky130_fd_sc_hd__nor2_4 _27186_ (.A(_20915_),
    .B(_20259_),
    .Y(_20916_));
 sky130_fd_sc_hd__a211o_4 _27187_ (.A1(\cpuregs[7][29] ),
    .A2(_20209_),
    .B1(_20210_),
    .C1(_20916_),
    .X(_20917_));
 sky130_vsdinv _27188_ (.A(\cpuregs[4][29] ),
    .Y(_20918_));
 sky130_fd_sc_hd__nor2_4 _27189_ (.A(_20918_),
    .B(_19841_),
    .Y(_20919_));
 sky130_fd_sc_hd__a211o_4 _27190_ (.A1(\cpuregs[5][29] ),
    .A2(_19839_),
    .B1(_19621_),
    .C1(_20919_),
    .X(_20920_));
 sky130_fd_sc_hd__a21o_4 _27191_ (.A1(_20917_),
    .A2(_20920_),
    .B1(_19627_),
    .X(_20921_));
 sky130_fd_sc_hd__nand3_4 _27192_ (.A(_20914_),
    .B(_19616_),
    .C(_20921_),
    .Y(_20922_));
 sky130_vsdinv _27193_ (.A(\cpuregs[18][29] ),
    .Y(_20923_));
 sky130_fd_sc_hd__nor2_4 _27194_ (.A(_20923_),
    .B(_19636_),
    .Y(_20924_));
 sky130_fd_sc_hd__a211o_4 _27195_ (.A1(\cpuregs[19][29] ),
    .A2(_19632_),
    .B1(_19634_),
    .C1(_20924_),
    .X(_20925_));
 sky130_vsdinv _27196_ (.A(\cpuregs[16][29] ),
    .Y(_20926_));
 sky130_fd_sc_hd__nor2_4 _27197_ (.A(_20926_),
    .B(_19856_),
    .Y(_20927_));
 sky130_fd_sc_hd__a211o_4 _27198_ (.A1(\cpuregs[17][29] ),
    .A2(_19854_),
    .B1(_19641_),
    .C1(_20927_),
    .X(_20928_));
 sky130_fd_sc_hd__a21oi_4 _27199_ (.A1(_20925_),
    .A2(_20928_),
    .B1(_19647_),
    .Y(_20929_));
 sky130_fd_sc_hd__a211o_4 _27200_ (.A1(_20908_),
    .A2(_20922_),
    .B1(_20031_),
    .C1(_20929_),
    .X(_20930_));
 sky130_fd_sc_hd__nand2_4 _27201_ (.A(_20930_),
    .B(_20429_),
    .Y(_20931_));
 sky130_fd_sc_hd__buf_1 _27202_ (.A(_18861_),
    .X(_20932_));
 sky130_fd_sc_hd__and3_4 _27203_ (.A(_20892_),
    .B(_20931_),
    .C(_20932_),
    .X(_00647_));
 sky130_vsdinv _27204_ (.A(\cpuregs[14][30] ),
    .Y(_20933_));
 sky130_fd_sc_hd__nor2_4 _27205_ (.A(_20933_),
    .B(_19580_),
    .Y(_20934_));
 sky130_fd_sc_hd__a211o_4 _27206_ (.A1(\cpuregs[15][30] ),
    .A2(_20480_),
    .B1(_20034_),
    .C1(_20934_),
    .X(_20935_));
 sky130_vsdinv _27207_ (.A(\cpuregs[12][30] ),
    .Y(_20936_));
 sky130_fd_sc_hd__nor2_4 _27208_ (.A(_20936_),
    .B(_19292_),
    .Y(_20937_));
 sky130_fd_sc_hd__a211o_4 _27209_ (.A1(\cpuregs[13][30] ),
    .A2(_20484_),
    .B1(_20082_),
    .C1(_20937_),
    .X(_20938_));
 sky130_fd_sc_hd__a21o_4 _27210_ (.A1(_20935_),
    .A2(_20938_),
    .B1(_19306_),
    .X(_20939_));
 sky130_vsdinv _27211_ (.A(\cpuregs[8][30] ),
    .Y(_20940_));
 sky130_fd_sc_hd__nor2_4 _27212_ (.A(_20940_),
    .B(_19596_),
    .Y(_20941_));
 sky130_fd_sc_hd__a211o_4 _27213_ (.A1(\cpuregs[9][30] ),
    .A2(_19593_),
    .B1(_19299_),
    .C1(_20941_),
    .X(_20942_));
 sky130_vsdinv _27214_ (.A(\cpuregs[10][30] ),
    .Y(_20943_));
 sky130_fd_sc_hd__nor2_4 _27215_ (.A(_20943_),
    .B(_19730_),
    .Y(_20944_));
 sky130_fd_sc_hd__a211o_4 _27216_ (.A1(\cpuregs[11][30] ),
    .A2(_19310_),
    .B1(_20492_),
    .C1(_20944_),
    .X(_20945_));
 sky130_fd_sc_hd__a21o_4 _27217_ (.A1(_20942_),
    .A2(_20945_),
    .B1(_20496_),
    .X(_20946_));
 sky130_fd_sc_hd__nand3_4 _27218_ (.A(_20939_),
    .B(_20946_),
    .C(_20498_),
    .Y(_20947_));
 sky130_fd_sc_hd__and2_4 _27219_ (.A(_20947_),
    .B(_19330_),
    .X(_20948_));
 sky130_fd_sc_hd__and2_4 _27220_ (.A(_19218_),
    .B(\cpuregs[0][30] ),
    .X(_20949_));
 sky130_fd_sc_hd__a211o_4 _27221_ (.A1(\cpuregs[1][30] ),
    .A2(_19610_),
    .B1(_20737_),
    .C1(_20949_),
    .X(_20950_));
 sky130_vsdinv _27222_ (.A(\cpuregs[2][30] ),
    .Y(_20951_));
 sky130_fd_sc_hd__nor2_4 _27223_ (.A(_20951_),
    .B(_19363_),
    .Y(_20952_));
 sky130_fd_sc_hd__a211o_4 _27224_ (.A1(\cpuregs[3][30] ),
    .A2(_19360_),
    .B1(_19361_),
    .C1(_20952_),
    .X(_20953_));
 sky130_fd_sc_hd__a21o_4 _27225_ (.A1(_20950_),
    .A2(_20953_),
    .B1(_19241_),
    .X(_20954_));
 sky130_vsdinv _27226_ (.A(\cpuregs[6][30] ),
    .Y(_20955_));
 sky130_fd_sc_hd__nor2_4 _27227_ (.A(_20955_),
    .B(_19624_),
    .Y(_20956_));
 sky130_fd_sc_hd__a211o_4 _27228_ (.A1(\cpuregs[7][30] ),
    .A2(_19620_),
    .B1(_19390_),
    .C1(_20956_),
    .X(_20957_));
 sky130_vsdinv _27229_ (.A(\cpuregs[4][30] ),
    .Y(_20958_));
 sky130_fd_sc_hd__nor2_4 _27230_ (.A(_20958_),
    .B(_19258_),
    .Y(_20959_));
 sky130_fd_sc_hd__a211o_4 _27231_ (.A1(\cpuregs[5][30] ),
    .A2(_20089_),
    .B1(_20611_),
    .C1(_20959_),
    .X(_20960_));
 sky130_fd_sc_hd__a21o_4 _27232_ (.A1(_20957_),
    .A2(_20960_),
    .B1(_19438_),
    .X(_20961_));
 sky130_fd_sc_hd__nand3_4 _27233_ (.A(_20954_),
    .B(_19255_),
    .C(_20961_),
    .Y(_20962_));
 sky130_vsdinv _27234_ (.A(\cpuregs[18][30] ),
    .Y(_20963_));
 sky130_fd_sc_hd__nor2_4 _27235_ (.A(_20963_),
    .B(_20518_),
    .Y(_20964_));
 sky130_fd_sc_hd__a211o_4 _27236_ (.A1(\cpuregs[19][30] ),
    .A2(_20516_),
    .B1(_19391_),
    .C1(_20964_),
    .X(_20965_));
 sky130_vsdinv _27237_ (.A(\cpuregs[16][30] ),
    .Y(_20966_));
 sky130_fd_sc_hd__nor2_4 _27238_ (.A(_20966_),
    .B(_19406_),
    .Y(_20967_));
 sky130_fd_sc_hd__a211o_4 _27239_ (.A1(\cpuregs[17][30] ),
    .A2(_19401_),
    .B1(_19402_),
    .C1(_20967_),
    .X(_20968_));
 sky130_fd_sc_hd__a21oi_4 _27240_ (.A1(_20965_),
    .A2(_20968_),
    .B1(_19410_),
    .Y(_20969_));
 sky130_fd_sc_hd__a2111o_4 _27241_ (.A1(_20948_),
    .A2(_20962_),
    .B1(_20785_),
    .C1(_20875_),
    .D1(_20969_),
    .X(_20970_));
 sky130_fd_sc_hd__nor2_4 _27242_ (.A(_20890_),
    .B(\timer[28] ),
    .Y(_20971_));
 sky130_vsdinv _27243_ (.A(\timer[30] ),
    .Y(_20972_));
 sky130_fd_sc_hd__a41oi_4 _27244_ (.A1(_20330_),
    .A2(_20233_),
    .A3(_20971_),
    .A4(_18931_),
    .B1(_20972_),
    .Y(_20973_));
 sky130_fd_sc_hd__and4_4 _27245_ (.A(_20378_),
    .B(_20972_),
    .C(_20971_),
    .D(_18931_),
    .X(_20974_));
 sky130_fd_sc_hd__o21ai_4 _27246_ (.A1(_20973_),
    .A2(_20974_),
    .B1(_19420_),
    .Y(_20975_));
 sky130_fd_sc_hd__a21oi_4 _27247_ (.A1(_20970_),
    .A2(_20975_),
    .B1(_20798_),
    .Y(_00649_));
 sky130_vsdinv _27248_ (.A(\cpuregs[14][31] ),
    .Y(_20976_));
 sky130_fd_sc_hd__nor2_4 _27249_ (.A(_20976_),
    .B(_19574_),
    .Y(_20977_));
 sky130_fd_sc_hd__a211o_4 _27250_ (.A1(\cpuregs[15][31] ),
    .A2(_19468_),
    .B1(_19571_),
    .C1(_20977_),
    .X(_20978_));
 sky130_vsdinv _27251_ (.A(\cpuregs[12][31] ),
    .Y(_20979_));
 sky130_fd_sc_hd__nor2_4 _27252_ (.A(_20979_),
    .B(_19429_),
    .Y(_20980_));
 sky130_fd_sc_hd__a211o_4 _27253_ (.A1(\cpuregs[13][31] ),
    .A2(_19804_),
    .B1(_19578_),
    .C1(_20980_),
    .X(_20981_));
 sky130_fd_sc_hd__a21o_4 _27254_ (.A1(_20978_),
    .A2(_20981_),
    .B1(_19584_),
    .X(_20982_));
 sky130_vsdinv _27255_ (.A(\cpuregs[8][31] ),
    .Y(_20983_));
 sky130_fd_sc_hd__nor2_4 _27256_ (.A(_20983_),
    .B(_19433_),
    .Y(_20984_));
 sky130_fd_sc_hd__a211o_4 _27257_ (.A1(\cpuregs[9][31] ),
    .A2(_19586_),
    .B1(_20812_),
    .C1(_20984_),
    .X(_20985_));
 sky130_vsdinv _27258_ (.A(\cpuregs[10][31] ),
    .Y(_20986_));
 sky130_fd_sc_hd__nor2_4 _27259_ (.A(_20986_),
    .B(_19819_),
    .Y(_20987_));
 sky130_fd_sc_hd__a211o_4 _27260_ (.A1(\cpuregs[11][31] ),
    .A2(_19507_),
    .B1(_19594_),
    .C1(_20987_),
    .X(_20988_));
 sky130_fd_sc_hd__a21o_4 _27261_ (.A1(_20985_),
    .A2(_20988_),
    .B1(_19354_),
    .X(_20989_));
 sky130_fd_sc_hd__nand3_4 _27262_ (.A(_20982_),
    .B(_20989_),
    .C(_19601_),
    .Y(_20990_));
 sky130_fd_sc_hd__and2_4 _27263_ (.A(_20990_),
    .B(_19603_),
    .X(_20991_));
 sky130_fd_sc_hd__and2_4 _27264_ (.A(_19338_),
    .B(\cpuregs[0][31] ),
    .X(_20992_));
 sky130_fd_sc_hd__a211o_4 _27265_ (.A1(\cpuregs[1][31] ),
    .A2(_19335_),
    .B1(_19606_),
    .C1(_20992_),
    .X(_20993_));
 sky130_vsdinv _27266_ (.A(\cpuregs[2][31] ),
    .Y(_20994_));
 sky130_fd_sc_hd__nor2_4 _27267_ (.A(_20994_),
    .B(_19350_),
    .Y(_20995_));
 sky130_fd_sc_hd__a211o_4 _27268_ (.A1(\cpuregs[3][31] ),
    .A2(_19343_),
    .B1(_19346_),
    .C1(_20995_),
    .X(_20996_));
 sky130_fd_sc_hd__a21o_4 _27269_ (.A1(_20993_),
    .A2(_20996_),
    .B1(_19355_),
    .X(_20997_));
 sky130_vsdinv _27270_ (.A(\cpuregs[6][31] ),
    .Y(_20998_));
 sky130_fd_sc_hd__nor2_4 _27271_ (.A(_20998_),
    .B(_19536_),
    .Y(_20999_));
 sky130_fd_sc_hd__a211o_4 _27272_ (.A1(\cpuregs[7][31] ),
    .A2(_19532_),
    .B1(_19534_),
    .C1(_20999_),
    .X(_21000_));
 sky130_vsdinv _27273_ (.A(\cpuregs[4][31] ),
    .Y(_21001_));
 sky130_fd_sc_hd__nor2_4 _27274_ (.A(_21001_),
    .B(_19841_),
    .Y(_21002_));
 sky130_fd_sc_hd__a211o_4 _27275_ (.A1(\cpuregs[5][31] ),
    .A2(_19839_),
    .B1(_19621_),
    .C1(_21002_),
    .X(_21003_));
 sky130_fd_sc_hd__a21o_4 _27276_ (.A1(_21000_),
    .A2(_21003_),
    .B1(_19627_),
    .X(_21004_));
 sky130_fd_sc_hd__nand3_4 _27277_ (.A(_20997_),
    .B(_19616_),
    .C(_21004_),
    .Y(_21005_));
 sky130_vsdinv _27278_ (.A(\cpuregs[18][31] ),
    .Y(_21006_));
 sky130_fd_sc_hd__nor2_4 _27279_ (.A(_21006_),
    .B(_20045_),
    .Y(_21007_));
 sky130_fd_sc_hd__a211o_4 _27280_ (.A1(\cpuregs[19][31] ),
    .A2(_20041_),
    .B1(_19788_),
    .C1(_21007_),
    .X(_21008_));
 sky130_vsdinv _27281_ (.A(\cpuregs[16][31] ),
    .Y(_21009_));
 sky130_fd_sc_hd__nor2_4 _27282_ (.A(_21009_),
    .B(_19396_),
    .Y(_21010_));
 sky130_fd_sc_hd__a211o_4 _27283_ (.A1(\cpuregs[17][31] ),
    .A2(_19388_),
    .B1(_19792_),
    .C1(_21010_),
    .X(_21011_));
 sky130_fd_sc_hd__a21oi_4 _27284_ (.A1(_21008_),
    .A2(_21011_),
    .B1(_19796_),
    .Y(_21012_));
 sky130_fd_sc_hd__a2111o_4 _27285_ (.A1(_20991_),
    .A2(_21005_),
    .B1(_20785_),
    .C1(_20875_),
    .D1(_21012_),
    .X(_21013_));
 sky130_vsdinv _27286_ (.A(_20974_),
    .Y(_21014_));
 sky130_fd_sc_hd__nand3_4 _27287_ (.A(_21014_),
    .B(\timer[31] ),
    .C(_19166_),
    .Y(_21015_));
 sky130_fd_sc_hd__a21oi_4 _27288_ (.A1(_21013_),
    .A2(_21015_),
    .B1(_20798_),
    .Y(_00650_));
 sky130_fd_sc_hd__buf_1 _27289_ (.A(instr_maskirq),
    .X(_21016_));
 sky130_fd_sc_hd__nand2_4 _27290_ (.A(_21016_),
    .B(_20230_),
    .Y(_21017_));
 sky130_fd_sc_hd__buf_1 _27291_ (.A(_21017_),
    .X(_21018_));
 sky130_fd_sc_hd__buf_1 _27292_ (.A(_21018_),
    .X(_21019_));
 sky130_fd_sc_hd__buf_1 _27293_ (.A(_21017_),
    .X(_21020_));
 sky130_fd_sc_hd__buf_1 _27294_ (.A(_21020_),
    .X(_21021_));
 sky130_fd_sc_hd__buf_1 _27295_ (.A(_18264_),
    .X(_21022_));
 sky130_fd_sc_hd__buf_1 _27296_ (.A(_21022_),
    .X(_21023_));
 sky130_fd_sc_hd__a21oi_4 _27297_ (.A1(_21021_),
    .A2(\irq_mask[0] ),
    .B1(_21023_),
    .Y(_21024_));
 sky130_fd_sc_hd__o41ai_4 _27298_ (.A1(_19281_),
    .A2(_19384_),
    .A3(_19226_),
    .A4(_21019_),
    .B1(_21024_),
    .Y(_00296_));
 sky130_fd_sc_hd__a2111o_4 _27299_ (.A1(_19332_),
    .A2(_19379_),
    .B1(_20157_),
    .C1(_19412_),
    .D1(_21020_),
    .X(_21025_));
 sky130_vsdinv _27300_ (.A(_21025_),
    .Y(_21026_));
 sky130_fd_sc_hd__a211o_4 _27301_ (.A1(\irq_mask[1] ),
    .A2(_21019_),
    .B1(_18286_),
    .C1(_21026_),
    .X(_00307_));
 sky130_fd_sc_hd__buf_1 _27302_ (.A(_21021_),
    .X(_21027_));
 sky130_fd_sc_hd__buf_1 _27303_ (.A(_20156_),
    .X(_21028_));
 sky130_fd_sc_hd__a211o_4 _27304_ (.A1(_19450_),
    .A2(_19478_),
    .B1(_21028_),
    .C1(_19489_),
    .X(_21029_));
 sky130_fd_sc_hd__buf_1 _27305_ (.A(_21018_),
    .X(_21030_));
 sky130_fd_sc_hd__buf_1 _27306_ (.A(_21022_),
    .X(_21031_));
 sky130_fd_sc_hd__a21oi_4 _27307_ (.A1(_21030_),
    .A2(_18311_),
    .B1(_21031_),
    .Y(_21032_));
 sky130_fd_sc_hd__o21ai_4 _27308_ (.A1(_21027_),
    .A2(_21029_),
    .B1(_21032_),
    .Y(_00318_));
 sky130_fd_sc_hd__a211o_4 _27309_ (.A1(_19523_),
    .A2(_19551_),
    .B1(_21028_),
    .C1(_19562_),
    .X(_21033_));
 sky130_fd_sc_hd__a21oi_4 _27310_ (.A1(_21030_),
    .A2(\irq_mask[3] ),
    .B1(_21031_),
    .Y(_21034_));
 sky130_fd_sc_hd__o21ai_4 _27311_ (.A1(_21027_),
    .A2(_21033_),
    .B1(_21034_),
    .Y(_00321_));
 sky130_fd_sc_hd__a211o_4 _27312_ (.A1(_19604_),
    .A2(_19629_),
    .B1(_21028_),
    .C1(_19648_),
    .X(_21035_));
 sky130_fd_sc_hd__a21oi_4 _27313_ (.A1(_21030_),
    .A2(\irq_mask[4] ),
    .B1(_21031_),
    .Y(_21036_));
 sky130_fd_sc_hd__o21ai_4 _27314_ (.A1(_21027_),
    .A2(_21035_),
    .B1(_21036_),
    .Y(_00322_));
 sky130_fd_sc_hd__buf_1 _27315_ (.A(_20649_),
    .X(_21037_));
 sky130_fd_sc_hd__a211o_4 _27316_ (.A1(_19671_),
    .A2(_19686_),
    .B1(_21037_),
    .C1(_19693_),
    .X(_21038_));
 sky130_fd_sc_hd__buf_1 _27317_ (.A(_18264_),
    .X(_21039_));
 sky130_fd_sc_hd__buf_1 _27318_ (.A(_21039_),
    .X(_21040_));
 sky130_fd_sc_hd__a21oi_4 _27319_ (.A1(_21030_),
    .A2(\irq_mask[5] ),
    .B1(_21040_),
    .Y(_21041_));
 sky130_fd_sc_hd__o21ai_4 _27320_ (.A1(_21027_),
    .A2(_21038_),
    .B1(_21041_),
    .Y(_00323_));
 sky130_fd_sc_hd__buf_1 _27321_ (.A(_21020_),
    .X(_21042_));
 sky130_fd_sc_hd__buf_1 _27322_ (.A(_21042_),
    .X(_21043_));
 sky130_fd_sc_hd__a211o_4 _27323_ (.A1(_19719_),
    .A2(_19738_),
    .B1(_21037_),
    .C1(_19749_),
    .X(_21044_));
 sky130_fd_sc_hd__buf_1 _27324_ (.A(_21018_),
    .X(_21045_));
 sky130_fd_sc_hd__a21oi_4 _27325_ (.A1(_21045_),
    .A2(\irq_mask[6] ),
    .B1(_21040_),
    .Y(_21046_));
 sky130_fd_sc_hd__o21ai_4 _27326_ (.A1(_21043_),
    .A2(_21044_),
    .B1(_21046_),
    .Y(_00324_));
 sky130_fd_sc_hd__a211o_4 _27327_ (.A1(_19770_),
    .A2(_19785_),
    .B1(_21037_),
    .C1(_19797_),
    .X(_21047_));
 sky130_fd_sc_hd__a21oi_4 _27328_ (.A1(_21045_),
    .A2(\irq_mask[7] ),
    .B1(_21040_),
    .Y(_21048_));
 sky130_fd_sc_hd__o21ai_4 _27329_ (.A1(_21043_),
    .A2(_21047_),
    .B1(_21048_),
    .Y(_00325_));
 sky130_fd_sc_hd__a211o_4 _27330_ (.A1(_19829_),
    .A2(_19853_),
    .B1(_21037_),
    .C1(_19862_),
    .X(_21049_));
 sky130_fd_sc_hd__a21oi_4 _27331_ (.A1(_21045_),
    .A2(\irq_mask[8] ),
    .B1(_21040_),
    .Y(_21050_));
 sky130_fd_sc_hd__o21ai_4 _27332_ (.A1(_21043_),
    .A2(_21049_),
    .B1(_21050_),
    .Y(_00326_));
 sky130_fd_sc_hd__buf_1 _27333_ (.A(_20103_),
    .X(_21051_));
 sky130_fd_sc_hd__a211o_4 _27334_ (.A1(_19888_),
    .A2(_19907_),
    .B1(_21051_),
    .C1(_19919_),
    .X(_21052_));
 sky130_fd_sc_hd__buf_1 _27335_ (.A(_21039_),
    .X(_21053_));
 sky130_fd_sc_hd__a21oi_4 _27336_ (.A1(_21045_),
    .A2(\irq_mask[9] ),
    .B1(_21053_),
    .Y(_21054_));
 sky130_fd_sc_hd__o21ai_4 _27337_ (.A1(_21043_),
    .A2(_21052_),
    .B1(_21054_),
    .Y(_00327_));
 sky130_fd_sc_hd__buf_1 _27338_ (.A(_21020_),
    .X(_21055_));
 sky130_fd_sc_hd__buf_1 _27339_ (.A(_18264_),
    .X(_21056_));
 sky130_fd_sc_hd__buf_1 _27340_ (.A(_21056_),
    .X(_21057_));
 sky130_fd_sc_hd__buf_1 _27341_ (.A(_21016_),
    .X(_21058_));
 sky130_fd_sc_hd__buf_1 _27342_ (.A(_21058_),
    .X(_21059_));
 sky130_fd_sc_hd__buf_1 _27343_ (.A(_21059_),
    .X(_21060_));
 sky130_fd_sc_hd__buf_1 _27344_ (.A(_18798_),
    .X(_21061_));
 sky130_fd_sc_hd__nand4_4 _27345_ (.A(_21060_),
    .B(_19965_),
    .C(_21061_),
    .D(_19974_),
    .Y(_21062_));
 sky130_vsdinv _27346_ (.A(_21062_),
    .Y(_21063_));
 sky130_fd_sc_hd__a211o_4 _27347_ (.A1(\irq_mask[10] ),
    .A2(_21055_),
    .B1(_21057_),
    .C1(_21063_),
    .X(_00297_));
 sky130_fd_sc_hd__buf_1 _27348_ (.A(_21042_),
    .X(_21064_));
 sky130_fd_sc_hd__buf_1 _27349_ (.A(_21017_),
    .X(_21065_));
 sky130_fd_sc_hd__buf_1 _27350_ (.A(_21065_),
    .X(_21066_));
 sky130_fd_sc_hd__a21oi_4 _27351_ (.A1(_21066_),
    .A2(\irq_mask[11] ),
    .B1(_21053_),
    .Y(_21067_));
 sky130_fd_sc_hd__o21ai_4 _27352_ (.A1(_21064_),
    .A2(_20050_),
    .B1(_21067_),
    .Y(_00298_));
 sky130_fd_sc_hd__a21oi_4 _27353_ (.A1(_21066_),
    .A2(\irq_mask[12] ),
    .B1(_21053_),
    .Y(_21068_));
 sky130_fd_sc_hd__o21ai_4 _27354_ (.A1(_21064_),
    .A2(_20111_),
    .B1(_21068_),
    .Y(_00299_));
 sky130_fd_sc_hd__a21oi_4 _27355_ (.A1(_21066_),
    .A2(\irq_mask[13] ),
    .B1(_21053_),
    .Y(_21069_));
 sky130_fd_sc_hd__o21ai_4 _27356_ (.A1(_21064_),
    .A2(_20170_),
    .B1(_21069_),
    .Y(_00300_));
 sky130_fd_sc_hd__buf_1 _27357_ (.A(_21039_),
    .X(_21070_));
 sky130_fd_sc_hd__a21oi_4 _27358_ (.A1(_21066_),
    .A2(\irq_mask[14] ),
    .B1(_21070_),
    .Y(_21071_));
 sky130_fd_sc_hd__o21ai_4 _27359_ (.A1(_21064_),
    .A2(_20226_),
    .B1(_21071_),
    .Y(_00301_));
 sky130_fd_sc_hd__buf_1 _27360_ (.A(_21042_),
    .X(_21072_));
 sky130_fd_sc_hd__buf_1 _27361_ (.A(_21065_),
    .X(_21073_));
 sky130_fd_sc_hd__a21oi_4 _27362_ (.A1(_21073_),
    .A2(\irq_mask[15] ),
    .B1(_21070_),
    .Y(_21074_));
 sky130_fd_sc_hd__o21ai_4 _27363_ (.A1(_21072_),
    .A2(_20275_),
    .B1(_21074_),
    .Y(_00302_));
 sky130_fd_sc_hd__buf_1 _27364_ (.A(_20649_),
    .X(_21075_));
 sky130_fd_sc_hd__a211o_4 _27365_ (.A1(_20297_),
    .A2(_20317_),
    .B1(_21075_),
    .C1(_20325_),
    .X(_21076_));
 sky130_fd_sc_hd__a21oi_4 _27366_ (.A1(_21073_),
    .A2(\irq_mask[16] ),
    .B1(_21070_),
    .Y(_21077_));
 sky130_fd_sc_hd__o21ai_4 _27367_ (.A1(_21072_),
    .A2(_21076_),
    .B1(_21077_),
    .Y(_00303_));
 sky130_fd_sc_hd__a21oi_4 _27368_ (.A1(_21073_),
    .A2(\irq_mask[17] ),
    .B1(_21070_),
    .Y(_21078_));
 sky130_fd_sc_hd__o21ai_4 _27369_ (.A1(_21072_),
    .A2(_20374_),
    .B1(_21078_),
    .Y(_00304_));
 sky130_fd_sc_hd__buf_1 _27370_ (.A(_21039_),
    .X(_21079_));
 sky130_fd_sc_hd__a21oi_4 _27371_ (.A1(_21073_),
    .A2(\irq_mask[18] ),
    .B1(_21079_),
    .Y(_21080_));
 sky130_fd_sc_hd__o21ai_4 _27372_ (.A1(_21072_),
    .A2(_20428_),
    .B1(_21080_),
    .Y(_00305_));
 sky130_fd_sc_hd__buf_1 _27373_ (.A(_21042_),
    .X(_21081_));
 sky130_fd_sc_hd__buf_1 _27374_ (.A(_21065_),
    .X(_21082_));
 sky130_fd_sc_hd__a21oi_4 _27375_ (.A1(_21082_),
    .A2(\irq_mask[19] ),
    .B1(_21079_),
    .Y(_21083_));
 sky130_fd_sc_hd__o21ai_4 _27376_ (.A1(_21081_),
    .A2(_20478_),
    .B1(_21083_),
    .Y(_00306_));
 sky130_fd_sc_hd__a211o_4 _27377_ (.A1(_20500_),
    .A2(_20514_),
    .B1(_21075_),
    .C1(_20524_),
    .X(_21084_));
 sky130_fd_sc_hd__a21oi_4 _27378_ (.A1(_21082_),
    .A2(\irq_mask[20] ),
    .B1(_21079_),
    .Y(_21085_));
 sky130_fd_sc_hd__o21ai_4 _27379_ (.A1(_21081_),
    .A2(_21084_),
    .B1(_21085_),
    .Y(_00308_));
 sky130_fd_sc_hd__a21oi_4 _27380_ (.A1(_21082_),
    .A2(\irq_mask[21] ),
    .B1(_21079_),
    .Y(_21086_));
 sky130_fd_sc_hd__o21ai_4 _27381_ (.A1(_21081_),
    .A2(_20573_),
    .B1(_21086_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand4_4 _27382_ (.A(_21060_),
    .B(_20607_),
    .C(_21061_),
    .D(_20616_),
    .Y(_21087_));
 sky130_vsdinv _27383_ (.A(_21087_),
    .Y(_21088_));
 sky130_fd_sc_hd__a211o_4 _27384_ (.A1(\irq_mask[22] ),
    .A2(_21055_),
    .B1(_21057_),
    .C1(_21088_),
    .X(_00310_));
 sky130_fd_sc_hd__buf_1 _27385_ (.A(_21022_),
    .X(_21089_));
 sky130_fd_sc_hd__a21oi_4 _27386_ (.A1(_21082_),
    .A2(\irq_mask[23] ),
    .B1(_21089_),
    .Y(_21090_));
 sky130_fd_sc_hd__o21ai_4 _27387_ (.A1(_21081_),
    .A2(_20657_),
    .B1(_21090_),
    .Y(_00311_));
 sky130_fd_sc_hd__a2111o_4 _27388_ (.A1(_20680_),
    .A2(_20695_),
    .B1(_20157_),
    .C1(_20703_),
    .D1(_21017_),
    .X(_21091_));
 sky130_vsdinv _27389_ (.A(_21091_),
    .Y(_21092_));
 sky130_fd_sc_hd__a211o_4 _27390_ (.A1(\irq_mask[24] ),
    .A2(_21055_),
    .B1(_21057_),
    .C1(_21092_),
    .X(_00312_));
 sky130_fd_sc_hd__buf_1 _27391_ (.A(_21018_),
    .X(_21093_));
 sky130_fd_sc_hd__a211o_4 _27392_ (.A1(_20727_),
    .A2(_20742_),
    .B1(_21051_),
    .C1(_20749_),
    .X(_21094_));
 sky130_fd_sc_hd__buf_1 _27393_ (.A(_21065_),
    .X(_21095_));
 sky130_fd_sc_hd__a21oi_4 _27394_ (.A1(_21095_),
    .A2(\irq_mask[25] ),
    .B1(_21089_),
    .Y(_21096_));
 sky130_fd_sc_hd__o21ai_4 _27395_ (.A1(_21093_),
    .A2(_21094_),
    .B1(_21096_),
    .Y(_00313_));
 sky130_fd_sc_hd__a211o_4 _27396_ (.A1(_20770_),
    .A2(_20784_),
    .B1(_21051_),
    .C1(_20792_),
    .X(_21097_));
 sky130_fd_sc_hd__a21oi_4 _27397_ (.A1(_21095_),
    .A2(\irq_mask[26] ),
    .B1(_21089_),
    .Y(_21098_));
 sky130_fd_sc_hd__o21ai_4 _27398_ (.A1(_21093_),
    .A2(_21097_),
    .B1(_21098_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand4_4 _27399_ (.A(_21060_),
    .B(_20833_),
    .C(_21061_),
    .D(_20841_),
    .Y(_21099_));
 sky130_vsdinv _27400_ (.A(_21099_),
    .Y(_21100_));
 sky130_fd_sc_hd__a211o_4 _27401_ (.A1(\irq_mask[27] ),
    .A2(_21055_),
    .B1(_21057_),
    .C1(_21100_),
    .X(_00315_));
 sky130_fd_sc_hd__a211o_4 _27402_ (.A1(_20859_),
    .A2(_20873_),
    .B1(_21075_),
    .C1(_20882_),
    .X(_21101_));
 sky130_fd_sc_hd__a21oi_4 _27403_ (.A1(_21095_),
    .A2(\irq_mask[28] ),
    .B1(_21089_),
    .Y(_21102_));
 sky130_fd_sc_hd__o21ai_4 _27404_ (.A1(_21093_),
    .A2(_21101_),
    .B1(_21102_),
    .Y(_00316_));
 sky130_fd_sc_hd__a21oi_4 _27405_ (.A1(_21095_),
    .A2(\irq_mask[29] ),
    .B1(_21023_),
    .Y(_21103_));
 sky130_fd_sc_hd__o21ai_4 _27406_ (.A1(_21093_),
    .A2(_20930_),
    .B1(_21103_),
    .Y(_00317_));
 sky130_fd_sc_hd__a211o_4 _27407_ (.A1(_20948_),
    .A2(_20962_),
    .B1(_21075_),
    .C1(_20969_),
    .X(_21104_));
 sky130_fd_sc_hd__a21oi_4 _27408_ (.A1(_21021_),
    .A2(\irq_mask[30] ),
    .B1(_21023_),
    .Y(_21105_));
 sky130_fd_sc_hd__o21ai_4 _27409_ (.A1(_21019_),
    .A2(_21104_),
    .B1(_21105_),
    .Y(_00319_));
 sky130_fd_sc_hd__a211o_4 _27410_ (.A1(_20991_),
    .A2(_21005_),
    .B1(_21051_),
    .C1(_21012_),
    .X(_21106_));
 sky130_fd_sc_hd__a21oi_4 _27411_ (.A1(_21021_),
    .A2(\irq_mask[31] ),
    .B1(_21023_),
    .Y(_21107_));
 sky130_fd_sc_hd__o21ai_4 _27412_ (.A1(_21019_),
    .A2(_21106_),
    .B1(_21107_),
    .Y(_00320_));
 sky130_vsdinv _27413_ (.A(mem_la_wdata[0]),
    .Y(_21108_));
 sky130_fd_sc_hd__buf_1 _27414_ (.A(_21108_),
    .X(_21109_));
 sky130_fd_sc_hd__buf_1 _27415_ (.A(_21109_),
    .X(_21110_));
 sky130_fd_sc_hd__o21a_4 _27416_ (.A1(_20230_),
    .A2(_18534_),
    .B1(_18248_),
    .X(_21111_));
 sky130_fd_sc_hd__buf_1 _27417_ (.A(_21111_),
    .X(_21112_));
 sky130_fd_sc_hd__buf_1 _27418_ (.A(_21112_),
    .X(_21113_));
 sky130_fd_sc_hd__buf_1 _27419_ (.A(is_slli_srli_srai),
    .X(_21114_));
 sky130_fd_sc_hd__buf_1 _27420_ (.A(_18289_),
    .X(_21115_));
 sky130_fd_sc_hd__buf_1 _27421_ (.A(_21115_),
    .X(_21116_));
 sky130_fd_sc_hd__buf_1 _27422_ (.A(is_slli_srli_srai),
    .X(_21117_));
 sky130_fd_sc_hd__buf_1 _27423_ (.A(\decoded_imm[0] ),
    .X(_21118_));
 sky130_fd_sc_hd__nor2_4 _27424_ (.A(_21117_),
    .B(_21118_),
    .Y(_21119_));
 sky130_fd_sc_hd__a211o_4 _27425_ (.A1(_19167_),
    .A2(_21114_),
    .B1(_21116_),
    .C1(_21119_),
    .X(_21120_));
 sky130_fd_sc_hd__o41ai_4 _27426_ (.A1(_18806_),
    .A2(_19384_),
    .A3(_19226_),
    .A4(_19281_),
    .B1(_21120_),
    .Y(_21121_));
 sky130_fd_sc_hd__a2bb2o_4 _27427_ (.A1_N(_21110_),
    .A2_N(_21113_),
    .B1(_19112_),
    .B2(_21121_),
    .X(_00562_));
 sky130_vsdinv _27428_ (.A(mem_la_wdata[1]),
    .Y(_21122_));
 sky130_fd_sc_hd__buf_1 _27429_ (.A(_21122_),
    .X(_21123_));
 sky130_fd_sc_hd__buf_1 _27430_ (.A(_21123_),
    .X(_21124_));
 sky130_fd_sc_hd__buf_1 _27431_ (.A(_21124_),
    .X(_21125_));
 sky130_fd_sc_hd__buf_1 _27432_ (.A(_21125_),
    .X(_21126_));
 sky130_fd_sc_hd__buf_1 _27433_ (.A(_21126_),
    .X(_21127_));
 sky130_fd_sc_hd__buf_1 _27434_ (.A(_19124_),
    .X(_21128_));
 sky130_fd_sc_hd__buf_1 _27435_ (.A(_21128_),
    .X(_21129_));
 sky130_fd_sc_hd__buf_1 _27436_ (.A(_18787_),
    .X(_21130_));
 sky130_fd_sc_hd__a2111o_4 _27437_ (.A1(_19332_),
    .A2(_19379_),
    .B1(_21130_),
    .C1(_20875_),
    .D1(_19412_),
    .X(_21131_));
 sky130_fd_sc_hd__buf_1 _27438_ (.A(_21117_),
    .X(_21132_));
 sky130_fd_sc_hd__buf_1 _27439_ (.A(_18290_),
    .X(_21133_));
 sky130_fd_sc_hd__buf_1 _27440_ (.A(_21133_),
    .X(_21134_));
 sky130_fd_sc_hd__buf_1 _27441_ (.A(\decoded_imm[1] ),
    .X(_21135_));
 sky130_fd_sc_hd__nor2_4 _27442_ (.A(_21117_),
    .B(_21135_),
    .Y(_21136_));
 sky130_fd_sc_hd__a211o_4 _27443_ (.A1(_19178_),
    .A2(_21132_),
    .B1(_21134_),
    .C1(_21136_),
    .X(_21137_));
 sky130_fd_sc_hd__nand2_4 _27444_ (.A(_21131_),
    .B(_21137_),
    .Y(_21138_));
 sky130_fd_sc_hd__a2bb2o_4 _27445_ (.A1_N(_21127_),
    .A2_N(_21113_),
    .B1(_21129_),
    .B2(_21138_),
    .X(_00573_));
 sky130_vsdinv _27446_ (.A(mem_la_wdata[2]),
    .Y(_21139_));
 sky130_fd_sc_hd__buf_1 _27447_ (.A(_21139_),
    .X(_21140_));
 sky130_fd_sc_hd__buf_1 _27448_ (.A(_21140_),
    .X(_21141_));
 sky130_fd_sc_hd__buf_1 _27449_ (.A(_21141_),
    .X(_21142_));
 sky130_fd_sc_hd__buf_1 _27450_ (.A(_21142_),
    .X(_21143_));
 sky130_fd_sc_hd__buf_1 _27451_ (.A(_21143_),
    .X(_21144_));
 sky130_fd_sc_hd__buf_1 _27452_ (.A(_21144_),
    .X(_21145_));
 sky130_fd_sc_hd__buf_1 _27453_ (.A(_18806_),
    .X(_21146_));
 sky130_fd_sc_hd__buf_1 _27454_ (.A(\decoded_imm[2] ),
    .X(_21147_));
 sky130_fd_sc_hd__nor2_4 _27455_ (.A(_21117_),
    .B(_21147_),
    .Y(_21148_));
 sky130_fd_sc_hd__a211o_4 _27456_ (.A1(_19173_),
    .A2(_21114_),
    .B1(_21134_),
    .C1(_21148_),
    .X(_21149_));
 sky130_fd_sc_hd__o21ai_4 _27457_ (.A1(_21146_),
    .A2(_21029_),
    .B1(_21149_),
    .Y(_21150_));
 sky130_fd_sc_hd__a2bb2o_4 _27458_ (.A1_N(_21145_),
    .A2_N(_21113_),
    .B1(_21129_),
    .B2(_21150_),
    .X(_00584_));
 sky130_vsdinv _27459_ (.A(mem_la_wdata[3]),
    .Y(_21151_));
 sky130_fd_sc_hd__buf_1 _27460_ (.A(_21151_),
    .X(_21152_));
 sky130_fd_sc_hd__buf_1 _27461_ (.A(_21152_),
    .X(_21153_));
 sky130_fd_sc_hd__buf_1 _27462_ (.A(_21153_),
    .X(_21154_));
 sky130_fd_sc_hd__buf_1 _27463_ (.A(_21154_),
    .X(_21155_));
 sky130_fd_sc_hd__buf_1 _27464_ (.A(_21155_),
    .X(_21156_));
 sky130_vsdinv _27465_ (.A(is_slli_srli_srai),
    .Y(_21157_));
 sky130_fd_sc_hd__buf_1 _27466_ (.A(_21157_),
    .X(_21158_));
 sky130_fd_sc_hd__buf_1 _27467_ (.A(\decoded_imm[3] ),
    .X(_21159_));
 sky130_vsdinv _27468_ (.A(_21159_),
    .Y(_21160_));
 sky130_fd_sc_hd__buf_1 _27469_ (.A(_21157_),
    .X(_21161_));
 sky130_fd_sc_hd__nor2_4 _27470_ (.A(\decoded_rs2[3] ),
    .B(_21161_),
    .Y(_21162_));
 sky130_fd_sc_hd__a211o_4 _27471_ (.A1(_21158_),
    .A2(_21160_),
    .B1(_21134_),
    .C1(_21162_),
    .X(_21163_));
 sky130_fd_sc_hd__o21ai_4 _27472_ (.A1(_21146_),
    .A2(_21033_),
    .B1(_21163_),
    .Y(_21164_));
 sky130_fd_sc_hd__a2bb2o_4 _27473_ (.A1_N(_21156_),
    .A2_N(_21113_),
    .B1(_21129_),
    .B2(_21164_),
    .X(_00587_));
 sky130_vsdinv _27474_ (.A(mem_la_wdata[4]),
    .Y(_21165_));
 sky130_fd_sc_hd__buf_1 _27475_ (.A(_21165_),
    .X(_21166_));
 sky130_fd_sc_hd__buf_1 _27476_ (.A(_21166_),
    .X(_21167_));
 sky130_fd_sc_hd__buf_1 _27477_ (.A(_21167_),
    .X(_21168_));
 sky130_fd_sc_hd__buf_1 _27478_ (.A(_21168_),
    .X(_21169_));
 sky130_fd_sc_hd__buf_1 _27479_ (.A(_21111_),
    .X(_21170_));
 sky130_fd_sc_hd__buf_1 _27480_ (.A(_21170_),
    .X(_21171_));
 sky130_fd_sc_hd__buf_1 _27481_ (.A(\decoded_imm[4] ),
    .X(_21172_));
 sky130_vsdinv _27482_ (.A(_21172_),
    .Y(_21173_));
 sky130_fd_sc_hd__nor2_4 _27483_ (.A(\decoded_rs2[4] ),
    .B(_21157_),
    .Y(_21174_));
 sky130_fd_sc_hd__a211o_4 _27484_ (.A1(_21158_),
    .A2(_21173_),
    .B1(_21134_),
    .C1(_21174_),
    .X(_21175_));
 sky130_fd_sc_hd__o21ai_4 _27485_ (.A1(_21146_),
    .A2(_21035_),
    .B1(_21175_),
    .Y(_21176_));
 sky130_fd_sc_hd__a2bb2o_4 _27486_ (.A1_N(_21169_),
    .A2_N(_21171_),
    .B1(_21129_),
    .B2(_21176_),
    .X(_00588_));
 sky130_vsdinv _27487_ (.A(mem_la_wdata[5]),
    .Y(_21177_));
 sky130_fd_sc_hd__buf_1 _27488_ (.A(_21177_),
    .X(_21178_));
 sky130_fd_sc_hd__buf_1 _27489_ (.A(_21178_),
    .X(_21179_));
 sky130_fd_sc_hd__buf_1 _27490_ (.A(_21128_),
    .X(_21180_));
 sky130_fd_sc_hd__buf_1 _27491_ (.A(_18788_),
    .X(_21181_));
 sky130_fd_sc_hd__buf_1 _27492_ (.A(_21181_),
    .X(_21182_));
 sky130_fd_sc_hd__buf_1 _27493_ (.A(_21161_),
    .X(_21183_));
 sky130_fd_sc_hd__buf_1 _27494_ (.A(_19097_),
    .X(_21184_));
 sky130_fd_sc_hd__buf_1 _27495_ (.A(\decoded_imm[5] ),
    .X(_21185_));
 sky130_fd_sc_hd__buf_1 _27496_ (.A(_21185_),
    .X(_21186_));
 sky130_fd_sc_hd__nand3_4 _27497_ (.A(_21183_),
    .B(_21184_),
    .C(_21186_),
    .Y(_21187_));
 sky130_fd_sc_hd__o21ai_4 _27498_ (.A1(_21182_),
    .A2(_21038_),
    .B1(_21187_),
    .Y(_21188_));
 sky130_fd_sc_hd__a2bb2o_4 _27499_ (.A1_N(_21179_),
    .A2_N(_21171_),
    .B1(_21180_),
    .B2(_21188_),
    .X(_00589_));
 sky130_vsdinv _27500_ (.A(mem_la_wdata[6]),
    .Y(_21189_));
 sky130_fd_sc_hd__buf_1 _27501_ (.A(_21189_),
    .X(_21190_));
 sky130_fd_sc_hd__buf_1 _27502_ (.A(_20231_),
    .X(_21191_));
 sky130_fd_sc_hd__buf_1 _27503_ (.A(\decoded_imm[6] ),
    .X(_21192_));
 sky130_fd_sc_hd__buf_1 _27504_ (.A(_21192_),
    .X(_21193_));
 sky130_fd_sc_hd__nand3_4 _27505_ (.A(_21183_),
    .B(_21191_),
    .C(_21193_),
    .Y(_21194_));
 sky130_fd_sc_hd__o21ai_4 _27506_ (.A1(_21182_),
    .A2(_21044_),
    .B1(_21194_),
    .Y(_21195_));
 sky130_fd_sc_hd__a2bb2o_4 _27507_ (.A1_N(_21190_),
    .A2_N(_21171_),
    .B1(_21180_),
    .B2(_21195_),
    .X(_00590_));
 sky130_vsdinv _27508_ (.A(mem_la_wdata[7]),
    .Y(_21196_));
 sky130_fd_sc_hd__buf_1 _27509_ (.A(_21196_),
    .X(_21197_));
 sky130_fd_sc_hd__buf_1 _27510_ (.A(_21197_),
    .X(_21198_));
 sky130_fd_sc_hd__buf_1 _27511_ (.A(_21158_),
    .X(_21199_));
 sky130_fd_sc_hd__buf_1 _27512_ (.A(\decoded_imm[7] ),
    .X(_21200_));
 sky130_fd_sc_hd__buf_1 _27513_ (.A(_21200_),
    .X(_21201_));
 sky130_fd_sc_hd__nand3_4 _27514_ (.A(_21199_),
    .B(_21191_),
    .C(_21201_),
    .Y(_21202_));
 sky130_fd_sc_hd__o21ai_4 _27515_ (.A1(_21182_),
    .A2(_21047_),
    .B1(_21202_),
    .Y(_21203_));
 sky130_fd_sc_hd__a2bb2o_4 _27516_ (.A1_N(_21198_),
    .A2_N(_21171_),
    .B1(_21180_),
    .B2(_21203_),
    .X(_00591_));
 sky130_vsdinv _27517_ (.A(pcpi_rs2[8]),
    .Y(_21204_));
 sky130_fd_sc_hd__buf_1 _27518_ (.A(_21170_),
    .X(_21205_));
 sky130_fd_sc_hd__buf_1 _27519_ (.A(\decoded_imm[8] ),
    .X(_21206_));
 sky130_fd_sc_hd__buf_1 _27520_ (.A(_21206_),
    .X(_21207_));
 sky130_fd_sc_hd__nand3_4 _27521_ (.A(_21199_),
    .B(_21191_),
    .C(_21207_),
    .Y(_21208_));
 sky130_fd_sc_hd__o21ai_4 _27522_ (.A1(_21182_),
    .A2(_21049_),
    .B1(_21208_),
    .Y(_21209_));
 sky130_fd_sc_hd__a2bb2o_4 _27523_ (.A1_N(_21204_),
    .A2_N(_21205_),
    .B1(_21180_),
    .B2(_21209_),
    .X(_00592_));
 sky130_vsdinv _27524_ (.A(pcpi_rs2[9]),
    .Y(_21210_));
 sky130_fd_sc_hd__buf_1 _27525_ (.A(_21210_),
    .X(_21211_));
 sky130_fd_sc_hd__buf_1 _27526_ (.A(_19124_),
    .X(_21212_));
 sky130_fd_sc_hd__buf_1 _27527_ (.A(_21212_),
    .X(_21213_));
 sky130_fd_sc_hd__buf_1 _27528_ (.A(_18289_),
    .X(_21214_));
 sky130_fd_sc_hd__buf_1 _27529_ (.A(_21214_),
    .X(_21215_));
 sky130_fd_sc_hd__buf_1 _27530_ (.A(_21215_),
    .X(_21216_));
 sky130_fd_sc_hd__buf_1 _27531_ (.A(_21114_),
    .X(_21217_));
 sky130_vsdinv _27532_ (.A(\decoded_imm[9] ),
    .Y(_21218_));
 sky130_fd_sc_hd__buf_1 _27533_ (.A(_21130_),
    .X(_21219_));
 sky130_fd_sc_hd__o32ai_4 _27534_ (.A1(_21216_),
    .A2(_21217_),
    .A3(_21218_),
    .B1(_21219_),
    .B2(_21052_),
    .Y(_21220_));
 sky130_fd_sc_hd__a2bb2o_4 _27535_ (.A1_N(_21211_),
    .A2_N(_21205_),
    .B1(_21213_),
    .B2(_21220_),
    .X(_00593_));
 sky130_fd_sc_hd__buf_1 _27536_ (.A(\decoded_imm[10] ),
    .X(_21221_));
 sky130_fd_sc_hd__buf_1 _27537_ (.A(_21221_),
    .X(_21222_));
 sky130_fd_sc_hd__nand3_4 _27538_ (.A(_21183_),
    .B(_21184_),
    .C(_21222_),
    .Y(_21223_));
 sky130_fd_sc_hd__o21ai_4 _27539_ (.A1(_21146_),
    .A2(_19975_),
    .B1(_21223_),
    .Y(_21224_));
 sky130_fd_sc_hd__nor2_4 _27540_ (.A(\cpu_state[2] ),
    .B(_18533_),
    .Y(_21225_));
 sky130_fd_sc_hd__buf_1 _27541_ (.A(_21225_),
    .X(_21226_));
 sky130_fd_sc_hd__buf_1 _27542_ (.A(_18654_),
    .X(_21227_));
 sky130_fd_sc_hd__buf_1 _27543_ (.A(_21227_),
    .X(_21228_));
 sky130_fd_sc_hd__o21a_4 _27544_ (.A1(_18805_),
    .A2(_21226_),
    .B1(_21228_),
    .X(_21229_));
 sky130_fd_sc_hd__a21o_4 _27545_ (.A1(_21224_),
    .A2(_19112_),
    .B1(_21229_),
    .X(_00563_));
 sky130_vsdinv _27546_ (.A(pcpi_rs2[11]),
    .Y(_21230_));
 sky130_fd_sc_hd__buf_1 _27547_ (.A(_21181_),
    .X(_21231_));
 sky130_fd_sc_hd__buf_1 _27548_ (.A(\decoded_imm[11] ),
    .X(_21232_));
 sky130_fd_sc_hd__nand3_4 _27549_ (.A(_21199_),
    .B(_21191_),
    .C(_21232_),
    .Y(_21233_));
 sky130_fd_sc_hd__o21ai_4 _27550_ (.A1(_21231_),
    .A2(_20050_),
    .B1(_21233_),
    .Y(_21234_));
 sky130_fd_sc_hd__a2bb2o_4 _27551_ (.A1_N(_21230_),
    .A2_N(_21205_),
    .B1(_21213_),
    .B2(_21234_),
    .X(_00564_));
 sky130_vsdinv _27552_ (.A(pcpi_rs2[12]),
    .Y(_21235_));
 sky130_fd_sc_hd__buf_1 _27553_ (.A(_21235_),
    .X(_21236_));
 sky130_fd_sc_hd__buf_1 _27554_ (.A(_20231_),
    .X(_21237_));
 sky130_fd_sc_hd__buf_1 _27555_ (.A(\decoded_imm[12] ),
    .X(_21238_));
 sky130_fd_sc_hd__buf_1 _27556_ (.A(_21238_),
    .X(_21239_));
 sky130_fd_sc_hd__nand3_4 _27557_ (.A(_21199_),
    .B(_21237_),
    .C(_21239_),
    .Y(_21240_));
 sky130_fd_sc_hd__o21ai_4 _27558_ (.A1(_21231_),
    .A2(_20111_),
    .B1(_21240_),
    .Y(_21241_));
 sky130_fd_sc_hd__a2bb2o_4 _27559_ (.A1_N(_21236_),
    .A2_N(_21205_),
    .B1(_21213_),
    .B2(_21241_),
    .X(_00565_));
 sky130_vsdinv _27560_ (.A(pcpi_rs2[13]),
    .Y(_21242_));
 sky130_fd_sc_hd__buf_1 _27561_ (.A(_21242_),
    .X(_21243_));
 sky130_fd_sc_hd__buf_1 _27562_ (.A(_21243_),
    .X(_21244_));
 sky130_fd_sc_hd__buf_1 _27563_ (.A(_21170_),
    .X(_21245_));
 sky130_vsdinv _27564_ (.A(\decoded_imm[13] ),
    .Y(_21246_));
 sky130_fd_sc_hd__o32ai_4 _27565_ (.A1(_21216_),
    .A2(_21217_),
    .A3(_21246_),
    .B1(_21219_),
    .B2(_20170_),
    .Y(_21247_));
 sky130_fd_sc_hd__a2bb2o_4 _27566_ (.A1_N(_21244_),
    .A2_N(_21245_),
    .B1(_21213_),
    .B2(_21247_),
    .X(_00566_));
 sky130_vsdinv _27567_ (.A(pcpi_rs2[14]),
    .Y(_21248_));
 sky130_fd_sc_hd__buf_1 _27568_ (.A(_21248_),
    .X(_21249_));
 sky130_fd_sc_hd__buf_1 _27569_ (.A(_21249_),
    .X(_21250_));
 sky130_fd_sc_hd__buf_1 _27570_ (.A(_21212_),
    .X(_21251_));
 sky130_fd_sc_hd__buf_1 _27571_ (.A(_21161_),
    .X(_21252_));
 sky130_fd_sc_hd__buf_1 _27572_ (.A(\decoded_imm[14] ),
    .X(_21253_));
 sky130_fd_sc_hd__nand3_4 _27573_ (.A(_21252_),
    .B(_21237_),
    .C(_21253_),
    .Y(_21254_));
 sky130_fd_sc_hd__o21ai_4 _27574_ (.A1(_21231_),
    .A2(_20226_),
    .B1(_21254_),
    .Y(_21255_));
 sky130_fd_sc_hd__a2bb2o_4 _27575_ (.A1_N(_21250_),
    .A2_N(_21245_),
    .B1(_21251_),
    .B2(_21255_),
    .X(_00567_));
 sky130_vsdinv _27576_ (.A(pcpi_rs2[15]),
    .Y(_21256_));
 sky130_fd_sc_hd__buf_1 _27577_ (.A(_21256_),
    .X(_21257_));
 sky130_fd_sc_hd__buf_1 _27578_ (.A(\decoded_imm[15] ),
    .X(_21258_));
 sky130_vsdinv _27579_ (.A(_21258_),
    .Y(_21259_));
 sky130_fd_sc_hd__buf_1 _27580_ (.A(_21181_),
    .X(_21260_));
 sky130_fd_sc_hd__o32ai_4 _27581_ (.A1(_21216_),
    .A2(_21217_),
    .A3(_21259_),
    .B1(_21260_),
    .B2(_20275_),
    .Y(_21261_));
 sky130_fd_sc_hd__a2bb2o_4 _27582_ (.A1_N(_21257_),
    .A2_N(_21245_),
    .B1(_21251_),
    .B2(_21261_),
    .X(_00568_));
 sky130_vsdinv _27583_ (.A(_18711_),
    .Y(_21262_));
 sky130_fd_sc_hd__buf_1 _27584_ (.A(\decoded_imm[16] ),
    .X(_21263_));
 sky130_fd_sc_hd__buf_1 _27585_ (.A(_21263_),
    .X(_21264_));
 sky130_fd_sc_hd__nand3_4 _27586_ (.A(_21252_),
    .B(_21237_),
    .C(_21264_),
    .Y(_21265_));
 sky130_fd_sc_hd__o21ai_4 _27587_ (.A1(_21231_),
    .A2(_21076_),
    .B1(_21265_),
    .Y(_21266_));
 sky130_fd_sc_hd__a2bb2o_4 _27588_ (.A1_N(_21262_),
    .A2_N(_21245_),
    .B1(_21251_),
    .B2(_21266_),
    .X(_00569_));
 sky130_vsdinv _27589_ (.A(pcpi_rs2[17]),
    .Y(_21267_));
 sky130_fd_sc_hd__buf_1 _27590_ (.A(_21170_),
    .X(_21268_));
 sky130_fd_sc_hd__buf_1 _27591_ (.A(_21181_),
    .X(_21269_));
 sky130_fd_sc_hd__buf_1 _27592_ (.A(\decoded_imm[17] ),
    .X(_21270_));
 sky130_fd_sc_hd__nand3_4 _27593_ (.A(_21252_),
    .B(_21237_),
    .C(_21270_),
    .Y(_21271_));
 sky130_fd_sc_hd__o21ai_4 _27594_ (.A1(_21269_),
    .A2(_20374_),
    .B1(_21271_),
    .Y(_21272_));
 sky130_fd_sc_hd__a2bb2o_4 _27595_ (.A1_N(_21267_),
    .A2_N(_21268_),
    .B1(_21251_),
    .B2(_21272_),
    .X(_00570_));
 sky130_fd_sc_hd__buf_1 _27596_ (.A(_21212_),
    .X(_21273_));
 sky130_fd_sc_hd__buf_1 _27597_ (.A(\decoded_imm[18] ),
    .X(_21274_));
 sky130_vsdinv _27598_ (.A(_21274_),
    .Y(_21275_));
 sky130_fd_sc_hd__o32ai_4 _27599_ (.A1(_21216_),
    .A2(_21217_),
    .A3(_21275_),
    .B1(_21260_),
    .B2(_20428_),
    .Y(_21276_));
 sky130_fd_sc_hd__a2bb2o_4 _27600_ (.A1_N(_18703_),
    .A2_N(_21268_),
    .B1(_21273_),
    .B2(_21276_),
    .X(_00571_));
 sky130_vsdinv _27601_ (.A(pcpi_rs2[19]),
    .Y(_21277_));
 sky130_fd_sc_hd__buf_1 _27602_ (.A(_18290_),
    .X(_21278_));
 sky130_fd_sc_hd__buf_1 _27603_ (.A(_21278_),
    .X(_21279_));
 sky130_fd_sc_hd__buf_1 _27604_ (.A(_21114_),
    .X(_21280_));
 sky130_fd_sc_hd__buf_1 _27605_ (.A(\decoded_imm[19] ),
    .X(_21281_));
 sky130_vsdinv _27606_ (.A(_21281_),
    .Y(_21282_));
 sky130_fd_sc_hd__o32ai_4 _27607_ (.A1(_21279_),
    .A2(_21280_),
    .A3(_21282_),
    .B1(_21260_),
    .B2(_20478_),
    .Y(_21283_));
 sky130_fd_sc_hd__a2bb2o_4 _27608_ (.A1_N(_21277_),
    .A2_N(_21268_),
    .B1(_21273_),
    .B2(_21283_),
    .X(_00572_));
 sky130_vsdinv _27609_ (.A(_18668_),
    .Y(_21284_));
 sky130_fd_sc_hd__buf_1 _27610_ (.A(_20231_),
    .X(_21285_));
 sky130_fd_sc_hd__buf_1 _27611_ (.A(\decoded_imm[20] ),
    .X(_21286_));
 sky130_fd_sc_hd__nand3_4 _27612_ (.A(_21252_),
    .B(_21285_),
    .C(_21286_),
    .Y(_21287_));
 sky130_fd_sc_hd__o21ai_4 _27613_ (.A1(_21269_),
    .A2(_21084_),
    .B1(_21287_),
    .Y(_21288_));
 sky130_fd_sc_hd__a2bb2o_4 _27614_ (.A1_N(_21284_),
    .A2_N(_21268_),
    .B1(_21273_),
    .B2(_21288_),
    .X(_00574_));
 sky130_vsdinv _27615_ (.A(pcpi_rs2[21]),
    .Y(_21289_));
 sky130_fd_sc_hd__buf_1 _27616_ (.A(_21111_),
    .X(_21290_));
 sky130_fd_sc_hd__buf_1 _27617_ (.A(_21161_),
    .X(_21291_));
 sky130_fd_sc_hd__buf_1 _27618_ (.A(\decoded_imm[21] ),
    .X(_21292_));
 sky130_fd_sc_hd__nand3_4 _27619_ (.A(_21291_),
    .B(_21285_),
    .C(_21292_),
    .Y(_21293_));
 sky130_fd_sc_hd__o21ai_4 _27620_ (.A1(_21269_),
    .A2(_20573_),
    .B1(_21293_),
    .Y(_21294_));
 sky130_fd_sc_hd__a2bb2o_4 _27621_ (.A1_N(_21289_),
    .A2_N(_21290_),
    .B1(_21273_),
    .B2(_21294_),
    .X(_00575_));
 sky130_fd_sc_hd__buf_1 _27622_ (.A(_21212_),
    .X(_21295_));
 sky130_fd_sc_hd__buf_1 _27623_ (.A(\decoded_imm[22] ),
    .X(_21296_));
 sky130_vsdinv _27624_ (.A(_21296_),
    .Y(_21297_));
 sky130_fd_sc_hd__o32ai_4 _27625_ (.A1(_21279_),
    .A2(_21280_),
    .A3(_21297_),
    .B1(_21260_),
    .B2(_20617_),
    .Y(_21298_));
 sky130_fd_sc_hd__a2bb2o_4 _27626_ (.A1_N(_18674_),
    .A2_N(_21290_),
    .B1(_21295_),
    .B2(_21298_),
    .X(_00576_));
 sky130_vsdinv _27627_ (.A(pcpi_rs2[23]),
    .Y(_21299_));
 sky130_fd_sc_hd__buf_1 _27628_ (.A(_21299_),
    .X(_21300_));
 sky130_vsdinv _27629_ (.A(\decoded_imm[23] ),
    .Y(_21301_));
 sky130_fd_sc_hd__buf_1 _27630_ (.A(_21130_),
    .X(_21302_));
 sky130_fd_sc_hd__o32ai_4 _27631_ (.A1(_21279_),
    .A2(_21280_),
    .A3(_21301_),
    .B1(_21302_),
    .B2(_20657_),
    .Y(_21303_));
 sky130_fd_sc_hd__a2bb2o_4 _27632_ (.A1_N(_21300_),
    .A2_N(_21290_),
    .B1(_21295_),
    .B2(_21303_),
    .X(_00577_));
 sky130_fd_sc_hd__a2111o_4 _27633_ (.A1(_20680_),
    .A2(_20695_),
    .B1(_21130_),
    .C1(_21028_),
    .D1(_20703_),
    .X(_21304_));
 sky130_fd_sc_hd__buf_1 _27634_ (.A(\decoded_imm[24] ),
    .X(_21305_));
 sky130_fd_sc_hd__nand3_4 _27635_ (.A(_21158_),
    .B(_20232_),
    .C(_21305_),
    .Y(_21306_));
 sky130_fd_sc_hd__nand2_4 _27636_ (.A(_21304_),
    .B(_21306_),
    .Y(_21307_));
 sky130_fd_sc_hd__a2bb2o_4 _27637_ (.A1_N(_18729_),
    .A2_N(_21290_),
    .B1(_21295_),
    .B2(_21307_),
    .X(_00578_));
 sky130_vsdinv _27638_ (.A(pcpi_rs2[25]),
    .Y(_21308_));
 sky130_fd_sc_hd__buf_1 _27639_ (.A(_21308_),
    .X(_21309_));
 sky130_fd_sc_hd__buf_1 _27640_ (.A(_21111_),
    .X(_21310_));
 sky130_fd_sc_hd__buf_1 _27641_ (.A(\decoded_imm[25] ),
    .X(_21311_));
 sky130_vsdinv _27642_ (.A(_21311_),
    .Y(_21312_));
 sky130_fd_sc_hd__o32ai_4 _27643_ (.A1(_21279_),
    .A2(_21280_),
    .A3(_21312_),
    .B1(_21302_),
    .B2(_21094_),
    .Y(_21313_));
 sky130_fd_sc_hd__a2bb2o_4 _27644_ (.A1_N(_21309_),
    .A2_N(_21310_),
    .B1(_21295_),
    .B2(_21313_),
    .X(_00579_));
 sky130_vsdinv _27645_ (.A(pcpi_rs2[26]),
    .Y(_21314_));
 sky130_fd_sc_hd__buf_1 _27646_ (.A(_21314_),
    .X(_21315_));
 sky130_fd_sc_hd__buf_1 _27647_ (.A(_18861_),
    .X(_21316_));
 sky130_fd_sc_hd__buf_1 _27648_ (.A(_21278_),
    .X(_21317_));
 sky130_fd_sc_hd__buf_1 _27649_ (.A(\decoded_imm[26] ),
    .X(_21318_));
 sky130_vsdinv _27650_ (.A(_21318_),
    .Y(_21319_));
 sky130_fd_sc_hd__o32ai_4 _27651_ (.A1(_21317_),
    .A2(_21132_),
    .A3(_21319_),
    .B1(_21302_),
    .B2(_21097_),
    .Y(_21320_));
 sky130_fd_sc_hd__a2bb2o_4 _27652_ (.A1_N(_21315_),
    .A2_N(_21310_),
    .B1(_21316_),
    .B2(_21320_),
    .X(_00580_));
 sky130_fd_sc_hd__buf_1 _27653_ (.A(\decoded_imm[27] ),
    .X(_21321_));
 sky130_vsdinv _27654_ (.A(_21321_),
    .Y(_21322_));
 sky130_fd_sc_hd__o32ai_4 _27655_ (.A1(_21317_),
    .A2(_21132_),
    .A3(_21322_),
    .B1(_21302_),
    .B2(_20842_),
    .Y(_21323_));
 sky130_fd_sc_hd__a2bb2o_4 _27656_ (.A1_N(_18760_),
    .A2_N(_21310_),
    .B1(_21316_),
    .B2(_21323_),
    .X(_00581_));
 sky130_vsdinv _27657_ (.A(pcpi_rs2[28]),
    .Y(_21324_));
 sky130_fd_sc_hd__buf_1 _27658_ (.A(_21324_),
    .X(_21325_));
 sky130_fd_sc_hd__buf_1 _27659_ (.A(\decoded_imm[28] ),
    .X(_21326_));
 sky130_fd_sc_hd__nand3_4 _27660_ (.A(_21291_),
    .B(_21285_),
    .C(_21326_),
    .Y(_21327_));
 sky130_fd_sc_hd__o21ai_4 _27661_ (.A1(_21269_),
    .A2(_21101_),
    .B1(_21327_),
    .Y(_21328_));
 sky130_fd_sc_hd__a2bb2o_4 _27662_ (.A1_N(_21325_),
    .A2_N(_21310_),
    .B1(_21316_),
    .B2(_21328_),
    .X(_00582_));
 sky130_vsdinv _27663_ (.A(pcpi_rs2[29]),
    .Y(_21329_));
 sky130_fd_sc_hd__buf_1 _27664_ (.A(\decoded_imm[29] ),
    .X(_21330_));
 sky130_fd_sc_hd__buf_1 _27665_ (.A(_21330_),
    .X(_21331_));
 sky130_fd_sc_hd__nand3_4 _27666_ (.A(_21291_),
    .B(_21285_),
    .C(_21331_),
    .Y(_21332_));
 sky130_fd_sc_hd__o21ai_4 _27667_ (.A1(_21219_),
    .A2(_20930_),
    .B1(_21332_),
    .Y(_21333_));
 sky130_fd_sc_hd__a2bb2o_4 _27668_ (.A1_N(_21329_),
    .A2_N(_21112_),
    .B1(_21316_),
    .B2(_21333_),
    .X(_00583_));
 sky130_vsdinv _27669_ (.A(pcpi_rs2[30]),
    .Y(_21334_));
 sky130_fd_sc_hd__buf_1 _27670_ (.A(_21128_),
    .X(_21335_));
 sky130_fd_sc_hd__buf_1 _27671_ (.A(\decoded_imm[30] ),
    .X(_21336_));
 sky130_fd_sc_hd__nand3_4 _27672_ (.A(_21291_),
    .B(_20232_),
    .C(_21336_),
    .Y(_21337_));
 sky130_fd_sc_hd__o21ai_4 _27673_ (.A1(_21219_),
    .A2(_21104_),
    .B1(_21337_),
    .Y(_21338_));
 sky130_fd_sc_hd__a2bb2o_4 _27674_ (.A1_N(_21334_),
    .A2_N(_21112_),
    .B1(_21335_),
    .B2(_21338_),
    .X(_00585_));
 sky130_fd_sc_hd__buf_1 _27675_ (.A(pcpi_rs2[31]),
    .X(_21339_));
 sky130_vsdinv _27676_ (.A(_21339_),
    .Y(_21340_));
 sky130_vsdinv _27677_ (.A(\decoded_imm[31] ),
    .Y(_21341_));
 sky130_fd_sc_hd__o32ai_4 _27678_ (.A1(_21317_),
    .A2(_21132_),
    .A3(_21341_),
    .B1(_18806_),
    .B2(_21106_),
    .Y(_21342_));
 sky130_fd_sc_hd__a2bb2o_4 _27679_ (.A1_N(_21340_),
    .A2_N(_21112_),
    .B1(_21335_),
    .B2(_21342_),
    .X(_00586_));
 sky130_vsdinv _27680_ (.A(_18296_),
    .Y(_21343_));
 sky130_fd_sc_hd__buf_1 _27681_ (.A(_21343_),
    .X(_21344_));
 sky130_fd_sc_hd__buf_1 _27682_ (.A(_21118_),
    .X(_21345_));
 sky130_fd_sc_hd__a21oi_4 _27683_ (.A1(_18272_),
    .A2(_18288_),
    .B1(_18224_),
    .Y(_21346_));
 sky130_vsdinv _27684_ (.A(_21346_),
    .Y(_21347_));
 sky130_fd_sc_hd__nor2_4 _27685_ (.A(_18281_),
    .B(_21347_),
    .Y(_21348_));
 sky130_fd_sc_hd__o21ai_4 _27686_ (.A1(_21345_),
    .A2(_18273_),
    .B1(_21348_),
    .Y(_21349_));
 sky130_fd_sc_hd__a21oi_4 _27687_ (.A1(_18259_),
    .A2(_18518_),
    .B1(_21349_),
    .Y(_21350_));
 sky130_fd_sc_hd__buf_1 _27688_ (.A(_18300_),
    .X(_21351_));
 sky130_vsdinv _27689_ (.A(_21345_),
    .Y(_21352_));
 sky130_fd_sc_hd__a22oi_4 _27690_ (.A1(_18245_),
    .A2(\cpu_state[5] ),
    .B1(_18236_),
    .B2(_18238_),
    .Y(_21353_));
 sky130_fd_sc_hd__nor4_4 _27691_ (.A(_21351_),
    .B(_21352_),
    .C(_21353_),
    .D(_18848_),
    .Y(_21354_));
 sky130_fd_sc_hd__buf_1 _27692_ (.A(_18795_),
    .X(_21355_));
 sky130_fd_sc_hd__buf_1 _27693_ (.A(_19193_),
    .X(_21356_));
 sky130_fd_sc_hd__or4_4 _27694_ (.A(_21355_),
    .B(_21356_),
    .C(_19226_),
    .D(_19281_),
    .X(_21357_));
 sky130_vsdinv _27695_ (.A(instr_lui),
    .Y(_21358_));
 sky130_fd_sc_hd__buf_1 _27696_ (.A(_21358_),
    .X(_21359_));
 sky130_fd_sc_hd__buf_1 _27697_ (.A(_21359_),
    .X(_21360_));
 sky130_fd_sc_hd__buf_1 _27698_ (.A(\reg_pc[0] ),
    .X(_21361_));
 sky130_fd_sc_hd__buf_1 _27699_ (.A(_21355_),
    .X(_21362_));
 sky130_fd_sc_hd__nand3_4 _27700_ (.A(_21360_),
    .B(_21361_),
    .C(_21362_),
    .Y(_21363_));
 sky130_fd_sc_hd__a21oi_4 _27701_ (.A1(_21357_),
    .A2(_21363_),
    .B1(_21317_),
    .Y(_21364_));
 sky130_fd_sc_hd__o21ai_4 _27702_ (.A1(_21354_),
    .A2(_21364_),
    .B1(_18862_),
    .Y(_21365_));
 sky130_fd_sc_hd__o21ai_4 _27703_ (.A1(_21344_),
    .A2(_21350_),
    .B1(_21365_),
    .Y(_00530_));
 sky130_vsdinv _27704_ (.A(pcpi_rs1[1]),
    .Y(_21366_));
 sky130_fd_sc_hd__buf_1 _27705_ (.A(_21366_),
    .X(_21367_));
 sky130_fd_sc_hd__buf_1 _27706_ (.A(_21367_),
    .X(_21368_));
 sky130_fd_sc_hd__buf_1 _27707_ (.A(_21368_),
    .X(_21369_));
 sky130_vsdinv _27708_ (.A(_18257_),
    .Y(_21370_));
 sky130_fd_sc_hd__buf_1 _27709_ (.A(_21370_),
    .X(_21371_));
 sky130_fd_sc_hd__nand2_4 _27710_ (.A(_18296_),
    .B(_21118_),
    .Y(_21372_));
 sky130_vsdinv _27711_ (.A(_21135_),
    .Y(_21373_));
 sky130_fd_sc_hd__nand2_4 _27712_ (.A(_21372_),
    .B(_21373_),
    .Y(_21374_));
 sky130_fd_sc_hd__nand3_4 _27713_ (.A(_18296_),
    .B(_21118_),
    .C(_21135_),
    .Y(_21375_));
 sky130_fd_sc_hd__and3_4 _27714_ (.A(_21371_),
    .B(_21374_),
    .C(_21375_),
    .X(_21376_));
 sky130_fd_sc_hd__o21a_4 _27715_ (.A1(_18273_),
    .A2(_21376_),
    .B1(_21348_),
    .X(_21377_));
 sky130_fd_sc_hd__buf_1 _27716_ (.A(_18620_),
    .X(_21378_));
 sky130_fd_sc_hd__buf_1 _27717_ (.A(_21378_),
    .X(_21379_));
 sky130_fd_sc_hd__buf_1 _27718_ (.A(_21379_),
    .X(_21380_));
 sky130_fd_sc_hd__nor2_4 _27719_ (.A(_21380_),
    .B(_21353_),
    .Y(_21381_));
 sky130_fd_sc_hd__and4_4 _27720_ (.A(_21371_),
    .B(_21374_),
    .C(_21375_),
    .D(_21381_),
    .X(_21382_));
 sky130_fd_sc_hd__buf_1 _27721_ (.A(_18795_),
    .X(_21383_));
 sky130_fd_sc_hd__a2111o_4 _27722_ (.A1(_19331_),
    .A2(_19378_),
    .B1(_21383_),
    .C1(_19194_),
    .D1(_19411_),
    .X(_21384_));
 sky130_fd_sc_hd__nand3_4 _27723_ (.A(_21360_),
    .B(_18304_),
    .C(_21362_),
    .Y(_21385_));
 sky130_fd_sc_hd__buf_1 _27724_ (.A(_21278_),
    .X(_21386_));
 sky130_fd_sc_hd__a21oi_4 _27725_ (.A1(_21384_),
    .A2(_21385_),
    .B1(_21386_),
    .Y(_21387_));
 sky130_fd_sc_hd__o21ai_4 _27726_ (.A1(_21382_),
    .A2(_21387_),
    .B1(_18862_),
    .Y(_21388_));
 sky130_fd_sc_hd__o21ai_4 _27727_ (.A1(_21369_),
    .A2(_21377_),
    .B1(_21388_),
    .Y(_00541_));
 sky130_vsdinv _27728_ (.A(_18613_),
    .Y(_21389_));
 sky130_fd_sc_hd__nand2_4 _27729_ (.A(_21370_),
    .B(_18245_),
    .Y(_21390_));
 sky130_fd_sc_hd__buf_1 _27730_ (.A(_18235_),
    .X(_21391_));
 sky130_fd_sc_hd__o21a_4 _27731_ (.A1(_21391_),
    .A2(_18257_),
    .B1(_18238_),
    .X(_21392_));
 sky130_fd_sc_hd__a211o_4 _27732_ (.A1(_21390_),
    .A2(_18242_),
    .B1(_21347_),
    .C1(_21392_),
    .X(_21393_));
 sky130_vsdinv _27733_ (.A(_21393_),
    .Y(_21394_));
 sky130_fd_sc_hd__buf_1 _27734_ (.A(_21394_),
    .X(_21395_));
 sky130_fd_sc_hd__buf_1 _27735_ (.A(_21395_),
    .X(_21396_));
 sky130_fd_sc_hd__buf_1 _27736_ (.A(_18613_),
    .X(_21397_));
 sky130_fd_sc_hd__xnor2_4 _27737_ (.A(_21397_),
    .B(_21147_),
    .Y(_21398_));
 sky130_fd_sc_hd__nand2_4 _27738_ (.A(_21375_),
    .B(_21366_),
    .Y(_21399_));
 sky130_fd_sc_hd__and2_4 _27739_ (.A(_21399_),
    .B(_21374_),
    .X(_21400_));
 sky130_fd_sc_hd__xor2_4 _27740_ (.A(_21398_),
    .B(_21400_),
    .X(_21401_));
 sky130_fd_sc_hd__nor3_4 _27741_ (.A(_21353_),
    .B(_21401_),
    .C(_18848_),
    .Y(_21402_));
 sky130_fd_sc_hd__a2111o_4 _27742_ (.A1(_19450_),
    .A2(_19478_),
    .B1(_21383_),
    .C1(_19194_),
    .D1(_19489_),
    .X(_21403_));
 sky130_fd_sc_hd__buf_1 _27743_ (.A(\reg_pc[2] ),
    .X(_21404_));
 sky130_fd_sc_hd__nand3_4 _27744_ (.A(_21360_),
    .B(_21362_),
    .C(_21404_),
    .Y(_21405_));
 sky130_fd_sc_hd__a21oi_4 _27745_ (.A1(_21403_),
    .A2(_21405_),
    .B1(_21386_),
    .Y(_21406_));
 sky130_fd_sc_hd__o21ai_4 _27746_ (.A1(_21402_),
    .A2(_21406_),
    .B1(_20932_),
    .Y(_21407_));
 sky130_fd_sc_hd__o21ai_4 _27747_ (.A1(_21389_),
    .A2(_21396_),
    .B1(_21407_),
    .Y(_00552_));
 sky130_fd_sc_hd__buf_1 _27748_ (.A(_18607_),
    .X(_21408_));
 sky130_vsdinv _27749_ (.A(_21408_),
    .Y(_21409_));
 sky130_fd_sc_hd__buf_1 _27750_ (.A(_18794_),
    .X(_21410_));
 sky130_fd_sc_hd__buf_1 _27751_ (.A(_20102_),
    .X(_21411_));
 sky130_fd_sc_hd__a2111o_4 _27752_ (.A1(_19523_),
    .A2(_19551_),
    .B1(_21410_),
    .C1(_21411_),
    .D1(_19562_),
    .X(_21412_));
 sky130_fd_sc_hd__buf_1 _27753_ (.A(_21358_),
    .X(_21413_));
 sky130_fd_sc_hd__buf_1 _27754_ (.A(_21413_),
    .X(_21414_));
 sky130_fd_sc_hd__buf_1 _27755_ (.A(_18794_),
    .X(_21415_));
 sky130_fd_sc_hd__buf_1 _27756_ (.A(_21415_),
    .X(_21416_));
 sky130_fd_sc_hd__buf_1 _27757_ (.A(\reg_pc[3] ),
    .X(_21417_));
 sky130_fd_sc_hd__buf_1 _27758_ (.A(_21417_),
    .X(_21418_));
 sky130_fd_sc_hd__nand3_4 _27759_ (.A(_21414_),
    .B(_21416_),
    .C(_21418_),
    .Y(_21419_));
 sky130_fd_sc_hd__a21o_4 _27760_ (.A1(_21412_),
    .A2(_21419_),
    .B1(_18292_),
    .X(_21420_));
 sky130_fd_sc_hd__buf_1 _27761_ (.A(_21408_),
    .X(_21421_));
 sky130_fd_sc_hd__xor2_4 _27762_ (.A(_21421_),
    .B(_21159_),
    .X(_21422_));
 sky130_fd_sc_hd__nor2_4 _27763_ (.A(_18612_),
    .B(_21147_),
    .Y(_21423_));
 sky130_fd_sc_hd__a22oi_4 _27764_ (.A1(_18612_),
    .A2(\decoded_imm[2] ),
    .B1(_21399_),
    .B2(_21374_),
    .Y(_21424_));
 sky130_fd_sc_hd__nor2_4 _27765_ (.A(_21423_),
    .B(_21424_),
    .Y(_21425_));
 sky130_fd_sc_hd__nor2_4 _27766_ (.A(_21353_),
    .B(_18258_),
    .Y(_21426_));
 sky130_fd_sc_hd__buf_1 _27767_ (.A(_21426_),
    .X(_21427_));
 sky130_fd_sc_hd__buf_1 _27768_ (.A(_21427_),
    .X(_21428_));
 sky130_fd_sc_hd__o21ai_4 _27769_ (.A1(_21422_),
    .A2(_21425_),
    .B1(_21428_),
    .Y(_21429_));
 sky130_fd_sc_hd__a21o_4 _27770_ (.A1(_21422_),
    .A2(_21425_),
    .B1(_21429_),
    .X(_21430_));
 sky130_fd_sc_hd__buf_1 _27771_ (.A(_18477_),
    .X(_21431_));
 sky130_fd_sc_hd__buf_1 _27772_ (.A(_21431_),
    .X(_21432_));
 sky130_fd_sc_hd__a21o_4 _27773_ (.A1(_21420_),
    .A2(_21430_),
    .B1(_21432_),
    .X(_21433_));
 sky130_fd_sc_hd__o21ai_4 _27774_ (.A1(_21409_),
    .A2(_21396_),
    .B1(_21433_),
    .Y(_00555_));
 sky130_fd_sc_hd__buf_1 _27775_ (.A(_18600_),
    .X(_21434_));
 sky130_vsdinv _27776_ (.A(_21434_),
    .Y(_21435_));
 sky130_fd_sc_hd__buf_1 _27777_ (.A(is_lui_auipc_jal),
    .X(_21436_));
 sky130_fd_sc_hd__buf_1 _27778_ (.A(_21436_),
    .X(_21437_));
 sky130_fd_sc_hd__a2111o_4 _27779_ (.A1(_19604_),
    .A2(_19629_),
    .B1(_21437_),
    .C1(_21411_),
    .D1(_19648_),
    .X(_21438_));
 sky130_fd_sc_hd__buf_1 _27780_ (.A(_18794_),
    .X(_21439_));
 sky130_fd_sc_hd__buf_1 _27781_ (.A(_21439_),
    .X(_21440_));
 sky130_fd_sc_hd__buf_1 _27782_ (.A(\reg_pc[4] ),
    .X(_21441_));
 sky130_fd_sc_hd__nand3_4 _27783_ (.A(_21414_),
    .B(_21440_),
    .C(_21441_),
    .Y(_21442_));
 sky130_fd_sc_hd__a21o_4 _27784_ (.A1(_21438_),
    .A2(_21442_),
    .B1(_18292_),
    .X(_21443_));
 sky130_fd_sc_hd__xnor2_4 _27785_ (.A(_21434_),
    .B(_21172_),
    .Y(_21444_));
 sky130_fd_sc_hd__nand2_4 _27786_ (.A(pcpi_rs1[3]),
    .B(_21159_),
    .Y(_21445_));
 sky130_fd_sc_hd__o21ai_4 _27787_ (.A1(_21423_),
    .A2(_21424_),
    .B1(_21445_),
    .Y(_21446_));
 sky130_fd_sc_hd__nor2_4 _27788_ (.A(pcpi_rs1[3]),
    .B(\decoded_imm[3] ),
    .Y(_21447_));
 sky130_vsdinv _27789_ (.A(_21447_),
    .Y(_21448_));
 sky130_fd_sc_hd__and2_4 _27790_ (.A(_21446_),
    .B(_21448_),
    .X(_21449_));
 sky130_vsdinv _27791_ (.A(_21449_),
    .Y(_21450_));
 sky130_fd_sc_hd__buf_1 _27792_ (.A(_21426_),
    .X(_21451_));
 sky130_fd_sc_hd__a21boi_4 _27793_ (.A1(_21444_),
    .A2(_21450_),
    .B1_N(_21451_),
    .Y(_21452_));
 sky130_fd_sc_hd__o21ai_4 _27794_ (.A1(_21444_),
    .A2(_21450_),
    .B1(_21452_),
    .Y(_21453_));
 sky130_fd_sc_hd__a21o_4 _27795_ (.A1(_21443_),
    .A2(_21453_),
    .B1(_21432_),
    .X(_21454_));
 sky130_fd_sc_hd__o21ai_4 _27796_ (.A1(_21435_),
    .A2(_21396_),
    .B1(_21454_),
    .Y(_00556_));
 sky130_vsdinv _27797_ (.A(_18581_),
    .Y(_21455_));
 sky130_fd_sc_hd__a2111o_4 _27798_ (.A1(_19671_),
    .A2(_19686_),
    .B1(_21437_),
    .C1(_21411_),
    .D1(_19693_),
    .X(_21456_));
 sky130_fd_sc_hd__buf_1 _27799_ (.A(\reg_pc[5] ),
    .X(_21457_));
 sky130_fd_sc_hd__buf_1 _27800_ (.A(_21457_),
    .X(_21458_));
 sky130_fd_sc_hd__nand3_4 _27801_ (.A(_21414_),
    .B(_21440_),
    .C(_21458_),
    .Y(_21459_));
 sky130_fd_sc_hd__buf_1 _27802_ (.A(_18291_),
    .X(_21460_));
 sky130_fd_sc_hd__a21o_4 _27803_ (.A1(_21456_),
    .A2(_21459_),
    .B1(_21460_),
    .X(_21461_));
 sky130_fd_sc_hd__buf_1 _27804_ (.A(_18582_),
    .X(_21462_));
 sky130_fd_sc_hd__xor2_4 _27805_ (.A(_21462_),
    .B(_21186_),
    .X(_21463_));
 sky130_fd_sc_hd__nor2_4 _27806_ (.A(_18599_),
    .B(_21172_),
    .Y(_21464_));
 sky130_fd_sc_hd__a22oi_4 _27807_ (.A1(_18599_),
    .A2(_21172_),
    .B1(_21446_),
    .B2(_21448_),
    .Y(_21465_));
 sky130_fd_sc_hd__nor2_4 _27808_ (.A(_21464_),
    .B(_21465_),
    .Y(_21466_));
 sky130_fd_sc_hd__o21ai_4 _27809_ (.A1(_21463_),
    .A2(_21466_),
    .B1(_21428_),
    .Y(_21467_));
 sky130_fd_sc_hd__a21o_4 _27810_ (.A1(_21463_),
    .A2(_21466_),
    .B1(_21467_),
    .X(_21468_));
 sky130_fd_sc_hd__a21o_4 _27811_ (.A1(_21461_),
    .A2(_21468_),
    .B1(_21432_),
    .X(_21469_));
 sky130_fd_sc_hd__o21ai_4 _27812_ (.A1(_21455_),
    .A2(_21396_),
    .B1(_21469_),
    .Y(_00557_));
 sky130_vsdinv _27813_ (.A(pcpi_rs1[6]),
    .Y(_21470_));
 sky130_fd_sc_hd__buf_1 _27814_ (.A(_21470_),
    .X(_21471_));
 sky130_fd_sc_hd__buf_1 _27815_ (.A(_21395_),
    .X(_21472_));
 sky130_fd_sc_hd__a2111o_4 _27816_ (.A1(_19719_),
    .A2(_19738_),
    .B1(_21437_),
    .C1(_20103_),
    .D1(_19749_),
    .X(_21473_));
 sky130_fd_sc_hd__buf_1 _27817_ (.A(\reg_pc[6] ),
    .X(_21474_));
 sky130_fd_sc_hd__buf_1 _27818_ (.A(_21474_),
    .X(_21475_));
 sky130_fd_sc_hd__buf_1 _27819_ (.A(_21475_),
    .X(_21476_));
 sky130_fd_sc_hd__nand3_4 _27820_ (.A(_21414_),
    .B(_21440_),
    .C(_21476_),
    .Y(_21477_));
 sky130_fd_sc_hd__a21o_4 _27821_ (.A1(_21473_),
    .A2(_21477_),
    .B1(_21460_),
    .X(_21478_));
 sky130_fd_sc_hd__buf_1 _27822_ (.A(_18594_),
    .X(_21479_));
 sky130_fd_sc_hd__xnor2_4 _27823_ (.A(_21479_),
    .B(_21192_),
    .Y(_21480_));
 sky130_fd_sc_hd__maj3_4 _27824_ (.A(_21462_),
    .B(_21466_),
    .C(_21185_),
    .X(_21481_));
 sky130_vsdinv _27825_ (.A(_21481_),
    .Y(_21482_));
 sky130_fd_sc_hd__a21boi_4 _27826_ (.A1(_21482_),
    .A2(_21480_),
    .B1_N(_21427_),
    .Y(_21483_));
 sky130_fd_sc_hd__o21ai_4 _27827_ (.A1(_21480_),
    .A2(_21482_),
    .B1(_21483_),
    .Y(_21484_));
 sky130_fd_sc_hd__a21o_4 _27828_ (.A1(_21478_),
    .A2(_21484_),
    .B1(_21432_),
    .X(_21485_));
 sky130_fd_sc_hd__o21ai_4 _27829_ (.A1(_21471_),
    .A2(_21472_),
    .B1(_21485_),
    .Y(_00558_));
 sky130_vsdinv _27830_ (.A(pcpi_rs1[7]),
    .Y(_21486_));
 sky130_fd_sc_hd__a2111o_4 _27831_ (.A1(_19770_),
    .A2(_19785_),
    .B1(_21437_),
    .C1(_20103_),
    .D1(_19797_),
    .X(_21487_));
 sky130_fd_sc_hd__buf_1 _27832_ (.A(_21413_),
    .X(_21488_));
 sky130_fd_sc_hd__buf_1 _27833_ (.A(\reg_pc[7] ),
    .X(_21489_));
 sky130_fd_sc_hd__buf_1 _27834_ (.A(_21489_),
    .X(_21490_));
 sky130_fd_sc_hd__nand3_4 _27835_ (.A(_21488_),
    .B(_21440_),
    .C(_21490_),
    .Y(_21491_));
 sky130_fd_sc_hd__a21o_4 _27836_ (.A1(_21487_),
    .A2(_21491_),
    .B1(_21460_),
    .X(_21492_));
 sky130_fd_sc_hd__buf_1 _27837_ (.A(_18588_),
    .X(_21493_));
 sky130_fd_sc_hd__xor2_4 _27838_ (.A(_21493_),
    .B(_21201_),
    .X(_21494_));
 sky130_fd_sc_hd__nor2_4 _27839_ (.A(_18594_),
    .B(_21192_),
    .Y(_21495_));
 sky130_fd_sc_hd__a2bb2o_4 _27840_ (.A1_N(_21464_),
    .A2_N(_21465_),
    .B1(_18581_),
    .B2(_21185_),
    .X(_21496_));
 sky130_fd_sc_hd__nor2_4 _27841_ (.A(pcpi_rs1[5]),
    .B(_21185_),
    .Y(_21497_));
 sky130_vsdinv _27842_ (.A(_21497_),
    .Y(_21498_));
 sky130_fd_sc_hd__a22oi_4 _27843_ (.A1(pcpi_rs1[6]),
    .A2(_21192_),
    .B1(_21496_),
    .B2(_21498_),
    .Y(_21499_));
 sky130_fd_sc_hd__nor2_4 _27844_ (.A(_21495_),
    .B(_21499_),
    .Y(_21500_));
 sky130_fd_sc_hd__o21ai_4 _27845_ (.A1(_21494_),
    .A2(_21500_),
    .B1(_21428_),
    .Y(_21501_));
 sky130_fd_sc_hd__a21o_4 _27846_ (.A1(_21494_),
    .A2(_21500_),
    .B1(_21501_),
    .X(_21502_));
 sky130_fd_sc_hd__buf_1 _27847_ (.A(_21431_),
    .X(_21503_));
 sky130_fd_sc_hd__a21o_4 _27848_ (.A1(_21492_),
    .A2(_21502_),
    .B1(_21503_),
    .X(_21504_));
 sky130_fd_sc_hd__o21ai_4 _27849_ (.A1(_21486_),
    .A2(_21472_),
    .B1(_21504_),
    .Y(_00559_));
 sky130_vsdinv _27850_ (.A(pcpi_rs1[8]),
    .Y(_21505_));
 sky130_fd_sc_hd__buf_1 _27851_ (.A(_21505_),
    .X(_21506_));
 sky130_fd_sc_hd__buf_1 _27852_ (.A(_18660_),
    .X(_21507_));
 sky130_fd_sc_hd__xnor2_4 _27853_ (.A(_21507_),
    .B(_21207_),
    .Y(_21508_));
 sky130_fd_sc_hd__nand2_4 _27854_ (.A(_18588_),
    .B(_21200_),
    .Y(_21509_));
 sky130_fd_sc_hd__o21ai_4 _27855_ (.A1(_21495_),
    .A2(_21499_),
    .B1(_21509_),
    .Y(_21510_));
 sky130_fd_sc_hd__nor2_4 _27856_ (.A(_18587_),
    .B(_21200_),
    .Y(_21511_));
 sky130_vsdinv _27857_ (.A(_21511_),
    .Y(_21512_));
 sky130_fd_sc_hd__and2_4 _27858_ (.A(_21510_),
    .B(_21512_),
    .X(_21513_));
 sky130_vsdinv _27859_ (.A(_21513_),
    .Y(_21514_));
 sky130_fd_sc_hd__buf_1 _27860_ (.A(_21426_),
    .X(_21515_));
 sky130_fd_sc_hd__a21boi_4 _27861_ (.A1(_21514_),
    .A2(_21508_),
    .B1_N(_21515_),
    .Y(_21516_));
 sky130_fd_sc_hd__o21ai_4 _27862_ (.A1(_21508_),
    .A2(_21514_),
    .B1(_21516_),
    .Y(_21517_));
 sky130_fd_sc_hd__buf_1 _27863_ (.A(_21436_),
    .X(_21518_));
 sky130_fd_sc_hd__buf_1 _27864_ (.A(_20155_),
    .X(_21519_));
 sky130_fd_sc_hd__a2111o_4 _27865_ (.A1(_19829_),
    .A2(_19853_),
    .B1(_21518_),
    .C1(_21519_),
    .D1(_19862_),
    .X(_21520_));
 sky130_fd_sc_hd__buf_1 _27866_ (.A(_21439_),
    .X(_21521_));
 sky130_fd_sc_hd__buf_1 _27867_ (.A(\reg_pc[8] ),
    .X(_21522_));
 sky130_fd_sc_hd__buf_1 _27868_ (.A(_21522_),
    .X(_21523_));
 sky130_fd_sc_hd__nand3_4 _27869_ (.A(_21488_),
    .B(_21521_),
    .C(_21523_),
    .Y(_21524_));
 sky130_fd_sc_hd__buf_1 _27870_ (.A(_18291_),
    .X(_21525_));
 sky130_fd_sc_hd__a21o_4 _27871_ (.A1(_21520_),
    .A2(_21524_),
    .B1(_21525_),
    .X(_21526_));
 sky130_fd_sc_hd__a21o_4 _27872_ (.A1(_21517_),
    .A2(_21526_),
    .B1(_21503_),
    .X(_21527_));
 sky130_fd_sc_hd__o21ai_4 _27873_ (.A1(_21506_),
    .A2(_21472_),
    .B1(_21527_),
    .Y(_00560_));
 sky130_vsdinv _27874_ (.A(_18651_),
    .Y(_21528_));
 sky130_fd_sc_hd__buf_1 _27875_ (.A(_21528_),
    .X(_21529_));
 sky130_fd_sc_hd__buf_1 _27876_ (.A(_18651_),
    .X(_21530_));
 sky130_fd_sc_hd__buf_1 _27877_ (.A(\decoded_imm[9] ),
    .X(_21531_));
 sky130_fd_sc_hd__xor2_4 _27878_ (.A(_21530_),
    .B(_21531_),
    .X(_21532_));
 sky130_fd_sc_hd__nor2_4 _27879_ (.A(pcpi_rs1[8]),
    .B(_21206_),
    .Y(_21533_));
 sky130_fd_sc_hd__a22oi_4 _27880_ (.A1(pcpi_rs1[8]),
    .A2(_21206_),
    .B1(_21510_),
    .B2(_21512_),
    .Y(_21534_));
 sky130_fd_sc_hd__nor2_4 _27881_ (.A(_21533_),
    .B(_21534_),
    .Y(_21535_));
 sky130_fd_sc_hd__buf_1 _27882_ (.A(_21427_),
    .X(_21536_));
 sky130_fd_sc_hd__o21ai_4 _27883_ (.A1(_21532_),
    .A2(_21535_),
    .B1(_21536_),
    .Y(_21537_));
 sky130_fd_sc_hd__a21o_4 _27884_ (.A1(_21532_),
    .A2(_21535_),
    .B1(_21537_),
    .X(_21538_));
 sky130_fd_sc_hd__a2111o_4 _27885_ (.A1(_19888_),
    .A2(_19907_),
    .B1(_21518_),
    .C1(_21519_),
    .D1(_19919_),
    .X(_21539_));
 sky130_fd_sc_hd__buf_1 _27886_ (.A(\reg_pc[9] ),
    .X(_21540_));
 sky130_fd_sc_hd__buf_1 _27887_ (.A(_21540_),
    .X(_21541_));
 sky130_fd_sc_hd__nand3_4 _27888_ (.A(_21488_),
    .B(_21521_),
    .C(_21541_),
    .Y(_21542_));
 sky130_fd_sc_hd__a21o_4 _27889_ (.A1(_21539_),
    .A2(_21542_),
    .B1(_21525_),
    .X(_21543_));
 sky130_fd_sc_hd__a21o_4 _27890_ (.A1(_21538_),
    .A2(_21543_),
    .B1(_21503_),
    .X(_21544_));
 sky130_fd_sc_hd__o21ai_4 _27891_ (.A1(_21529_),
    .A2(_21472_),
    .B1(_21544_),
    .Y(_00561_));
 sky130_fd_sc_hd__buf_1 _27892_ (.A(_18653_),
    .X(_21545_));
 sky130_vsdinv _27893_ (.A(_21545_),
    .Y(_21546_));
 sky130_fd_sc_hd__buf_1 _27894_ (.A(_21395_),
    .X(_21547_));
 sky130_fd_sc_hd__xnor2_4 _27895_ (.A(_21545_),
    .B(_21222_),
    .Y(_21548_));
 sky130_fd_sc_hd__nand2_4 _27896_ (.A(_18650_),
    .B(_21531_),
    .Y(_21549_));
 sky130_fd_sc_hd__o21ai_4 _27897_ (.A1(_21533_),
    .A2(_21534_),
    .B1(_21549_),
    .Y(_21550_));
 sky130_fd_sc_hd__nor2_4 _27898_ (.A(_18650_),
    .B(_21531_),
    .Y(_21551_));
 sky130_vsdinv _27899_ (.A(_21551_),
    .Y(_21552_));
 sky130_fd_sc_hd__and2_4 _27900_ (.A(_21550_),
    .B(_21552_),
    .X(_21553_));
 sky130_vsdinv _27901_ (.A(_21553_),
    .Y(_21554_));
 sky130_fd_sc_hd__a21boi_4 _27902_ (.A1(_21554_),
    .A2(_21548_),
    .B1_N(_21515_),
    .Y(_21555_));
 sky130_fd_sc_hd__o21ai_4 _27903_ (.A1(_21548_),
    .A2(_21554_),
    .B1(_21555_),
    .Y(_21556_));
 sky130_fd_sc_hd__or2_4 _27904_ (.A(_21410_),
    .B(_19975_),
    .X(_21557_));
 sky130_fd_sc_hd__buf_1 _27905_ (.A(\reg_pc[10] ),
    .X(_21558_));
 sky130_fd_sc_hd__buf_1 _27906_ (.A(_21558_),
    .X(_21559_));
 sky130_fd_sc_hd__nand3_4 _27907_ (.A(_21488_),
    .B(_21521_),
    .C(_21559_),
    .Y(_21560_));
 sky130_fd_sc_hd__a21o_4 _27908_ (.A1(_21557_),
    .A2(_21560_),
    .B1(_21525_),
    .X(_21561_));
 sky130_fd_sc_hd__a21o_4 _27909_ (.A1(_21556_),
    .A2(_21561_),
    .B1(_21503_),
    .X(_21562_));
 sky130_fd_sc_hd__o21ai_4 _27910_ (.A1(_21546_),
    .A2(_21547_),
    .B1(_21562_),
    .Y(_00531_));
 sky130_vsdinv _27911_ (.A(_18657_),
    .Y(_21563_));
 sky130_fd_sc_hd__buf_1 _27912_ (.A(_21563_),
    .X(_21564_));
 sky130_fd_sc_hd__buf_1 _27913_ (.A(_18657_),
    .X(_21565_));
 sky130_fd_sc_hd__xor2_4 _27914_ (.A(_21565_),
    .B(_21232_),
    .X(_21566_));
 sky130_fd_sc_hd__nor2_4 _27915_ (.A(_18653_),
    .B(_21221_),
    .Y(_21567_));
 sky130_fd_sc_hd__a22oi_4 _27916_ (.A1(_18653_),
    .A2(_21221_),
    .B1(_21550_),
    .B2(_21552_),
    .Y(_21568_));
 sky130_fd_sc_hd__nor2_4 _27917_ (.A(_21567_),
    .B(_21568_),
    .Y(_21569_));
 sky130_fd_sc_hd__o21ai_4 _27918_ (.A1(_21566_),
    .A2(_21569_),
    .B1(_21536_),
    .Y(_21570_));
 sky130_fd_sc_hd__a21o_4 _27919_ (.A1(_21566_),
    .A2(_21569_),
    .B1(_21570_),
    .X(_21571_));
 sky130_fd_sc_hd__a2111o_4 _27920_ (.A1(_20004_),
    .A2(_20028_),
    .B1(_21518_),
    .C1(_21519_),
    .D1(_20049_),
    .X(_21572_));
 sky130_fd_sc_hd__buf_1 _27921_ (.A(_21413_),
    .X(_21573_));
 sky130_fd_sc_hd__buf_1 _27922_ (.A(\reg_pc[11] ),
    .X(_21574_));
 sky130_fd_sc_hd__nand3_4 _27923_ (.A(_21573_),
    .B(_21521_),
    .C(_21574_),
    .Y(_21575_));
 sky130_fd_sc_hd__a21o_4 _27924_ (.A1(_21572_),
    .A2(_21575_),
    .B1(_21525_),
    .X(_21576_));
 sky130_fd_sc_hd__buf_1 _27925_ (.A(_21431_),
    .X(_21577_));
 sky130_fd_sc_hd__a21o_4 _27926_ (.A1(_21571_),
    .A2(_21576_),
    .B1(_21577_),
    .X(_21578_));
 sky130_fd_sc_hd__o21ai_4 _27927_ (.A1(_21564_),
    .A2(_21547_),
    .B1(_21578_),
    .Y(_00532_));
 sky130_vsdinv _27928_ (.A(_18646_),
    .Y(_21579_));
 sky130_fd_sc_hd__buf_1 _27929_ (.A(_21579_),
    .X(_21580_));
 sky130_fd_sc_hd__buf_1 _27930_ (.A(_21394_),
    .X(_21581_));
 sky130_fd_sc_hd__buf_1 _27931_ (.A(_21581_),
    .X(_21582_));
 sky130_fd_sc_hd__buf_1 _27932_ (.A(_19097_),
    .X(_21583_));
 sky130_fd_sc_hd__buf_1 _27933_ (.A(_21355_),
    .X(_21584_));
 sky130_fd_sc_hd__buf_1 _27934_ (.A(_21359_),
    .X(_21585_));
 sky130_fd_sc_hd__buf_1 _27935_ (.A(\reg_pc[12] ),
    .X(_21586_));
 sky130_fd_sc_hd__buf_1 _27936_ (.A(_21586_),
    .X(_21587_));
 sky130_fd_sc_hd__nand3_4 _27937_ (.A(_21585_),
    .B(_21416_),
    .C(_21587_),
    .Y(_21588_));
 sky130_fd_sc_hd__o21ai_4 _27938_ (.A1(_21584_),
    .A2(_20111_),
    .B1(_21588_),
    .Y(_21589_));
 sky130_fd_sc_hd__buf_1 _27939_ (.A(_18646_),
    .X(_21590_));
 sky130_fd_sc_hd__xnor2_4 _27940_ (.A(_21590_),
    .B(_21239_),
    .Y(_21591_));
 sky130_fd_sc_hd__nand2_4 _27941_ (.A(_18656_),
    .B(_21232_),
    .Y(_21592_));
 sky130_fd_sc_hd__o21ai_4 _27942_ (.A1(_21567_),
    .A2(_21568_),
    .B1(_21592_),
    .Y(_21593_));
 sky130_fd_sc_hd__nor2_4 _27943_ (.A(_18656_),
    .B(\decoded_imm[11] ),
    .Y(_21594_));
 sky130_vsdinv _27944_ (.A(_21594_),
    .Y(_21595_));
 sky130_fd_sc_hd__nand2_4 _27945_ (.A(_21593_),
    .B(_21595_),
    .Y(_21596_));
 sky130_fd_sc_hd__buf_1 _27946_ (.A(_21427_),
    .X(_21597_));
 sky130_fd_sc_hd__o21ai_4 _27947_ (.A1(_21591_),
    .A2(_21596_),
    .B1(_21597_),
    .Y(_21598_));
 sky130_fd_sc_hd__a21oi_4 _27948_ (.A1(_21591_),
    .A2(_21596_),
    .B1(_21598_),
    .Y(_21599_));
 sky130_fd_sc_hd__a21o_4 _27949_ (.A1(_21583_),
    .A2(_21589_),
    .B1(_21599_),
    .X(_21600_));
 sky130_fd_sc_hd__a2bb2o_4 _27950_ (.A1_N(_21580_),
    .A2_N(_21582_),
    .B1(_21335_),
    .B2(_21600_),
    .X(_00533_));
 sky130_fd_sc_hd__buf_1 _27951_ (.A(_18640_),
    .X(_21601_));
 sky130_vsdinv _27952_ (.A(_21601_),
    .Y(_21602_));
 sky130_fd_sc_hd__buf_1 _27953_ (.A(\decoded_imm[13] ),
    .X(_21603_));
 sky130_fd_sc_hd__nor2_4 _27954_ (.A(_18640_),
    .B(_21603_),
    .Y(_21604_));
 sky130_fd_sc_hd__buf_1 _27955_ (.A(_21601_),
    .X(_21605_));
 sky130_fd_sc_hd__nand2_4 _27956_ (.A(_21605_),
    .B(_21603_),
    .Y(_21606_));
 sky130_vsdinv _27957_ (.A(_21606_),
    .Y(_21607_));
 sky130_fd_sc_hd__nor2_4 _27958_ (.A(_21604_),
    .B(_21607_),
    .Y(_21608_));
 sky130_fd_sc_hd__nand2_4 _27959_ (.A(_18645_),
    .B(_21238_),
    .Y(_21609_));
 sky130_fd_sc_hd__nor2_4 _27960_ (.A(_18645_),
    .B(_21238_),
    .Y(_21610_));
 sky130_fd_sc_hd__a21oi_4 _27961_ (.A1(_21596_),
    .A2(_21609_),
    .B1(_21610_),
    .Y(_21611_));
 sky130_fd_sc_hd__a21boi_4 _27962_ (.A1(_21611_),
    .A2(_21608_),
    .B1_N(_21515_),
    .Y(_21612_));
 sky130_fd_sc_hd__o21ai_4 _27963_ (.A1(_21608_),
    .A2(_21611_),
    .B1(_21612_),
    .Y(_21613_));
 sky130_fd_sc_hd__buf_1 _27964_ (.A(_20102_),
    .X(_21614_));
 sky130_fd_sc_hd__a2111o_4 _27965_ (.A1(_20134_),
    .A2(_20154_),
    .B1(_21518_),
    .C1(_21614_),
    .D1(_20169_),
    .X(_21615_));
 sky130_fd_sc_hd__buf_1 _27966_ (.A(_21439_),
    .X(_21616_));
 sky130_fd_sc_hd__buf_1 _27967_ (.A(\reg_pc[13] ),
    .X(_21617_));
 sky130_fd_sc_hd__nand3_4 _27968_ (.A(_21573_),
    .B(_21616_),
    .C(_21617_),
    .Y(_21618_));
 sky130_fd_sc_hd__buf_1 _27969_ (.A(_21115_),
    .X(_21619_));
 sky130_fd_sc_hd__a21o_4 _27970_ (.A1(_21615_),
    .A2(_21618_),
    .B1(_21619_),
    .X(_21620_));
 sky130_fd_sc_hd__a21o_4 _27971_ (.A1(_21613_),
    .A2(_21620_),
    .B1(_21577_),
    .X(_21621_));
 sky130_fd_sc_hd__o21ai_4 _27972_ (.A1(_21602_),
    .A2(_21547_),
    .B1(_21621_),
    .Y(_00534_));
 sky130_vsdinv _27973_ (.A(_18638_),
    .Y(_21622_));
 sky130_vsdinv _27974_ (.A(_21604_),
    .Y(_21623_));
 sky130_fd_sc_hd__nand2_4 _27975_ (.A(_18637_),
    .B(_21253_),
    .Y(_21624_));
 sky130_fd_sc_hd__buf_1 _27976_ (.A(_21624_),
    .X(_21625_));
 sky130_fd_sc_hd__nor2_4 _27977_ (.A(_18637_),
    .B(_21253_),
    .Y(_21626_));
 sky130_vsdinv _27978_ (.A(_21626_),
    .Y(_21627_));
 sky130_fd_sc_hd__a21o_4 _27979_ (.A1(_18640_),
    .A2(_21603_),
    .B1(_21611_),
    .X(_21628_));
 sky130_fd_sc_hd__o21ai_4 _27980_ (.A1(_21607_),
    .A2(_21611_),
    .B1(_21623_),
    .Y(_21629_));
 sky130_fd_sc_hd__a21bo_4 _27981_ (.A1(_21625_),
    .A2(_21627_),
    .B1_N(_21629_),
    .X(_21630_));
 sky130_fd_sc_hd__nand2_4 _27982_ (.A(_21630_),
    .B(_21451_),
    .Y(_21631_));
 sky130_fd_sc_hd__a41o_4 _27983_ (.A1(_21623_),
    .A2(_21625_),
    .A3(_21627_),
    .A4(_21628_),
    .B1(_21631_),
    .X(_21632_));
 sky130_fd_sc_hd__buf_1 _27984_ (.A(_21436_),
    .X(_21633_));
 sky130_fd_sc_hd__a2111o_4 _27985_ (.A1(_20201_),
    .A2(_20218_),
    .B1(_21633_),
    .C1(_21614_),
    .D1(_20225_),
    .X(_21634_));
 sky130_fd_sc_hd__buf_1 _27986_ (.A(\reg_pc[14] ),
    .X(_21635_));
 sky130_fd_sc_hd__nand3_4 _27987_ (.A(_21573_),
    .B(_21616_),
    .C(_21635_),
    .Y(_21636_));
 sky130_fd_sc_hd__a21o_4 _27988_ (.A1(_21634_),
    .A2(_21636_),
    .B1(_21619_),
    .X(_21637_));
 sky130_fd_sc_hd__a21o_4 _27989_ (.A1(_21632_),
    .A2(_21637_),
    .B1(_21577_),
    .X(_21638_));
 sky130_fd_sc_hd__o21ai_4 _27990_ (.A1(_21622_),
    .A2(_21547_),
    .B1(_21638_),
    .Y(_00535_));
 sky130_vsdinv _27991_ (.A(_18642_),
    .Y(_21639_));
 sky130_fd_sc_hd__buf_1 _27992_ (.A(_21639_),
    .X(_21640_));
 sky130_fd_sc_hd__buf_1 _27993_ (.A(_21581_),
    .X(_21641_));
 sky130_fd_sc_hd__and2_4 _27994_ (.A(_21629_),
    .B(_21625_),
    .X(_21642_));
 sky130_fd_sc_hd__xor2_4 _27995_ (.A(pcpi_rs1[15]),
    .B(_21258_),
    .X(_21643_));
 sky130_vsdinv _27996_ (.A(_21643_),
    .Y(_21644_));
 sky130_fd_sc_hd__o21ai_4 _27997_ (.A1(_21626_),
    .A2(_21642_),
    .B1(_21644_),
    .Y(_21645_));
 sky130_fd_sc_hd__a211o_4 _27998_ (.A1(_21629_),
    .A2(_21625_),
    .B1(_21626_),
    .C1(_21644_),
    .X(_21646_));
 sky130_fd_sc_hd__nand3_4 _27999_ (.A(_21645_),
    .B(_21646_),
    .C(_21597_),
    .Y(_21647_));
 sky130_fd_sc_hd__a2111o_4 _28000_ (.A1(_20251_),
    .A2(_20266_),
    .B1(_21633_),
    .C1(_21614_),
    .D1(_20274_),
    .X(_21648_));
 sky130_fd_sc_hd__buf_1 _28001_ (.A(\reg_pc[15] ),
    .X(_21649_));
 sky130_fd_sc_hd__buf_1 _28002_ (.A(_21649_),
    .X(_21650_));
 sky130_fd_sc_hd__nand3_4 _28003_ (.A(_21573_),
    .B(_21616_),
    .C(_21650_),
    .Y(_21651_));
 sky130_fd_sc_hd__a21o_4 _28004_ (.A1(_21648_),
    .A2(_21651_),
    .B1(_21619_),
    .X(_21652_));
 sky130_fd_sc_hd__a21o_4 _28005_ (.A1(_21647_),
    .A2(_21652_),
    .B1(_21577_),
    .X(_21653_));
 sky130_fd_sc_hd__o21ai_4 _28006_ (.A1(_21640_),
    .A2(_21641_),
    .B1(_21653_),
    .Y(_00536_));
 sky130_vsdinv _28007_ (.A(_18710_),
    .Y(_21654_));
 sky130_fd_sc_hd__xor2_4 _28008_ (.A(pcpi_rs1[16]),
    .B(_21263_),
    .X(_21655_));
 sky130_fd_sc_hd__and3_4 _28009_ (.A(_21643_),
    .B(_21624_),
    .C(_21627_),
    .X(_21656_));
 sky130_fd_sc_hd__nand3_4 _28010_ (.A(_21628_),
    .B(_21623_),
    .C(_21656_),
    .Y(_21657_));
 sky130_fd_sc_hd__maj3_4 _28011_ (.A(_21639_),
    .B(_21624_),
    .C(_21259_),
    .X(_21658_));
 sky130_fd_sc_hd__nand2_4 _28012_ (.A(_21657_),
    .B(_21658_),
    .Y(_21659_));
 sky130_fd_sc_hd__a21boi_4 _28013_ (.A1(_21659_),
    .A2(_21655_),
    .B1_N(_21515_),
    .Y(_21660_));
 sky130_fd_sc_hd__o21ai_4 _28014_ (.A1(_21655_),
    .A2(_21659_),
    .B1(_21660_),
    .Y(_21661_));
 sky130_fd_sc_hd__a2111o_4 _28015_ (.A1(_20297_),
    .A2(_20317_),
    .B1(_21633_),
    .C1(_21614_),
    .D1(_20325_),
    .X(_21662_));
 sky130_fd_sc_hd__buf_1 _28016_ (.A(_21413_),
    .X(_21663_));
 sky130_fd_sc_hd__buf_1 _28017_ (.A(\reg_pc[16] ),
    .X(_21664_));
 sky130_fd_sc_hd__buf_1 _28018_ (.A(_21664_),
    .X(_21665_));
 sky130_fd_sc_hd__nand3_4 _28019_ (.A(_21663_),
    .B(_21616_),
    .C(_21665_),
    .Y(_21666_));
 sky130_fd_sc_hd__a21o_4 _28020_ (.A1(_21662_),
    .A2(_21666_),
    .B1(_21619_),
    .X(_21667_));
 sky130_fd_sc_hd__buf_1 _28021_ (.A(_21431_),
    .X(_21668_));
 sky130_fd_sc_hd__a21o_4 _28022_ (.A1(_21661_),
    .A2(_21667_),
    .B1(_21668_),
    .X(_21669_));
 sky130_fd_sc_hd__o21ai_4 _28023_ (.A1(_21654_),
    .A2(_21641_),
    .B1(_21669_),
    .Y(_00537_));
 sky130_vsdinv _28024_ (.A(pcpi_rs1[17]),
    .Y(_21670_));
 sky130_fd_sc_hd__buf_1 _28025_ (.A(_21670_),
    .X(_21671_));
 sky130_fd_sc_hd__a2111o_4 _28026_ (.A1(_20351_),
    .A2(_20365_),
    .B1(_21383_),
    .C1(_21356_),
    .D1(_20373_),
    .X(_21672_));
 sky130_fd_sc_hd__buf_1 _28027_ (.A(_21359_),
    .X(_21673_));
 sky130_fd_sc_hd__buf_1 _28028_ (.A(\reg_pc[17] ),
    .X(_21674_));
 sky130_fd_sc_hd__nand3_4 _28029_ (.A(_21673_),
    .B(_21362_),
    .C(_21674_),
    .Y(_21675_));
 sky130_fd_sc_hd__a21oi_4 _28030_ (.A1(_21672_),
    .A2(_21675_),
    .B1(_21386_),
    .Y(_21676_));
 sky130_fd_sc_hd__xor2_4 _28031_ (.A(_18714_),
    .B(_21270_),
    .X(_21677_));
 sky130_fd_sc_hd__buf_1 _28032_ (.A(_18710_),
    .X(_21678_));
 sky130_fd_sc_hd__maj3_4 _28033_ (.A(_21678_),
    .B(_21659_),
    .C(_21264_),
    .X(_21679_));
 sky130_fd_sc_hd__a22oi_4 _28034_ (.A1(_18246_),
    .A2(\cpu_state[5] ),
    .B1(_18237_),
    .B2(_18239_),
    .Y(_21680_));
 sky130_fd_sc_hd__nor2_4 _28035_ (.A(_21680_),
    .B(_18258_),
    .Y(_21681_));
 sky130_fd_sc_hd__buf_1 _28036_ (.A(_21681_),
    .X(_21682_));
 sky130_fd_sc_hd__o21ai_4 _28037_ (.A1(_21677_),
    .A2(_21679_),
    .B1(_21682_),
    .Y(_21683_));
 sky130_fd_sc_hd__a21oi_4 _28038_ (.A1(_21677_),
    .A2(_21679_),
    .B1(_21683_),
    .Y(_21684_));
 sky130_fd_sc_hd__buf_1 _28039_ (.A(_21346_),
    .X(_21685_));
 sky130_fd_sc_hd__o21ai_4 _28040_ (.A1(_21676_),
    .A2(_21684_),
    .B1(_21685_),
    .Y(_21686_));
 sky130_fd_sc_hd__o21ai_4 _28041_ (.A1(_21671_),
    .A2(_21641_),
    .B1(_21686_),
    .Y(_00538_));
 sky130_fd_sc_hd__buf_1 _28042_ (.A(_18701_),
    .X(_21687_));
 sky130_fd_sc_hd__xor2_4 _28043_ (.A(_18700_),
    .B(_21274_),
    .X(_21688_));
 sky130_vsdinv _28044_ (.A(_21688_),
    .Y(_21689_));
 sky130_fd_sc_hd__and2_4 _28045_ (.A(_21677_),
    .B(_21655_),
    .X(_21690_));
 sky130_fd_sc_hd__nand2_4 _28046_ (.A(_18709_),
    .B(_21263_),
    .Y(_21691_));
 sky130_vsdinv _28047_ (.A(_21691_),
    .Y(_21692_));
 sky130_fd_sc_hd__maj3_4 _28048_ (.A(_18714_),
    .B(_21692_),
    .C(_21270_),
    .X(_21693_));
 sky130_fd_sc_hd__a21oi_4 _28049_ (.A1(_21659_),
    .A2(_21690_),
    .B1(_21693_),
    .Y(_21694_));
 sky130_fd_sc_hd__o21ai_4 _28050_ (.A1(_21689_),
    .A2(_21694_),
    .B1(_21536_),
    .Y(_21695_));
 sky130_fd_sc_hd__a21o_4 _28051_ (.A1(_21689_),
    .A2(_21694_),
    .B1(_21695_),
    .X(_21696_));
 sky130_fd_sc_hd__buf_1 _28052_ (.A(_20155_),
    .X(_21697_));
 sky130_fd_sc_hd__a2111o_4 _28053_ (.A1(_20406_),
    .A2(_20420_),
    .B1(_21633_),
    .C1(_21697_),
    .D1(_20427_),
    .X(_21698_));
 sky130_fd_sc_hd__buf_1 _28054_ (.A(_21439_),
    .X(_21699_));
 sky130_fd_sc_hd__buf_1 _28055_ (.A(\reg_pc[18] ),
    .X(_21700_));
 sky130_fd_sc_hd__buf_1 _28056_ (.A(_21700_),
    .X(_21701_));
 sky130_fd_sc_hd__nand3_4 _28057_ (.A(_21663_),
    .B(_21699_),
    .C(_21701_),
    .Y(_21702_));
 sky130_fd_sc_hd__buf_1 _28058_ (.A(_21115_),
    .X(_21703_));
 sky130_fd_sc_hd__a21o_4 _28059_ (.A1(_21698_),
    .A2(_21702_),
    .B1(_21703_),
    .X(_21704_));
 sky130_fd_sc_hd__a21o_4 _28060_ (.A1(_21696_),
    .A2(_21704_),
    .B1(_21668_),
    .X(_21705_));
 sky130_fd_sc_hd__o21ai_4 _28061_ (.A1(_21687_),
    .A2(_21641_),
    .B1(_21705_),
    .Y(_00539_));
 sky130_vsdinv _28062_ (.A(_18693_),
    .Y(_21706_));
 sky130_fd_sc_hd__buf_1 _28063_ (.A(_21706_),
    .X(_21707_));
 sky130_fd_sc_hd__buf_1 _28064_ (.A(_21685_),
    .X(_21708_));
 sky130_fd_sc_hd__xor2_4 _28065_ (.A(_18693_),
    .B(_21281_),
    .X(_21709_));
 sky130_vsdinv _28066_ (.A(_21709_),
    .Y(_21710_));
 sky130_fd_sc_hd__maj3_4 _28067_ (.A(_21687_),
    .B(_21694_),
    .C(_21275_),
    .X(_21711_));
 sky130_fd_sc_hd__nor2_4 _28068_ (.A(_21710_),
    .B(_21711_),
    .Y(_21712_));
 sky130_vsdinv _28069_ (.A(_21681_),
    .Y(_21713_));
 sky130_fd_sc_hd__a21o_4 _28070_ (.A1(_21711_),
    .A2(_21710_),
    .B1(_21713_),
    .X(_21714_));
 sky130_fd_sc_hd__buf_1 _28071_ (.A(_21415_),
    .X(_21715_));
 sky130_fd_sc_hd__buf_1 _28072_ (.A(\reg_pc[19] ),
    .X(_21716_));
 sky130_fd_sc_hd__buf_1 _28073_ (.A(_21716_),
    .X(_21717_));
 sky130_fd_sc_hd__nand3_4 _28074_ (.A(_21673_),
    .B(_21715_),
    .C(_21717_),
    .Y(_21718_));
 sky130_fd_sc_hd__o21ai_4 _28075_ (.A1(_21584_),
    .A2(_20478_),
    .B1(_21718_),
    .Y(_21719_));
 sky130_fd_sc_hd__a2bb2o_4 _28076_ (.A1_N(_21712_),
    .A2_N(_21714_),
    .B1(_21583_),
    .B2(_21719_),
    .X(_21720_));
 sky130_fd_sc_hd__a2bb2o_4 _28077_ (.A1_N(_21707_),
    .A2_N(_21582_),
    .B1(_21708_),
    .B2(_21720_),
    .X(_00540_));
 sky130_fd_sc_hd__buf_1 _28078_ (.A(_18666_),
    .X(_21721_));
 sky130_vsdinv _28079_ (.A(_21721_),
    .Y(_21722_));
 sky130_fd_sc_hd__buf_1 _28080_ (.A(_21581_),
    .X(_21723_));
 sky130_fd_sc_hd__xor2_4 _28081_ (.A(pcpi_rs1[20]),
    .B(\decoded_imm[20] ),
    .X(_21724_));
 sky130_fd_sc_hd__a21boi_4 _28082_ (.A1(_21657_),
    .A2(_21658_),
    .B1_N(_21690_),
    .Y(_21725_));
 sky130_fd_sc_hd__and2_4 _28083_ (.A(_21688_),
    .B(_21709_),
    .X(_21726_));
 sky130_fd_sc_hd__o21ai_4 _28084_ (.A1(_21693_),
    .A2(_21725_),
    .B1(_21726_),
    .Y(_21727_));
 sky130_fd_sc_hd__nand2_4 _28085_ (.A(_18700_),
    .B(_21274_),
    .Y(_21728_));
 sky130_fd_sc_hd__maj3_4 _28086_ (.A(_21706_),
    .B(_21728_),
    .C(_21282_),
    .X(_21729_));
 sky130_fd_sc_hd__nand2_4 _28087_ (.A(_21727_),
    .B(_21729_),
    .Y(_21730_));
 sky130_fd_sc_hd__a21boi_4 _28088_ (.A1(_21730_),
    .A2(_21724_),
    .B1_N(_21451_),
    .Y(_21731_));
 sky130_fd_sc_hd__o21ai_4 _28089_ (.A1(_21724_),
    .A2(_21730_),
    .B1(_21731_),
    .Y(_21732_));
 sky130_fd_sc_hd__buf_1 _28090_ (.A(_21436_),
    .X(_21733_));
 sky130_fd_sc_hd__a2111o_4 _28091_ (.A1(_20500_),
    .A2(_20514_),
    .B1(_21733_),
    .C1(_21697_),
    .D1(_20524_),
    .X(_21734_));
 sky130_fd_sc_hd__buf_1 _28092_ (.A(\reg_pc[20] ),
    .X(_21735_));
 sky130_fd_sc_hd__nand3_4 _28093_ (.A(_21663_),
    .B(_21699_),
    .C(_21735_),
    .Y(_21736_));
 sky130_fd_sc_hd__a21o_4 _28094_ (.A1(_21734_),
    .A2(_21736_),
    .B1(_21703_),
    .X(_21737_));
 sky130_fd_sc_hd__a21o_4 _28095_ (.A1(_21732_),
    .A2(_21737_),
    .B1(_21668_),
    .X(_21738_));
 sky130_fd_sc_hd__o21ai_4 _28096_ (.A1(_21722_),
    .A2(_21723_),
    .B1(_21738_),
    .Y(_00542_));
 sky130_fd_sc_hd__buf_1 _28097_ (.A(_18680_),
    .X(_21739_));
 sky130_vsdinv _28098_ (.A(_21739_),
    .Y(_21740_));
 sky130_fd_sc_hd__a2111o_4 _28099_ (.A1(_20551_),
    .A2(_20565_),
    .B1(_21383_),
    .C1(_21356_),
    .D1(_20572_),
    .X(_21741_));
 sky130_fd_sc_hd__buf_1 _28100_ (.A(\reg_pc[21] ),
    .X(_21742_));
 sky130_fd_sc_hd__buf_1 _28101_ (.A(_21742_),
    .X(_21743_));
 sky130_fd_sc_hd__nand3_4 _28102_ (.A(_21673_),
    .B(_21715_),
    .C(_21743_),
    .Y(_21744_));
 sky130_fd_sc_hd__a21oi_4 _28103_ (.A1(_21741_),
    .A2(_21744_),
    .B1(_21386_),
    .Y(_21745_));
 sky130_fd_sc_hd__xor2_4 _28104_ (.A(pcpi_rs1[21]),
    .B(\decoded_imm[21] ),
    .X(_21746_));
 sky130_fd_sc_hd__maj3_4 _28105_ (.A(_21721_),
    .B(_21730_),
    .C(_21286_),
    .X(_21747_));
 sky130_fd_sc_hd__o21ai_4 _28106_ (.A1(_21746_),
    .A2(_21747_),
    .B1(_21682_),
    .Y(_21748_));
 sky130_fd_sc_hd__a21oi_4 _28107_ (.A1(_21746_),
    .A2(_21747_),
    .B1(_21748_),
    .Y(_21749_));
 sky130_fd_sc_hd__o21ai_4 _28108_ (.A1(_21745_),
    .A2(_21749_),
    .B1(_21685_),
    .Y(_21750_));
 sky130_fd_sc_hd__o21ai_4 _28109_ (.A1(_21740_),
    .A2(_21723_),
    .B1(_21750_),
    .Y(_00543_));
 sky130_fd_sc_hd__buf_1 _28110_ (.A(_18673_),
    .X(_21751_));
 sky130_fd_sc_hd__xor2_4 _28111_ (.A(pcpi_rs1[22]),
    .B(\decoded_imm[22] ),
    .X(_21752_));
 sky130_vsdinv _28112_ (.A(_21752_),
    .Y(_21753_));
 sky130_fd_sc_hd__and2_4 _28113_ (.A(_21746_),
    .B(_21724_),
    .X(_21754_));
 sky130_fd_sc_hd__nand2_4 _28114_ (.A(_18665_),
    .B(_21286_),
    .Y(_21755_));
 sky130_vsdinv _28115_ (.A(_21755_),
    .Y(_21756_));
 sky130_fd_sc_hd__maj3_4 _28116_ (.A(pcpi_rs1[21]),
    .B(_21756_),
    .C(_21292_),
    .X(_21757_));
 sky130_fd_sc_hd__a21oi_4 _28117_ (.A1(_21730_),
    .A2(_21754_),
    .B1(_21757_),
    .Y(_21758_));
 sky130_fd_sc_hd__o21ai_4 _28118_ (.A1(_21753_),
    .A2(_21758_),
    .B1(_21536_),
    .Y(_21759_));
 sky130_fd_sc_hd__a21o_4 _28119_ (.A1(_21753_),
    .A2(_21758_),
    .B1(_21759_),
    .X(_21760_));
 sky130_fd_sc_hd__or2_4 _28120_ (.A(_21410_),
    .B(_20617_),
    .X(_21761_));
 sky130_fd_sc_hd__buf_1 _28121_ (.A(\reg_pc[22] ),
    .X(_21762_));
 sky130_fd_sc_hd__nand3_4 _28122_ (.A(_21663_),
    .B(_21699_),
    .C(_21762_),
    .Y(_21763_));
 sky130_fd_sc_hd__a21o_4 _28123_ (.A1(_21761_),
    .A2(_21763_),
    .B1(_21703_),
    .X(_21764_));
 sky130_fd_sc_hd__a21o_4 _28124_ (.A1(_21760_),
    .A2(_21764_),
    .B1(_21668_),
    .X(_21765_));
 sky130_fd_sc_hd__o21ai_4 _28125_ (.A1(_21751_),
    .A2(_21723_),
    .B1(_21765_),
    .Y(_00544_));
 sky130_vsdinv _28126_ (.A(pcpi_rs1[23]),
    .Y(_21766_));
 sky130_fd_sc_hd__xor2_4 _28127_ (.A(pcpi_rs1[23]),
    .B(\decoded_imm[23] ),
    .X(_21767_));
 sky130_vsdinv _28128_ (.A(_21767_),
    .Y(_21768_));
 sky130_fd_sc_hd__maj3_4 _28129_ (.A(_21751_),
    .B(_21758_),
    .C(_21297_),
    .X(_21769_));
 sky130_fd_sc_hd__nor2_4 _28130_ (.A(_21768_),
    .B(_21769_),
    .Y(_21770_));
 sky130_fd_sc_hd__a21o_4 _28131_ (.A1(_21769_),
    .A2(_21768_),
    .B1(_21713_),
    .X(_21771_));
 sky130_fd_sc_hd__buf_1 _28132_ (.A(\reg_pc[23] ),
    .X(_21772_));
 sky130_fd_sc_hd__nand3_4 _28133_ (.A(_21585_),
    .B(_21715_),
    .C(_21772_),
    .Y(_21773_));
 sky130_fd_sc_hd__o21ai_4 _28134_ (.A1(_21584_),
    .A2(_20657_),
    .B1(_21773_),
    .Y(_21774_));
 sky130_fd_sc_hd__a2bb2o_4 _28135_ (.A1_N(_21770_),
    .A2_N(_21771_),
    .B1(_21184_),
    .B2(_21774_),
    .X(_21775_));
 sky130_fd_sc_hd__a2bb2o_4 _28136_ (.A1_N(_21766_),
    .A2_N(_21582_),
    .B1(_21708_),
    .B2(_21775_),
    .X(_00545_));
 sky130_fd_sc_hd__xor2_4 _28137_ (.A(pcpi_rs1[24]),
    .B(\decoded_imm[24] ),
    .X(_21776_));
 sky130_vsdinv _28138_ (.A(_21754_),
    .Y(_21777_));
 sky130_fd_sc_hd__a21oi_4 _28139_ (.A1(_21727_),
    .A2(_21729_),
    .B1(_21777_),
    .Y(_21778_));
 sky130_fd_sc_hd__and2_4 _28140_ (.A(_21752_),
    .B(_21767_),
    .X(_21779_));
 sky130_fd_sc_hd__o21ai_4 _28141_ (.A1(_21757_),
    .A2(_21778_),
    .B1(_21779_),
    .Y(_21780_));
 sky130_fd_sc_hd__nand2_4 _28142_ (.A(_18672_),
    .B(_21296_),
    .Y(_21781_));
 sky130_fd_sc_hd__maj3_4 _28143_ (.A(_21766_),
    .B(_21781_),
    .C(_21301_),
    .X(_21782_));
 sky130_fd_sc_hd__nand2_4 _28144_ (.A(_21780_),
    .B(_21782_),
    .Y(_21783_));
 sky130_fd_sc_hd__a21boi_4 _28145_ (.A1(_21783_),
    .A2(_21776_),
    .B1_N(_21451_),
    .Y(_21784_));
 sky130_fd_sc_hd__o21ai_4 _28146_ (.A1(_21776_),
    .A2(_21783_),
    .B1(_21784_),
    .Y(_21785_));
 sky130_fd_sc_hd__a2111o_4 _28147_ (.A1(_20679_),
    .A2(_20694_),
    .B1(_21733_),
    .C1(_21697_),
    .D1(_20702_),
    .X(_21786_));
 sky130_fd_sc_hd__buf_1 _28148_ (.A(_21358_),
    .X(_21787_));
 sky130_fd_sc_hd__buf_1 _28149_ (.A(\reg_pc[24] ),
    .X(_21788_));
 sky130_fd_sc_hd__nand3_4 _28150_ (.A(_21787_),
    .B(_21699_),
    .C(_21788_),
    .Y(_21789_));
 sky130_fd_sc_hd__a21o_4 _28151_ (.A1(_21786_),
    .A2(_21789_),
    .B1(_21703_),
    .X(_21790_));
 sky130_fd_sc_hd__buf_1 _28152_ (.A(_19494_),
    .X(_21791_));
 sky130_fd_sc_hd__a21o_4 _28153_ (.A1(_21785_),
    .A2(_21790_),
    .B1(_21791_),
    .X(_21792_));
 sky130_fd_sc_hd__o21ai_4 _28154_ (.A1(_18728_),
    .A2(_21723_),
    .B1(_21792_),
    .Y(_00546_));
 sky130_vsdinv _28155_ (.A(_18765_),
    .Y(_21793_));
 sky130_fd_sc_hd__buf_1 _28156_ (.A(_21581_),
    .X(_21794_));
 sky130_fd_sc_hd__a2111o_4 _28157_ (.A1(_20727_),
    .A2(_20742_),
    .B1(_21355_),
    .C1(_21356_),
    .D1(_20749_),
    .X(_21795_));
 sky130_fd_sc_hd__buf_1 _28158_ (.A(\reg_pc[25] ),
    .X(_21796_));
 sky130_fd_sc_hd__nand3_4 _28159_ (.A(_21673_),
    .B(_21715_),
    .C(_21796_),
    .Y(_21797_));
 sky130_fd_sc_hd__a21oi_4 _28160_ (.A1(_21795_),
    .A2(_21797_),
    .B1(_18292_),
    .Y(_21798_));
 sky130_fd_sc_hd__xor2_4 _28161_ (.A(pcpi_rs1[25]),
    .B(\decoded_imm[25] ),
    .X(_21799_));
 sky130_fd_sc_hd__maj3_4 _28162_ (.A(_18732_),
    .B(_21783_),
    .C(_21305_),
    .X(_21800_));
 sky130_fd_sc_hd__o21ai_4 _28163_ (.A1(_21799_),
    .A2(_21800_),
    .B1(_21682_),
    .Y(_21801_));
 sky130_fd_sc_hd__a21oi_4 _28164_ (.A1(_21799_),
    .A2(_21800_),
    .B1(_21801_),
    .Y(_21802_));
 sky130_fd_sc_hd__o21ai_4 _28165_ (.A1(_21798_),
    .A2(_21802_),
    .B1(_21685_),
    .Y(_21803_));
 sky130_fd_sc_hd__o21ai_4 _28166_ (.A1(_21793_),
    .A2(_21794_),
    .B1(_21803_),
    .Y(_00547_));
 sky130_vsdinv _28167_ (.A(_18724_),
    .Y(_21804_));
 sky130_fd_sc_hd__xor2_4 _28168_ (.A(pcpi_rs1[26]),
    .B(\decoded_imm[26] ),
    .X(_21805_));
 sky130_vsdinv _28169_ (.A(_21805_),
    .Y(_21806_));
 sky130_fd_sc_hd__and2_4 _28170_ (.A(_21799_),
    .B(_21776_),
    .X(_21807_));
 sky130_fd_sc_hd__nand2_4 _28171_ (.A(pcpi_rs1[24]),
    .B(\decoded_imm[24] ),
    .Y(_21808_));
 sky130_vsdinv _28172_ (.A(_21808_),
    .Y(_21809_));
 sky130_fd_sc_hd__maj3_4 _28173_ (.A(_18764_),
    .B(_21809_),
    .C(_21311_),
    .X(_21810_));
 sky130_fd_sc_hd__a21oi_4 _28174_ (.A1(_21783_),
    .A2(_21807_),
    .B1(_21810_),
    .Y(_21811_));
 sky130_fd_sc_hd__o21ai_4 _28175_ (.A1(_21806_),
    .A2(_21811_),
    .B1(_21428_),
    .Y(_21812_));
 sky130_fd_sc_hd__a21o_4 _28176_ (.A1(_21806_),
    .A2(_21811_),
    .B1(_21812_),
    .X(_21813_));
 sky130_fd_sc_hd__a2111o_4 _28177_ (.A1(_20770_),
    .A2(_20784_),
    .B1(_21733_),
    .C1(_21697_),
    .D1(_20792_),
    .X(_21814_));
 sky130_fd_sc_hd__buf_1 _28178_ (.A(_18795_),
    .X(_21815_));
 sky130_fd_sc_hd__buf_1 _28179_ (.A(\reg_pc[26] ),
    .X(_21816_));
 sky130_fd_sc_hd__buf_1 _28180_ (.A(_21816_),
    .X(_21817_));
 sky130_fd_sc_hd__nand3_4 _28181_ (.A(_21787_),
    .B(_21815_),
    .C(_21817_),
    .Y(_21818_));
 sky130_fd_sc_hd__buf_1 _28182_ (.A(_21115_),
    .X(_21819_));
 sky130_fd_sc_hd__a21o_4 _28183_ (.A1(_21814_),
    .A2(_21818_),
    .B1(_21819_),
    .X(_21820_));
 sky130_fd_sc_hd__a21o_4 _28184_ (.A1(_21813_),
    .A2(_21820_),
    .B1(_21791_),
    .X(_21821_));
 sky130_fd_sc_hd__o21ai_4 _28185_ (.A1(_21804_),
    .A2(_21794_),
    .B1(_21821_),
    .Y(_00548_));
 sky130_fd_sc_hd__buf_1 _28186_ (.A(_18758_),
    .X(_21822_));
 sky130_fd_sc_hd__xor2_4 _28187_ (.A(pcpi_rs1[27]),
    .B(\decoded_imm[27] ),
    .X(_21823_));
 sky130_vsdinv _28188_ (.A(_21823_),
    .Y(_21824_));
 sky130_fd_sc_hd__maj3_4 _28189_ (.A(_21804_),
    .B(_21811_),
    .C(_21319_),
    .X(_21825_));
 sky130_fd_sc_hd__nor2_4 _28190_ (.A(_21824_),
    .B(_21825_),
    .Y(_21826_));
 sky130_fd_sc_hd__a21o_4 _28191_ (.A1(_21825_),
    .A2(_21824_),
    .B1(_21713_),
    .X(_21827_));
 sky130_fd_sc_hd__buf_1 _28192_ (.A(\reg_pc[27] ),
    .X(_21828_));
 sky130_fd_sc_hd__buf_1 _28193_ (.A(_21828_),
    .X(_21829_));
 sky130_fd_sc_hd__nand3_4 _28194_ (.A(_21585_),
    .B(_21416_),
    .C(_21829_),
    .Y(_21830_));
 sky130_fd_sc_hd__o21ai_4 _28195_ (.A1(_21584_),
    .A2(_20842_),
    .B1(_21830_),
    .Y(_21831_));
 sky130_fd_sc_hd__a2bb2o_4 _28196_ (.A1_N(_21826_),
    .A2_N(_21827_),
    .B1(_21184_),
    .B2(_21831_),
    .X(_21832_));
 sky130_fd_sc_hd__a2bb2o_4 _28197_ (.A1_N(_21822_),
    .A2_N(_21395_),
    .B1(_21708_),
    .B2(_21832_),
    .X(_00549_));
 sky130_fd_sc_hd__buf_1 _28198_ (.A(pcpi_rs1[28]),
    .X(_21833_));
 sky130_vsdinv _28199_ (.A(_21833_),
    .Y(_21834_));
 sky130_fd_sc_hd__nand2_4 _28200_ (.A(_18746_),
    .B(\decoded_imm[28] ),
    .Y(_21835_));
 sky130_fd_sc_hd__nor2_4 _28201_ (.A(_21833_),
    .B(\decoded_imm[28] ),
    .Y(_21836_));
 sky130_vsdinv _28202_ (.A(_21836_),
    .Y(_21837_));
 sky130_vsdinv _28203_ (.A(_21807_),
    .Y(_21838_));
 sky130_fd_sc_hd__a21oi_4 _28204_ (.A1(_21780_),
    .A2(_21782_),
    .B1(_21838_),
    .Y(_21839_));
 sky130_fd_sc_hd__and2_4 _28205_ (.A(_21805_),
    .B(_21823_),
    .X(_21840_));
 sky130_fd_sc_hd__o21ai_4 _28206_ (.A1(_21810_),
    .A2(_21839_),
    .B1(_21840_),
    .Y(_21841_));
 sky130_fd_sc_hd__nand2_4 _28207_ (.A(_18720_),
    .B(_21318_),
    .Y(_21842_));
 sky130_fd_sc_hd__maj3_4 _28208_ (.A(_18758_),
    .B(_21842_),
    .C(_21322_),
    .X(_21843_));
 sky130_fd_sc_hd__nand2_4 _28209_ (.A(_21841_),
    .B(_21843_),
    .Y(_21844_));
 sky130_fd_sc_hd__a21o_4 _28210_ (.A1(_21835_),
    .A2(_21837_),
    .B1(_21844_),
    .X(_21845_));
 sky130_fd_sc_hd__nand3_4 _28211_ (.A(_21844_),
    .B(_21835_),
    .C(_21837_),
    .Y(_21846_));
 sky130_fd_sc_hd__nand3_4 _28212_ (.A(_21845_),
    .B(_21597_),
    .C(_21846_),
    .Y(_21847_));
 sky130_fd_sc_hd__a2111o_4 _28213_ (.A1(_20859_),
    .A2(_20873_),
    .B1(_21733_),
    .C1(_19382_),
    .D1(_20882_),
    .X(_21848_));
 sky130_fd_sc_hd__buf_1 _28214_ (.A(\reg_pc[28] ),
    .X(_21849_));
 sky130_fd_sc_hd__buf_1 _28215_ (.A(_21849_),
    .X(_21850_));
 sky130_fd_sc_hd__nand3_4 _28216_ (.A(_21787_),
    .B(_21815_),
    .C(_21850_),
    .Y(_21851_));
 sky130_fd_sc_hd__a21o_4 _28217_ (.A1(_21848_),
    .A2(_21851_),
    .B1(_21819_),
    .X(_21852_));
 sky130_fd_sc_hd__a21o_4 _28218_ (.A1(_21847_),
    .A2(_21852_),
    .B1(_21791_),
    .X(_21853_));
 sky130_fd_sc_hd__o21ai_4 _28219_ (.A1(_21834_),
    .A2(_21794_),
    .B1(_21853_),
    .Y(_00550_));
 sky130_vsdinv _28220_ (.A(pcpi_rs1[29]),
    .Y(_21854_));
 sky130_fd_sc_hd__buf_1 _28221_ (.A(_18751_),
    .X(_21855_));
 sky130_fd_sc_hd__xor2_4 _28222_ (.A(_21855_),
    .B(_21330_),
    .X(_21856_));
 sky130_vsdinv _28223_ (.A(_21856_),
    .Y(_21857_));
 sky130_vsdinv _28224_ (.A(_21835_),
    .Y(_21858_));
 sky130_fd_sc_hd__a21oi_4 _28225_ (.A1(_21844_),
    .A2(_21837_),
    .B1(_21858_),
    .Y(_21859_));
 sky130_fd_sc_hd__o21ai_4 _28226_ (.A1(_21857_),
    .A2(_21859_),
    .B1(_21681_),
    .Y(_21860_));
 sky130_fd_sc_hd__a21o_4 _28227_ (.A1(_21857_),
    .A2(_21859_),
    .B1(_21860_),
    .X(_21861_));
 sky130_fd_sc_hd__a2111o_4 _28228_ (.A1(_20908_),
    .A2(_20922_),
    .B1(_21415_),
    .C1(_19382_),
    .D1(_20929_),
    .X(_21862_));
 sky130_fd_sc_hd__buf_1 _28229_ (.A(\reg_pc[29] ),
    .X(_21863_));
 sky130_fd_sc_hd__buf_1 _28230_ (.A(_21863_),
    .X(_21864_));
 sky130_fd_sc_hd__buf_1 _28231_ (.A(_21864_),
    .X(_21865_));
 sky130_fd_sc_hd__nand3_4 _28232_ (.A(_21787_),
    .B(_21815_),
    .C(_21865_),
    .Y(_21866_));
 sky130_fd_sc_hd__a21o_4 _28233_ (.A1(_21862_),
    .A2(_21866_),
    .B1(_21819_),
    .X(_21867_));
 sky130_fd_sc_hd__a21o_4 _28234_ (.A1(_21861_),
    .A2(_21867_),
    .B1(_21347_),
    .X(_21868_));
 sky130_fd_sc_hd__o21ai_4 _28235_ (.A1(_21854_),
    .A2(_21794_),
    .B1(_21868_),
    .Y(_00551_));
 sky130_fd_sc_hd__buf_1 _28236_ (.A(pcpi_rs1[30]),
    .X(_21869_));
 sky130_vsdinv _28237_ (.A(_21869_),
    .Y(_21870_));
 sky130_fd_sc_hd__buf_1 _28238_ (.A(_21869_),
    .X(_21871_));
 sky130_fd_sc_hd__nand2_4 _28239_ (.A(_21871_),
    .B(_21336_),
    .Y(_21872_));
 sky130_fd_sc_hd__nor2_4 _28240_ (.A(_21869_),
    .B(\decoded_imm[30] ),
    .Y(_21873_));
 sky130_vsdinv _28241_ (.A(_21873_),
    .Y(_21874_));
 sky130_fd_sc_hd__a21oi_4 _28242_ (.A1(_21841_),
    .A2(_21843_),
    .B1(_21836_),
    .Y(_21875_));
 sky130_fd_sc_hd__nor2_4 _28243_ (.A(_21855_),
    .B(\decoded_imm[29] ),
    .Y(_21876_));
 sky130_vsdinv _28244_ (.A(_21876_),
    .Y(_21877_));
 sky130_fd_sc_hd__o21ai_4 _28245_ (.A1(_21858_),
    .A2(_21875_),
    .B1(_21877_),
    .Y(_21878_));
 sky130_fd_sc_hd__buf_1 _28246_ (.A(_21855_),
    .X(_21879_));
 sky130_fd_sc_hd__nand2_4 _28247_ (.A(_21879_),
    .B(_21330_),
    .Y(_21880_));
 sky130_fd_sc_hd__nand2_4 _28248_ (.A(_21878_),
    .B(_21880_),
    .Y(_21881_));
 sky130_fd_sc_hd__a21o_4 _28249_ (.A1(_21872_),
    .A2(_21874_),
    .B1(_21881_),
    .X(_21882_));
 sky130_fd_sc_hd__nand3_4 _28250_ (.A(_21881_),
    .B(_21872_),
    .C(_21874_),
    .Y(_21883_));
 sky130_fd_sc_hd__nand3_4 _28251_ (.A(_21882_),
    .B(_21597_),
    .C(_21883_),
    .Y(_21884_));
 sky130_fd_sc_hd__a2111o_4 _28252_ (.A1(_20948_),
    .A2(_20962_),
    .B1(_21415_),
    .C1(_19382_),
    .D1(_20969_),
    .X(_21885_));
 sky130_fd_sc_hd__buf_1 _28253_ (.A(\reg_pc[30] ),
    .X(_21886_));
 sky130_fd_sc_hd__buf_1 _28254_ (.A(_21886_),
    .X(_21887_));
 sky130_fd_sc_hd__nand3_4 _28255_ (.A(_21359_),
    .B(_21815_),
    .C(_21887_),
    .Y(_21888_));
 sky130_fd_sc_hd__a21o_4 _28256_ (.A1(_21885_),
    .A2(_21888_),
    .B1(_21819_),
    .X(_21889_));
 sky130_fd_sc_hd__a21o_4 _28257_ (.A1(_21884_),
    .A2(_21889_),
    .B1(_21791_),
    .X(_21890_));
 sky130_fd_sc_hd__o21ai_4 _28258_ (.A1(_21870_),
    .A2(_21582_),
    .B1(_21890_),
    .Y(_00553_));
 sky130_vsdinv _28259_ (.A(_21872_),
    .Y(_21891_));
 sky130_fd_sc_hd__a21oi_4 _28260_ (.A1(_21878_),
    .A2(_21880_),
    .B1(_21873_),
    .Y(_21892_));
 sky130_fd_sc_hd__xor2_4 _28261_ (.A(_18741_),
    .B(\decoded_imm[31] ),
    .X(_21893_));
 sky130_fd_sc_hd__o21ai_4 _28262_ (.A1(_21891_),
    .A2(_21892_),
    .B1(_21893_),
    .Y(_21894_));
 sky130_fd_sc_hd__nand2_4 _28263_ (.A(_21881_),
    .B(_21874_),
    .Y(_21895_));
 sky130_vsdinv _28264_ (.A(_21893_),
    .Y(_21896_));
 sky130_fd_sc_hd__nand3_4 _28265_ (.A(_21895_),
    .B(_21872_),
    .C(_21896_),
    .Y(_21897_));
 sky130_fd_sc_hd__nand3_4 _28266_ (.A(_21894_),
    .B(_21682_),
    .C(_21897_),
    .Y(_21898_));
 sky130_fd_sc_hd__a2111o_4 _28267_ (.A1(_20991_),
    .A2(_21005_),
    .B1(_21410_),
    .C1(_21411_),
    .D1(_21012_),
    .X(_21899_));
 sky130_fd_sc_hd__buf_1 _28268_ (.A(\reg_pc[31] ),
    .X(_21900_));
 sky130_fd_sc_hd__nand3_4 _28269_ (.A(_21585_),
    .B(_21416_),
    .C(_21900_),
    .Y(_21901_));
 sky130_fd_sc_hd__a21o_4 _28270_ (.A1(_21899_),
    .A2(_21901_),
    .B1(_21460_),
    .X(_21902_));
 sky130_fd_sc_hd__nand2_4 _28271_ (.A(_21898_),
    .B(_21902_),
    .Y(_21903_));
 sky130_fd_sc_hd__nand2_4 _28272_ (.A(_21903_),
    .B(_21708_),
    .Y(_21904_));
 sky130_fd_sc_hd__buf_1 _28273_ (.A(_18741_),
    .X(_21905_));
 sky130_fd_sc_hd__buf_1 _28274_ (.A(_21905_),
    .X(_21906_));
 sky130_fd_sc_hd__nand2_4 _28275_ (.A(_21393_),
    .B(_21906_),
    .Y(_21907_));
 sky130_fd_sc_hd__nand2_4 _28276_ (.A(_21904_),
    .B(_21907_),
    .Y(_00554_));
 sky130_vsdinv _28277_ (.A(latched_branch),
    .Y(_21908_));
 sky130_vsdinv _28278_ (.A(\reg_next_pc[0] ),
    .Y(_21909_));
 sky130_fd_sc_hd__nand2_4 _28279_ (.A(latched_branch),
    .B(latched_store),
    .Y(_21910_));
 sky130_vsdinv _28280_ (.A(_21910_),
    .Y(_21911_));
 sky130_fd_sc_hd__buf_1 _28281_ (.A(_21911_),
    .X(_21912_));
 sky130_fd_sc_hd__buf_1 _28282_ (.A(_21912_),
    .X(_21913_));
 sky130_fd_sc_hd__buf_1 _28283_ (.A(_21913_),
    .X(_21914_));
 sky130_fd_sc_hd__buf_1 _28284_ (.A(_21914_),
    .X(_21915_));
 sky130_fd_sc_hd__buf_1 _28285_ (.A(_21915_),
    .X(_21916_));
 sky130_fd_sc_hd__buf_1 _28286_ (.A(_21916_),
    .X(_21917_));
 sky130_fd_sc_hd__buf_1 _28287_ (.A(_21917_),
    .X(_21918_));
 sky130_fd_sc_hd__buf_1 _28288_ (.A(_21918_),
    .X(_21919_));
 sky130_fd_sc_hd__a211o_4 _28289_ (.A1(_19077_),
    .A2(_21908_),
    .B1(_21909_),
    .C1(_21919_),
    .X(_21920_));
 sky130_vsdinv _28290_ (.A(_18539_),
    .Y(_21921_));
 sky130_fd_sc_hd__buf_1 _28291_ (.A(_21921_),
    .X(_21922_));
 sky130_fd_sc_hd__buf_1 _28292_ (.A(_21922_),
    .X(_21923_));
 sky130_fd_sc_hd__buf_1 _28293_ (.A(\decoded_imm_uj[0] ),
    .X(_21924_));
 sky130_vsdinv _28294_ (.A(_21924_),
    .Y(_21925_));
 sky130_fd_sc_hd__buf_1 _28295_ (.A(_19136_),
    .X(_21926_));
 sky130_fd_sc_hd__buf_1 _28296_ (.A(_18566_),
    .X(_21927_));
 sky130_fd_sc_hd__buf_1 _28297_ (.A(_18544_),
    .X(_21928_));
 sky130_fd_sc_hd__nand3_4 _28298_ (.A(_18778_),
    .B(_21927_),
    .C(_21928_),
    .Y(_21929_));
 sky130_fd_sc_hd__nor4_4 _28299_ (.A(_21923_),
    .B(_21925_),
    .C(_21926_),
    .D(_21929_),
    .Y(_21930_));
 sky130_fd_sc_hd__o21a_4 _28300_ (.A1(_21920_),
    .A2(_21930_),
    .B1(_19102_),
    .X(_21931_));
 sky130_fd_sc_hd__nand4_4 _28301_ (.A(_18777_),
    .B(_18781_),
    .C(_21924_),
    .D(_21920_),
    .Y(_21932_));
 sky130_fd_sc_hd__buf_1 _28302_ (.A(_19125_),
    .X(_21933_));
 sky130_fd_sc_hd__o21ai_4 _28303_ (.A1(_19116_),
    .A2(\reg_next_pc[0] ),
    .B1(_21933_),
    .Y(_21934_));
 sky130_fd_sc_hd__a21oi_4 _28304_ (.A1(_21931_),
    .A2(_21932_),
    .B1(_21934_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_4 _28305_ (.A(_21908_),
    .B(\irq_state[0] ),
    .Y(_21935_));
 sky130_fd_sc_hd__and4_4 _28306_ (.A(_21935_),
    .B(\reg_next_pc[0] ),
    .C(\decoded_imm_uj[0] ),
    .D(_21910_),
    .X(_21936_));
 sky130_fd_sc_hd__buf_1 _28307_ (.A(_21910_),
    .X(_21937_));
 sky130_vsdinv _28308_ (.A(latched_stalu),
    .Y(_21938_));
 sky130_fd_sc_hd__buf_1 _28309_ (.A(_21938_),
    .X(_21939_));
 sky130_fd_sc_hd__or2_4 _28310_ (.A(\reg_out[1] ),
    .B(latched_stalu),
    .X(_21940_));
 sky130_fd_sc_hd__o21ai_4 _28311_ (.A1(\alu_out_q[1] ),
    .A2(_21939_),
    .B1(_21940_),
    .Y(_21941_));
 sky130_fd_sc_hd__nand3_4 _28312_ (.A(_21935_),
    .B(\reg_next_pc[1] ),
    .C(_21910_),
    .Y(_21942_));
 sky130_fd_sc_hd__o21ai_4 _28313_ (.A1(_21937_),
    .A2(_21941_),
    .B1(_21942_),
    .Y(_21943_));
 sky130_fd_sc_hd__xor2_4 _28314_ (.A(\decoded_imm_uj[1] ),
    .B(_21943_),
    .X(_21944_));
 sky130_fd_sc_hd__or2_4 _28315_ (.A(_21936_),
    .B(_21944_),
    .X(_21945_));
 sky130_fd_sc_hd__nand2_4 _28316_ (.A(_21944_),
    .B(_21936_),
    .Y(_21946_));
 sky130_fd_sc_hd__a41oi_4 _28317_ (.A1(_18777_),
    .A2(_18780_),
    .A3(_21945_),
    .A4(_21946_),
    .B1(_18579_),
    .Y(_21947_));
 sky130_fd_sc_hd__buf_1 _28318_ (.A(_18484_),
    .X(_21948_));
 sky130_fd_sc_hd__buf_1 _28319_ (.A(_18540_),
    .X(_21949_));
 sky130_fd_sc_hd__buf_1 _28320_ (.A(_21949_),
    .X(_21950_));
 sky130_fd_sc_hd__buf_1 _28321_ (.A(_18542_),
    .X(_21951_));
 sky130_fd_sc_hd__buf_1 _28322_ (.A(_21951_),
    .X(_21952_));
 sky130_fd_sc_hd__buf_1 _28323_ (.A(_18557_),
    .X(_21953_));
 sky130_fd_sc_hd__buf_1 _28324_ (.A(_21953_),
    .X(_21954_));
 sky130_vsdinv _28325_ (.A(_21943_),
    .Y(_21955_));
 sky130_fd_sc_hd__a41o_4 _28326_ (.A1(_21948_),
    .A2(_21950_),
    .A3(_21952_),
    .A4(_21954_),
    .B1(_21955_),
    .X(_21956_));
 sky130_fd_sc_hd__o21ai_4 _28327_ (.A1(_19116_),
    .A2(\reg_next_pc[1] ),
    .B1(_21933_),
    .Y(_21957_));
 sky130_fd_sc_hd__a21oi_4 _28328_ (.A1(_21947_),
    .A2(_21956_),
    .B1(_21957_),
    .Y(_00509_));
 sky130_fd_sc_hd__buf_1 _28329_ (.A(_19134_),
    .X(_21958_));
 sky130_fd_sc_hd__buf_1 _28330_ (.A(_21958_),
    .X(_21959_));
 sky130_fd_sc_hd__buf_1 _28331_ (.A(latched_branch),
    .X(_21960_));
 sky130_fd_sc_hd__nor2_4 _28332_ (.A(\irq_state[0] ),
    .B(_21960_),
    .Y(_21961_));
 sky130_vsdinv _28333_ (.A(latched_store),
    .Y(_21962_));
 sky130_fd_sc_hd__or2_4 _28334_ (.A(latched_stalu),
    .B(\reg_out[2] ),
    .X(_21963_));
 sky130_fd_sc_hd__o21a_4 _28335_ (.A1(_21939_),
    .A2(\alu_out_q[2] ),
    .B1(_21963_),
    .X(_21964_));
 sky130_fd_sc_hd__o21a_4 _28336_ (.A1(_21962_),
    .A2(_21964_),
    .B1(_21960_),
    .X(_21965_));
 sky130_fd_sc_hd__o21ai_4 _28337_ (.A1(_21961_),
    .A2(_21965_),
    .B1(\reg_next_pc[2] ),
    .Y(_21966_));
 sky130_fd_sc_hd__buf_1 _28338_ (.A(_21960_),
    .X(_21967_));
 sky130_fd_sc_hd__buf_1 _28339_ (.A(latched_store),
    .X(_21968_));
 sky130_fd_sc_hd__nand3_4 _28340_ (.A(_21964_),
    .B(_21967_),
    .C(_21968_),
    .Y(_21969_));
 sky130_fd_sc_hd__nand2_4 _28341_ (.A(_21966_),
    .B(_21969_),
    .Y(_21970_));
 sky130_fd_sc_hd__buf_1 _28342_ (.A(_21970_),
    .X(_21971_));
 sky130_fd_sc_hd__buf_1 _28343_ (.A(_21971_),
    .X(_21972_));
 sky130_fd_sc_hd__buf_1 _28344_ (.A(_18404_),
    .X(_21973_));
 sky130_fd_sc_hd__buf_1 _28345_ (.A(_21973_),
    .X(_21974_));
 sky130_fd_sc_hd__buf_1 _28346_ (.A(_21974_),
    .X(_21975_));
 sky130_vsdinv _28347_ (.A(\decoded_imm_uj[2] ),
    .Y(_21976_));
 sky130_fd_sc_hd__a21oi_4 _28348_ (.A1(_21966_),
    .A2(_21969_),
    .B1(_21976_),
    .Y(_21977_));
 sky130_vsdinv _28349_ (.A(_21977_),
    .Y(_21978_));
 sky130_fd_sc_hd__nand3_4 _28350_ (.A(_21966_),
    .B(_21976_),
    .C(_21969_),
    .Y(_21979_));
 sky130_fd_sc_hd__maj3_4 _28351_ (.A(\decoded_imm_uj[1] ),
    .B(_21943_),
    .C(_21936_),
    .X(_21980_));
 sky130_vsdinv _28352_ (.A(_21980_),
    .Y(_21981_));
 sky130_fd_sc_hd__a21o_4 _28353_ (.A1(_21978_),
    .A2(_21979_),
    .B1(_21981_),
    .X(_21982_));
 sky130_fd_sc_hd__nand3_4 _28354_ (.A(_21978_),
    .B(_21979_),
    .C(_21981_),
    .Y(_21983_));
 sky130_fd_sc_hd__nand3_4 _28355_ (.A(_21982_),
    .B(_18540_),
    .C(_21983_),
    .Y(_21984_));
 sky130_fd_sc_hd__buf_1 _28356_ (.A(_18566_),
    .X(_21985_));
 sky130_fd_sc_hd__buf_1 _28357_ (.A(_21921_),
    .X(_21986_));
 sky130_fd_sc_hd__nand2_4 _28358_ (.A(_21971_),
    .B(_21986_),
    .Y(_21987_));
 sky130_fd_sc_hd__and3_4 _28359_ (.A(_21984_),
    .B(_21985_),
    .C(_21987_),
    .X(_21988_));
 sky130_fd_sc_hd__a211o_4 _28360_ (.A1(_21959_),
    .A2(_21972_),
    .B1(_21975_),
    .C1(_21988_),
    .X(_21989_));
 sky130_fd_sc_hd__buf_1 _28361_ (.A(_18485_),
    .X(_21990_));
 sky130_fd_sc_hd__buf_1 _28362_ (.A(\irq_pending[2] ),
    .X(_21991_));
 sky130_fd_sc_hd__or2_4 _28363_ (.A(_21991_),
    .B(_18946_),
    .X(_21992_));
 sky130_vsdinv _28364_ (.A(\irq_pending[4] ),
    .Y(_21993_));
 sky130_vsdinv _28365_ (.A(\irq_pending[5] ),
    .Y(_21994_));
 sky130_vsdinv _28366_ (.A(\irq_pending[6] ),
    .Y(_21995_));
 sky130_vsdinv _28367_ (.A(\irq_pending[7] ),
    .Y(_21996_));
 sky130_fd_sc_hd__nand4_4 _28368_ (.A(_21993_),
    .B(_21994_),
    .C(_21995_),
    .D(_21996_),
    .Y(_21997_));
 sky130_fd_sc_hd__nor4_4 _28369_ (.A(_18907_),
    .B(\irq_pending[1] ),
    .C(_21992_),
    .D(_21997_),
    .Y(_21998_));
 sky130_vsdinv _28370_ (.A(\irq_pending[20] ),
    .Y(_21999_));
 sky130_vsdinv _28371_ (.A(\irq_pending[21] ),
    .Y(_22000_));
 sky130_vsdinv _28372_ (.A(\irq_pending[22] ),
    .Y(_22001_));
 sky130_vsdinv _28373_ (.A(\irq_pending[23] ),
    .Y(_22002_));
 sky130_fd_sc_hd__nand4_4 _28374_ (.A(_21999_),
    .B(_22000_),
    .C(_22001_),
    .D(_22002_),
    .Y(_22003_));
 sky130_vsdinv _28375_ (.A(\irq_pending[16] ),
    .Y(_22004_));
 sky130_vsdinv _28376_ (.A(\irq_pending[17] ),
    .Y(_22005_));
 sky130_vsdinv _28377_ (.A(\irq_pending[18] ),
    .Y(_22006_));
 sky130_vsdinv _28378_ (.A(\irq_pending[19] ),
    .Y(_22007_));
 sky130_fd_sc_hd__nand4_4 _28379_ (.A(_22004_),
    .B(_22005_),
    .C(_22006_),
    .D(_22007_),
    .Y(_22008_));
 sky130_fd_sc_hd__nor2_4 _28380_ (.A(_22003_),
    .B(_22008_),
    .Y(_22009_));
 sky130_vsdinv _28381_ (.A(\irq_pending[28] ),
    .Y(_22010_));
 sky130_vsdinv _28382_ (.A(\irq_pending[29] ),
    .Y(_22011_));
 sky130_vsdinv _28383_ (.A(\irq_pending[30] ),
    .Y(_22012_));
 sky130_vsdinv _28384_ (.A(\irq_pending[31] ),
    .Y(_22013_));
 sky130_fd_sc_hd__nand4_4 _28385_ (.A(_22010_),
    .B(_22011_),
    .C(_22012_),
    .D(_22013_),
    .Y(_22014_));
 sky130_vsdinv _28386_ (.A(\irq_pending[24] ),
    .Y(_22015_));
 sky130_vsdinv _28387_ (.A(\irq_pending[25] ),
    .Y(_22016_));
 sky130_vsdinv _28388_ (.A(\irq_pending[26] ),
    .Y(_22017_));
 sky130_vsdinv _28389_ (.A(\irq_pending[27] ),
    .Y(_22018_));
 sky130_fd_sc_hd__nand4_4 _28390_ (.A(_22015_),
    .B(_22016_),
    .C(_22017_),
    .D(_22018_),
    .Y(_22019_));
 sky130_fd_sc_hd__nor2_4 _28391_ (.A(_22014_),
    .B(_22019_),
    .Y(_22020_));
 sky130_vsdinv _28392_ (.A(\irq_pending[12] ),
    .Y(_22021_));
 sky130_vsdinv _28393_ (.A(\irq_pending[13] ),
    .Y(_22022_));
 sky130_vsdinv _28394_ (.A(\irq_pending[14] ),
    .Y(_22023_));
 sky130_vsdinv _28395_ (.A(\irq_pending[15] ),
    .Y(_22024_));
 sky130_fd_sc_hd__nand4_4 _28396_ (.A(_22021_),
    .B(_22022_),
    .C(_22023_),
    .D(_22024_),
    .Y(_22025_));
 sky130_vsdinv _28397_ (.A(\irq_pending[8] ),
    .Y(_22026_));
 sky130_vsdinv _28398_ (.A(\irq_pending[9] ),
    .Y(_22027_));
 sky130_vsdinv _28399_ (.A(\irq_pending[10] ),
    .Y(_22028_));
 sky130_vsdinv _28400_ (.A(\irq_pending[11] ),
    .Y(_22029_));
 sky130_fd_sc_hd__nand4_4 _28401_ (.A(_22026_),
    .B(_22027_),
    .C(_22028_),
    .D(_22029_),
    .Y(_22030_));
 sky130_fd_sc_hd__nor2_4 _28402_ (.A(_22025_),
    .B(_22030_),
    .Y(_22031_));
 sky130_fd_sc_hd__and4_4 _28403_ (.A(_21998_),
    .B(_22009_),
    .C(_22020_),
    .D(_22031_),
    .X(_22032_));
 sky130_fd_sc_hd__buf_1 _28404_ (.A(_22032_),
    .X(_22033_));
 sky130_fd_sc_hd__buf_1 _28405_ (.A(_22033_),
    .X(_22034_));
 sky130_fd_sc_hd__buf_1 _28406_ (.A(_18553_),
    .X(_22035_));
 sky130_fd_sc_hd__a21oi_4 _28407_ (.A1(_21971_),
    .A2(_22034_),
    .B1(_22035_),
    .Y(_22036_));
 sky130_fd_sc_hd__o21ai_4 _28408_ (.A1(_21972_),
    .A2(_22034_),
    .B1(_22036_),
    .Y(_22037_));
 sky130_fd_sc_hd__nand3_4 _28409_ (.A(_21989_),
    .B(_21990_),
    .C(_22037_),
    .Y(_22038_));
 sky130_fd_sc_hd__buf_1 _28410_ (.A(_18547_),
    .X(_22039_));
 sky130_fd_sc_hd__a21oi_4 _28411_ (.A1(_22039_),
    .A2(_21972_),
    .B1(_19092_),
    .Y(_22040_));
 sky130_fd_sc_hd__buf_1 _28412_ (.A(_19115_),
    .X(_22041_));
 sky130_fd_sc_hd__o21ai_4 _28413_ (.A1(_22041_),
    .A2(\reg_next_pc[2] ),
    .B1(_21933_),
    .Y(_22042_));
 sky130_fd_sc_hd__a21oi_4 _28414_ (.A1(_22038_),
    .A2(_22040_),
    .B1(_22042_),
    .Y(_00520_));
 sky130_fd_sc_hd__buf_1 _28415_ (.A(_21938_),
    .X(_22043_));
 sky130_fd_sc_hd__buf_1 _28416_ (.A(latched_stalu),
    .X(_22044_));
 sky130_fd_sc_hd__or2_4 _28417_ (.A(_22044_),
    .B(\reg_out[3] ),
    .X(_22045_));
 sky130_fd_sc_hd__o21a_4 _28418_ (.A1(_22043_),
    .A2(\alu_out_q[3] ),
    .B1(_22045_),
    .X(_22046_));
 sky130_fd_sc_hd__nand2_4 _28419_ (.A(_22046_),
    .B(_21911_),
    .Y(_22047_));
 sky130_fd_sc_hd__buf_1 _28420_ (.A(_21935_),
    .X(_22048_));
 sky130_fd_sc_hd__buf_1 _28421_ (.A(_21937_),
    .X(_22049_));
 sky130_fd_sc_hd__nand3_4 _28422_ (.A(_22048_),
    .B(\reg_next_pc[3] ),
    .C(_22049_),
    .Y(_22050_));
 sky130_vsdinv _28423_ (.A(\decoded_imm_uj[3] ),
    .Y(_22051_));
 sky130_fd_sc_hd__a21oi_4 _28424_ (.A1(_22047_),
    .A2(_22050_),
    .B1(_22051_),
    .Y(_22052_));
 sky130_fd_sc_hd__nand3_4 _28425_ (.A(_22047_),
    .B(_22051_),
    .C(_22050_),
    .Y(_22053_));
 sky130_vsdinv _28426_ (.A(_22053_),
    .Y(_22054_));
 sky130_fd_sc_hd__nor2_4 _28427_ (.A(_22052_),
    .B(_22054_),
    .Y(_22055_));
 sky130_fd_sc_hd__a21oi_4 _28428_ (.A1(_21979_),
    .A2(_21980_),
    .B1(_21977_),
    .Y(_22056_));
 sky130_fd_sc_hd__buf_1 _28429_ (.A(_18774_),
    .X(_22057_));
 sky130_fd_sc_hd__o21ai_4 _28430_ (.A1(_22055_),
    .A2(_22056_),
    .B1(_22057_),
    .Y(_22058_));
 sky130_fd_sc_hd__a21o_4 _28431_ (.A1(_22055_),
    .A2(_22056_),
    .B1(_22058_),
    .X(_22059_));
 sky130_fd_sc_hd__nand2_4 _28432_ (.A(_22047_),
    .B(_22050_),
    .Y(_22060_));
 sky130_fd_sc_hd__buf_1 _28433_ (.A(_22060_),
    .X(_22061_));
 sky130_vsdinv _28434_ (.A(_22061_),
    .Y(_22062_));
 sky130_fd_sc_hd__xor2_4 _28435_ (.A(_22062_),
    .B(_21971_),
    .X(_22063_));
 sky130_fd_sc_hd__buf_1 _28436_ (.A(_21986_),
    .X(_22064_));
 sky130_fd_sc_hd__nor2_4 _28437_ (.A(_18342_),
    .B(_19133_),
    .Y(_22065_));
 sky130_vsdinv _28438_ (.A(_22065_),
    .Y(_22066_));
 sky130_fd_sc_hd__buf_1 _28439_ (.A(_22066_),
    .X(_22067_));
 sky130_fd_sc_hd__a21oi_4 _28440_ (.A1(_22063_),
    .A2(_22064_),
    .B1(_22067_),
    .Y(_22068_));
 sky130_fd_sc_hd__nand2_4 _28441_ (.A(_22059_),
    .B(_22068_),
    .Y(_22069_));
 sky130_vsdinv _28442_ (.A(_22032_),
    .Y(_22070_));
 sky130_fd_sc_hd__buf_1 _28443_ (.A(_22070_),
    .X(_22071_));
 sky130_fd_sc_hd__buf_1 _28444_ (.A(_18407_),
    .X(_22072_));
 sky130_fd_sc_hd__and2_4 _28445_ (.A(_21998_),
    .B(_22031_),
    .X(_22073_));
 sky130_fd_sc_hd__buf_1 _28446_ (.A(_22073_),
    .X(_22074_));
 sky130_fd_sc_hd__buf_1 _28447_ (.A(_22074_),
    .X(_22075_));
 sky130_fd_sc_hd__and2_4 _28448_ (.A(_22009_),
    .B(_22020_),
    .X(_22076_));
 sky130_fd_sc_hd__buf_1 _28449_ (.A(_22076_),
    .X(_22077_));
 sky130_fd_sc_hd__buf_1 _28450_ (.A(_22077_),
    .X(_22078_));
 sky130_fd_sc_hd__nand3_4 _28451_ (.A(_22075_),
    .B(_22078_),
    .C(_22062_),
    .Y(_22079_));
 sky130_vsdinv _28452_ (.A(_22079_),
    .Y(_22080_));
 sky130_fd_sc_hd__a211o_4 _28453_ (.A1(_22063_),
    .A2(_22071_),
    .B1(_22072_),
    .C1(_22080_),
    .X(_22081_));
 sky130_fd_sc_hd__a21o_4 _28454_ (.A1(_22069_),
    .A2(_22081_),
    .B1(_22039_),
    .X(_22082_));
 sky130_fd_sc_hd__o21ai_4 _28455_ (.A1(_18542_),
    .A2(_21973_),
    .B1(_18483_),
    .Y(_22083_));
 sky130_fd_sc_hd__buf_1 _28456_ (.A(_22083_),
    .X(_22084_));
 sky130_fd_sc_hd__buf_1 _28457_ (.A(_22084_),
    .X(_22085_));
 sky130_fd_sc_hd__a21oi_4 _28458_ (.A1(_22085_),
    .A2(_22061_),
    .B1(_19092_),
    .Y(_22086_));
 sky130_fd_sc_hd__o21ai_4 _28459_ (.A1(_22041_),
    .A2(\reg_next_pc[3] ),
    .B1(_21933_),
    .Y(_22087_));
 sky130_fd_sc_hd__a21oi_4 _28460_ (.A1(_22082_),
    .A2(_22086_),
    .B1(_22087_),
    .Y(_00523_));
 sky130_fd_sc_hd__or2_4 _28461_ (.A(_22044_),
    .B(\reg_out[4] ),
    .X(_22088_));
 sky130_fd_sc_hd__o21a_4 _28462_ (.A1(_22043_),
    .A2(\alu_out_q[4] ),
    .B1(_22088_),
    .X(_22089_));
 sky130_fd_sc_hd__a21o_4 _28463_ (.A1(_21960_),
    .A2(_21968_),
    .B1(\reg_next_pc[4] ),
    .X(_22090_));
 sky130_fd_sc_hd__o21ai_4 _28464_ (.A1(_21937_),
    .A2(_22089_),
    .B1(_22090_),
    .Y(_22091_));
 sky130_vsdinv _28465_ (.A(\irq_state[0] ),
    .Y(_22092_));
 sky130_fd_sc_hd__buf_1 _28466_ (.A(_22092_),
    .X(_22093_));
 sky130_fd_sc_hd__and2_4 _28467_ (.A(_22091_),
    .B(_22093_),
    .X(_22094_));
 sky130_fd_sc_hd__buf_1 _28468_ (.A(_22094_),
    .X(_22095_));
 sky130_vsdinv _28469_ (.A(_22095_),
    .Y(_22096_));
 sky130_fd_sc_hd__a21oi_4 _28470_ (.A1(_21970_),
    .A2(_22061_),
    .B1(_22096_),
    .Y(_22097_));
 sky130_fd_sc_hd__and3_4 _28471_ (.A(_21970_),
    .B(_22060_),
    .C(_22096_),
    .X(_22098_));
 sky130_fd_sc_hd__or2_4 _28472_ (.A(_22097_),
    .B(_22098_),
    .X(_22099_));
 sky130_fd_sc_hd__buf_1 _28473_ (.A(_22070_),
    .X(_22100_));
 sky130_fd_sc_hd__buf_1 _28474_ (.A(_22100_),
    .X(_22101_));
 sky130_fd_sc_hd__buf_1 _28475_ (.A(_18562_),
    .X(_22102_));
 sky130_fd_sc_hd__buf_1 _28476_ (.A(_22102_),
    .X(_22103_));
 sky130_fd_sc_hd__nor2_4 _28477_ (.A(_18541_),
    .B(do_waitirq),
    .Y(_22104_));
 sky130_fd_sc_hd__buf_1 _28478_ (.A(_22104_),
    .X(_22105_));
 sky130_fd_sc_hd__buf_1 _28479_ (.A(_22105_),
    .X(_22106_));
 sky130_fd_sc_hd__buf_1 _28480_ (.A(_22033_),
    .X(_22107_));
 sky130_fd_sc_hd__and2_4 _28481_ (.A(_22107_),
    .B(_22095_),
    .X(_22108_));
 sky130_fd_sc_hd__a2111oi_4 _28482_ (.A1(_22099_),
    .A2(_22101_),
    .B1(_22103_),
    .C1(_22106_),
    .D1(_22108_),
    .Y(_22109_));
 sky130_fd_sc_hd__buf_1 _28483_ (.A(_21921_),
    .X(_22110_));
 sky130_fd_sc_hd__buf_1 _28484_ (.A(_22110_),
    .X(_22111_));
 sky130_fd_sc_hd__buf_1 _28485_ (.A(_22111_),
    .X(_22112_));
 sky130_fd_sc_hd__buf_1 _28486_ (.A(_21974_),
    .X(_22113_));
 sky130_vsdinv _28487_ (.A(\decoded_imm_uj[4] ),
    .Y(_22114_));
 sky130_fd_sc_hd__a21o_4 _28488_ (.A1(_22091_),
    .A2(_22092_),
    .B1(_22114_),
    .X(_22115_));
 sky130_fd_sc_hd__buf_1 _28489_ (.A(_22115_),
    .X(_22116_));
 sky130_fd_sc_hd__nand3_4 _28490_ (.A(_22091_),
    .B(_22093_),
    .C(_22114_),
    .Y(_22117_));
 sky130_fd_sc_hd__and2_4 _28491_ (.A(_22116_),
    .B(_22117_),
    .X(_22118_));
 sky130_fd_sc_hd__nor2_4 _28492_ (.A(_22054_),
    .B(_22056_),
    .Y(_22119_));
 sky130_fd_sc_hd__a211o_4 _28493_ (.A1(\decoded_imm_uj[3] ),
    .A2(_22061_),
    .B1(_22118_),
    .C1(_22119_),
    .X(_22120_));
 sky130_fd_sc_hd__o21ai_4 _28494_ (.A1(_22052_),
    .A2(_22119_),
    .B1(_22118_),
    .Y(_22121_));
 sky130_fd_sc_hd__buf_1 _28495_ (.A(_21922_),
    .X(_22122_));
 sky130_fd_sc_hd__a21oi_4 _28496_ (.A1(_22120_),
    .A2(_22121_),
    .B1(_22122_),
    .Y(_22123_));
 sky130_fd_sc_hd__a2111oi_4 _28497_ (.A1(_22112_),
    .A2(_22099_),
    .B1(_21959_),
    .C1(_22113_),
    .D1(_22123_),
    .Y(_22124_));
 sky130_fd_sc_hd__buf_1 _28498_ (.A(_18485_),
    .X(_22125_));
 sky130_fd_sc_hd__o21ai_4 _28499_ (.A1(_22109_),
    .A2(_22124_),
    .B1(_22125_),
    .Y(_22126_));
 sky130_fd_sc_hd__buf_1 _28500_ (.A(_18551_),
    .X(_22127_));
 sky130_fd_sc_hd__a21oi_4 _28501_ (.A1(_22085_),
    .A2(_22096_),
    .B1(_22127_),
    .Y(_22128_));
 sky130_fd_sc_hd__buf_1 _28502_ (.A(_19125_),
    .X(_22129_));
 sky130_fd_sc_hd__o21ai_4 _28503_ (.A1(_22041_),
    .A2(\reg_next_pc[4] ),
    .B1(_22129_),
    .Y(_22130_));
 sky130_fd_sc_hd__a21oi_4 _28504_ (.A1(_22126_),
    .A2(_22128_),
    .B1(_22130_),
    .Y(_00524_));
 sky130_fd_sc_hd__buf_1 _28505_ (.A(_22044_),
    .X(_22131_));
 sky130_fd_sc_hd__or2_4 _28506_ (.A(\alu_out_q[5] ),
    .B(_21939_),
    .X(_22132_));
 sky130_fd_sc_hd__o21a_4 _28507_ (.A1(_22131_),
    .A2(\reg_out[5] ),
    .B1(_22132_),
    .X(_22133_));
 sky130_fd_sc_hd__nand2_4 _28508_ (.A(_22133_),
    .B(_21911_),
    .Y(_22134_));
 sky130_fd_sc_hd__nand3_4 _28509_ (.A(_22048_),
    .B(\reg_next_pc[5] ),
    .C(_21937_),
    .Y(_22135_));
 sky130_fd_sc_hd__nand2_4 _28510_ (.A(_22134_),
    .B(_22135_),
    .Y(_22136_));
 sky130_fd_sc_hd__nand2_4 _28511_ (.A(_22136_),
    .B(\decoded_imm_uj[5] ),
    .Y(_22137_));
 sky130_vsdinv _28512_ (.A(\decoded_imm_uj[5] ),
    .Y(_22138_));
 sky130_fd_sc_hd__nand3_4 _28513_ (.A(_22134_),
    .B(_22138_),
    .C(_22135_),
    .Y(_22139_));
 sky130_fd_sc_hd__a22oi_4 _28514_ (.A1(_22137_),
    .A2(_22139_),
    .B1(_22121_),
    .B2(_22116_),
    .Y(_22140_));
 sky130_fd_sc_hd__a41o_4 _28515_ (.A1(_22121_),
    .A2(_22116_),
    .A3(_22137_),
    .A4(_22139_),
    .B1(_22111_),
    .X(_22141_));
 sky130_vsdinv _28516_ (.A(_22136_),
    .Y(_22142_));
 sky130_fd_sc_hd__xor2_4 _28517_ (.A(_22142_),
    .B(_22098_),
    .X(_22143_));
 sky130_fd_sc_hd__buf_1 _28518_ (.A(_21986_),
    .X(_22144_));
 sky130_fd_sc_hd__buf_1 _28519_ (.A(_22066_),
    .X(_22145_));
 sky130_fd_sc_hd__a21oi_4 _28520_ (.A1(_22143_),
    .A2(_22144_),
    .B1(_22145_),
    .Y(_22146_));
 sky130_fd_sc_hd__o21ai_4 _28521_ (.A1(_22140_),
    .A2(_22141_),
    .B1(_22146_),
    .Y(_22147_));
 sky130_fd_sc_hd__buf_1 _28522_ (.A(_22074_),
    .X(_22148_));
 sky130_fd_sc_hd__buf_1 _28523_ (.A(_22077_),
    .X(_22149_));
 sky130_fd_sc_hd__nand3_4 _28524_ (.A(_22142_),
    .B(_22148_),
    .C(_22149_),
    .Y(_22150_));
 sky130_vsdinv _28525_ (.A(_22150_),
    .Y(_22151_));
 sky130_fd_sc_hd__a211o_4 _28526_ (.A1(_22143_),
    .A2(_22071_),
    .B1(_22072_),
    .C1(_22151_),
    .X(_22152_));
 sky130_fd_sc_hd__a21o_4 _28527_ (.A1(_22147_),
    .A2(_22152_),
    .B1(_22039_),
    .X(_22153_));
 sky130_fd_sc_hd__a21oi_4 _28528_ (.A1(_22085_),
    .A2(_22136_),
    .B1(_22127_),
    .Y(_22154_));
 sky130_fd_sc_hd__o21ai_4 _28529_ (.A1(_22041_),
    .A2(\reg_next_pc[5] ),
    .B1(_22129_),
    .Y(_22155_));
 sky130_fd_sc_hd__a21oi_4 _28530_ (.A1(_22153_),
    .A2(_22154_),
    .B1(_22155_),
    .Y(_00525_));
 sky130_fd_sc_hd__or2_4 _28531_ (.A(\alu_out_q[6] ),
    .B(_21939_),
    .X(_22156_));
 sky130_fd_sc_hd__o21a_4 _28532_ (.A1(_22131_),
    .A2(\reg_out[6] ),
    .B1(_22156_),
    .X(_22157_));
 sky130_fd_sc_hd__nand2_4 _28533_ (.A(_22157_),
    .B(_21911_),
    .Y(_22158_));
 sky130_fd_sc_hd__nand3_4 _28534_ (.A(_22048_),
    .B(\reg_next_pc[6] ),
    .C(_22049_),
    .Y(_22159_));
 sky130_fd_sc_hd__nand2_4 _28535_ (.A(_22158_),
    .B(_22159_),
    .Y(_22160_));
 sky130_fd_sc_hd__nand4_4 _28536_ (.A(_21970_),
    .B(_22060_),
    .C(_22096_),
    .D(_22136_),
    .Y(_22161_));
 sky130_fd_sc_hd__xor2_4 _28537_ (.A(_22160_),
    .B(_22161_),
    .X(_22162_));
 sky130_vsdinv _28538_ (.A(_22160_),
    .Y(_22163_));
 sky130_fd_sc_hd__buf_1 _28539_ (.A(_22163_),
    .X(_22164_));
 sky130_fd_sc_hd__nand3_4 _28540_ (.A(_22164_),
    .B(_22075_),
    .C(_22078_),
    .Y(_22165_));
 sky130_vsdinv _28541_ (.A(_22165_),
    .Y(_22166_));
 sky130_fd_sc_hd__a2111oi_4 _28542_ (.A1(_22162_),
    .A2(_22101_),
    .B1(_22103_),
    .C1(_22106_),
    .D1(_22166_),
    .Y(_22167_));
 sky130_fd_sc_hd__nand4_4 _28543_ (.A(_22115_),
    .B(_22117_),
    .C(_22137_),
    .D(_22139_),
    .Y(_22168_));
 sky130_vsdinv _28544_ (.A(_22168_),
    .Y(_22169_));
 sky130_fd_sc_hd__o21ai_4 _28545_ (.A1(_22052_),
    .A2(_22119_),
    .B1(_22169_),
    .Y(_22170_));
 sky130_fd_sc_hd__maj3_4 _28546_ (.A(_22138_),
    .B(_22116_),
    .C(_22142_),
    .X(_22171_));
 sky130_fd_sc_hd__xor2_4 _28547_ (.A(\decoded_imm_uj[6] ),
    .B(_22160_),
    .X(_22172_));
 sky130_vsdinv _28548_ (.A(_22172_),
    .Y(_22173_));
 sky130_fd_sc_hd__a21oi_4 _28549_ (.A1(_22170_),
    .A2(_22171_),
    .B1(_22173_),
    .Y(_22174_));
 sky130_fd_sc_hd__and3_4 _28550_ (.A(_22170_),
    .B(_22173_),
    .C(_22171_),
    .X(_22175_));
 sky130_fd_sc_hd__buf_1 _28551_ (.A(_18540_),
    .X(_22176_));
 sky130_fd_sc_hd__o21a_4 _28552_ (.A1(_22174_),
    .A2(_22175_),
    .B1(_22176_),
    .X(_22177_));
 sky130_fd_sc_hd__a2111oi_4 _28553_ (.A1(_22112_),
    .A2(_22162_),
    .B1(_21959_),
    .C1(_22113_),
    .D1(_22177_),
    .Y(_22178_));
 sky130_fd_sc_hd__o21ai_4 _28554_ (.A1(_22167_),
    .A2(_22178_),
    .B1(_22125_),
    .Y(_22179_));
 sky130_fd_sc_hd__a21oi_4 _28555_ (.A1(_22085_),
    .A2(_22160_),
    .B1(_22127_),
    .Y(_22180_));
 sky130_fd_sc_hd__buf_1 _28556_ (.A(_19115_),
    .X(_22181_));
 sky130_fd_sc_hd__o21ai_4 _28557_ (.A1(_22181_),
    .A2(\reg_next_pc[6] ),
    .B1(_22129_),
    .Y(_22182_));
 sky130_fd_sc_hd__a21oi_4 _28558_ (.A1(_22179_),
    .A2(_22180_),
    .B1(_22182_),
    .Y(_00526_));
 sky130_fd_sc_hd__buf_1 _28559_ (.A(_21922_),
    .X(_22183_));
 sky130_fd_sc_hd__buf_1 _28560_ (.A(_22043_),
    .X(_22184_));
 sky130_fd_sc_hd__or2_4 _28561_ (.A(_22044_),
    .B(\reg_out[7] ),
    .X(_22185_));
 sky130_fd_sc_hd__o21a_4 _28562_ (.A1(_22184_),
    .A2(\alu_out_q[7] ),
    .B1(_22185_),
    .X(_22186_));
 sky130_fd_sc_hd__nand2_4 _28563_ (.A(_22186_),
    .B(_21912_),
    .Y(_22187_));
 sky130_fd_sc_hd__buf_1 _28564_ (.A(_22048_),
    .X(_22188_));
 sky130_fd_sc_hd__nand3_4 _28565_ (.A(_22188_),
    .B(\reg_next_pc[7] ),
    .C(_22049_),
    .Y(_22189_));
 sky130_fd_sc_hd__nand2_4 _28566_ (.A(_22187_),
    .B(_22189_),
    .Y(_22190_));
 sky130_fd_sc_hd__buf_1 _28567_ (.A(_22190_),
    .X(_22191_));
 sky130_vsdinv _28568_ (.A(_22191_),
    .Y(_22192_));
 sky130_fd_sc_hd__nor2_4 _28569_ (.A(_22164_),
    .B(_22161_),
    .Y(_22193_));
 sky130_fd_sc_hd__xor2_4 _28570_ (.A(_22192_),
    .B(_22193_),
    .X(_22194_));
 sky130_fd_sc_hd__buf_1 _28571_ (.A(_22066_),
    .X(_22195_));
 sky130_fd_sc_hd__buf_1 _28572_ (.A(_22195_),
    .X(_22196_));
 sky130_fd_sc_hd__buf_1 _28573_ (.A(_22110_),
    .X(_22197_));
 sky130_vsdinv _28574_ (.A(\decoded_imm_uj[6] ),
    .Y(_22198_));
 sky130_fd_sc_hd__a21oi_4 _28575_ (.A1(_22158_),
    .A2(_22159_),
    .B1(_22198_),
    .Y(_22199_));
 sky130_fd_sc_hd__xor2_4 _28576_ (.A(\decoded_imm_uj[7] ),
    .B(_22190_),
    .X(_22200_));
 sky130_vsdinv _28577_ (.A(_22200_),
    .Y(_22201_));
 sky130_fd_sc_hd__nor3_4 _28578_ (.A(_22199_),
    .B(_22201_),
    .C(_22174_),
    .Y(_22202_));
 sky130_fd_sc_hd__o21a_4 _28579_ (.A1(_22199_),
    .A2(_22174_),
    .B1(_22201_),
    .X(_22203_));
 sky130_fd_sc_hd__nor3_4 _28580_ (.A(_22197_),
    .B(_22202_),
    .C(_22203_),
    .Y(_22204_));
 sky130_fd_sc_hd__a211o_4 _28581_ (.A1(_22183_),
    .A2(_22194_),
    .B1(_22196_),
    .C1(_22204_),
    .X(_22205_));
 sky130_fd_sc_hd__buf_1 _28582_ (.A(_18407_),
    .X(_22206_));
 sky130_fd_sc_hd__buf_1 _28583_ (.A(_22074_),
    .X(_22207_));
 sky130_fd_sc_hd__buf_1 _28584_ (.A(_22077_),
    .X(_22208_));
 sky130_fd_sc_hd__nand3_4 _28585_ (.A(_22207_),
    .B(_22208_),
    .C(_22192_),
    .Y(_22209_));
 sky130_vsdinv _28586_ (.A(_22209_),
    .Y(_22210_));
 sky130_fd_sc_hd__a211o_4 _28587_ (.A1(_22194_),
    .A2(_22071_),
    .B1(_22206_),
    .C1(_22210_),
    .X(_22211_));
 sky130_fd_sc_hd__a21o_4 _28588_ (.A1(_22205_),
    .A2(_22211_),
    .B1(_22039_),
    .X(_22212_));
 sky130_fd_sc_hd__buf_1 _28589_ (.A(_22084_),
    .X(_22213_));
 sky130_fd_sc_hd__a21oi_4 _28590_ (.A1(_22213_),
    .A2(_22191_),
    .B1(_22127_),
    .Y(_22214_));
 sky130_fd_sc_hd__o21ai_4 _28591_ (.A1(_22181_),
    .A2(\reg_next_pc[7] ),
    .B1(_22129_),
    .Y(_22215_));
 sky130_fd_sc_hd__a21oi_4 _28592_ (.A1(_22212_),
    .A2(_22214_),
    .B1(_22215_),
    .Y(_00527_));
 sky130_fd_sc_hd__buf_1 _28593_ (.A(_21962_),
    .X(_22216_));
 sky130_fd_sc_hd__or2_4 _28594_ (.A(_22131_),
    .B(\reg_out[8] ),
    .X(_22217_));
 sky130_fd_sc_hd__o21a_4 _28595_ (.A1(_22184_),
    .A2(\alu_out_q[8] ),
    .B1(_22217_),
    .X(_22218_));
 sky130_fd_sc_hd__o21a_4 _28596_ (.A1(_22216_),
    .A2(_22218_),
    .B1(_21967_),
    .X(_22219_));
 sky130_fd_sc_hd__o21ai_4 _28597_ (.A1(_21961_),
    .A2(_22219_),
    .B1(\reg_next_pc[8] ),
    .Y(_22220_));
 sky130_fd_sc_hd__buf_1 _28598_ (.A(_21967_),
    .X(_22221_));
 sky130_fd_sc_hd__nand3_4 _28599_ (.A(_22218_),
    .B(_22221_),
    .C(_21968_),
    .Y(_22222_));
 sky130_fd_sc_hd__and2_4 _28600_ (.A(_22220_),
    .B(_22222_),
    .X(_22223_));
 sky130_fd_sc_hd__buf_1 _28601_ (.A(_22223_),
    .X(_22224_));
 sky130_fd_sc_hd__nor3_4 _28602_ (.A(_22163_),
    .B(_22192_),
    .C(_22161_),
    .Y(_22225_));
 sky130_fd_sc_hd__xor2_4 _28603_ (.A(_22224_),
    .B(_22225_),
    .X(_22226_));
 sky130_fd_sc_hd__and3_4 _28604_ (.A(_22220_),
    .B(_22107_),
    .C(_22222_),
    .X(_22227_));
 sky130_fd_sc_hd__a2111oi_4 _28605_ (.A1(_22226_),
    .A2(_22101_),
    .B1(_22103_),
    .C1(_22106_),
    .D1(_22227_),
    .Y(_22228_));
 sky130_fd_sc_hd__buf_1 _28606_ (.A(_21958_),
    .X(_22229_));
 sky130_vsdinv _28607_ (.A(\decoded_imm_uj[8] ),
    .Y(_22230_));
 sky130_fd_sc_hd__a21o_4 _28608_ (.A1(_22220_),
    .A2(_22222_),
    .B1(_22230_),
    .X(_22231_));
 sky130_fd_sc_hd__buf_1 _28609_ (.A(_22231_),
    .X(_22232_));
 sky130_fd_sc_hd__nand3_4 _28610_ (.A(_22220_),
    .B(_22230_),
    .C(_22222_),
    .Y(_22233_));
 sky130_fd_sc_hd__maj3_4 _28611_ (.A(\decoded_imm_uj[7] ),
    .B(_22199_),
    .C(_22191_),
    .X(_22234_));
 sky130_fd_sc_hd__and2_4 _28612_ (.A(_22172_),
    .B(_22200_),
    .X(_22235_));
 sky130_fd_sc_hd__a21boi_4 _28613_ (.A1(_22170_),
    .A2(_22171_),
    .B1_N(_22235_),
    .Y(_22236_));
 sky130_fd_sc_hd__a211o_4 _28614_ (.A1(_22232_),
    .A2(_22233_),
    .B1(_22234_),
    .C1(_22236_),
    .X(_22237_));
 sky130_fd_sc_hd__and2_4 _28615_ (.A(_22231_),
    .B(_22233_),
    .X(_22238_));
 sky130_fd_sc_hd__o21ai_4 _28616_ (.A1(_22234_),
    .A2(_22236_),
    .B1(_22238_),
    .Y(_22239_));
 sky130_fd_sc_hd__a21oi_4 _28617_ (.A1(_22237_),
    .A2(_22239_),
    .B1(_22122_),
    .Y(_22240_));
 sky130_fd_sc_hd__a2111oi_4 _28618_ (.A1(_22112_),
    .A2(_22226_),
    .B1(_22229_),
    .C1(_22113_),
    .D1(_22240_),
    .Y(_22241_));
 sky130_fd_sc_hd__o21ai_4 _28619_ (.A1(_22228_),
    .A2(_22241_),
    .B1(_22125_),
    .Y(_22242_));
 sky130_vsdinv _28620_ (.A(_22224_),
    .Y(_22243_));
 sky130_fd_sc_hd__buf_1 _28621_ (.A(_18551_),
    .X(_22244_));
 sky130_fd_sc_hd__a21oi_4 _28622_ (.A1(_22213_),
    .A2(_22243_),
    .B1(_22244_),
    .Y(_22245_));
 sky130_fd_sc_hd__buf_1 _28623_ (.A(_19125_),
    .X(_22246_));
 sky130_fd_sc_hd__o21ai_4 _28624_ (.A1(_22181_),
    .A2(\reg_next_pc[8] ),
    .B1(_22246_),
    .Y(_22247_));
 sky130_fd_sc_hd__a21oi_4 _28625_ (.A1(_22242_),
    .A2(_22245_),
    .B1(_22247_),
    .Y(_00528_));
 sky130_fd_sc_hd__buf_1 _28626_ (.A(_22131_),
    .X(_22248_));
 sky130_fd_sc_hd__or2_4 _28627_ (.A(\alu_out_q[9] ),
    .B(_22043_),
    .X(_22249_));
 sky130_fd_sc_hd__o21a_4 _28628_ (.A1(_22248_),
    .A2(\reg_out[9] ),
    .B1(_22249_),
    .X(_22250_));
 sky130_fd_sc_hd__nand2_4 _28629_ (.A(_22250_),
    .B(_21912_),
    .Y(_22251_));
 sky130_fd_sc_hd__buf_1 _28630_ (.A(_22049_),
    .X(_22252_));
 sky130_fd_sc_hd__nand3_4 _28631_ (.A(_22188_),
    .B(\reg_next_pc[9] ),
    .C(_22252_),
    .Y(_22253_));
 sky130_fd_sc_hd__nand2_4 _28632_ (.A(_22251_),
    .B(_22253_),
    .Y(_22254_));
 sky130_fd_sc_hd__nand2_4 _28633_ (.A(_22254_),
    .B(\decoded_imm_uj[9] ),
    .Y(_22255_));
 sky130_vsdinv _28634_ (.A(\decoded_imm_uj[9] ),
    .Y(_22256_));
 sky130_fd_sc_hd__nand3_4 _28635_ (.A(_22251_),
    .B(_22256_),
    .C(_22253_),
    .Y(_22257_));
 sky130_fd_sc_hd__and2_4 _28636_ (.A(_22255_),
    .B(_22257_),
    .X(_22258_));
 sky130_fd_sc_hd__a21oi_4 _28637_ (.A1(_22239_),
    .A2(_22232_),
    .B1(_22258_),
    .Y(_22259_));
 sky130_fd_sc_hd__buf_1 _28638_ (.A(_22110_),
    .X(_22260_));
 sky130_fd_sc_hd__a41o_4 _28639_ (.A1(_22239_),
    .A2(_22232_),
    .A3(_22255_),
    .A4(_22257_),
    .B1(_22260_),
    .X(_22261_));
 sky130_vsdinv _28640_ (.A(_22254_),
    .Y(_22262_));
 sky130_fd_sc_hd__buf_1 _28641_ (.A(_22262_),
    .X(_22263_));
 sky130_fd_sc_hd__a2111oi_4 _28642_ (.A1(_22187_),
    .A2(_22189_),
    .B1(_22164_),
    .C1(_22224_),
    .D1(_22161_),
    .Y(_22264_));
 sky130_fd_sc_hd__xor2_4 _28643_ (.A(_22263_),
    .B(_22264_),
    .X(_22265_));
 sky130_fd_sc_hd__buf_1 _28644_ (.A(_21986_),
    .X(_22266_));
 sky130_fd_sc_hd__a21oi_4 _28645_ (.A1(_22265_),
    .A2(_22266_),
    .B1(_22145_),
    .Y(_22267_));
 sky130_fd_sc_hd__o21ai_4 _28646_ (.A1(_22259_),
    .A2(_22261_),
    .B1(_22267_),
    .Y(_22268_));
 sky130_fd_sc_hd__buf_1 _28647_ (.A(_22074_),
    .X(_22269_));
 sky130_fd_sc_hd__buf_1 _28648_ (.A(_22077_),
    .X(_22270_));
 sky130_fd_sc_hd__nand3_4 _28649_ (.A(_22263_),
    .B(_22269_),
    .C(_22270_),
    .Y(_22271_));
 sky130_vsdinv _28650_ (.A(_22271_),
    .Y(_22272_));
 sky130_fd_sc_hd__a211o_4 _28651_ (.A1(_22265_),
    .A2(_22071_),
    .B1(_22206_),
    .C1(_22272_),
    .X(_22273_));
 sky130_fd_sc_hd__buf_1 _28652_ (.A(_18547_),
    .X(_22274_));
 sky130_fd_sc_hd__a21o_4 _28653_ (.A1(_22268_),
    .A2(_22273_),
    .B1(_22274_),
    .X(_22275_));
 sky130_fd_sc_hd__buf_1 _28654_ (.A(_22254_),
    .X(_22276_));
 sky130_fd_sc_hd__a21oi_4 _28655_ (.A1(_22213_),
    .A2(_22276_),
    .B1(_22244_),
    .Y(_22277_));
 sky130_fd_sc_hd__o21ai_4 _28656_ (.A1(_22181_),
    .A2(\reg_next_pc[9] ),
    .B1(_22246_),
    .Y(_22278_));
 sky130_fd_sc_hd__a21oi_4 _28657_ (.A1(_22275_),
    .A2(_22277_),
    .B1(_22278_),
    .Y(_00529_));
 sky130_fd_sc_hd__buf_1 _28658_ (.A(_22248_),
    .X(_22279_));
 sky130_fd_sc_hd__buf_1 _28659_ (.A(_22184_),
    .X(_22280_));
 sky130_fd_sc_hd__or2_4 _28660_ (.A(\alu_out_q[10] ),
    .B(_22280_),
    .X(_22281_));
 sky130_fd_sc_hd__o21a_4 _28661_ (.A1(_22279_),
    .A2(\reg_out[10] ),
    .B1(_22281_),
    .X(_22282_));
 sky130_fd_sc_hd__nand2_4 _28662_ (.A(_22282_),
    .B(_21912_),
    .Y(_22283_));
 sky130_fd_sc_hd__nand3_4 _28663_ (.A(_22188_),
    .B(\reg_next_pc[10] ),
    .C(_22252_),
    .Y(_22284_));
 sky130_fd_sc_hd__nand2_4 _28664_ (.A(_22283_),
    .B(_22284_),
    .Y(_22285_));
 sky130_fd_sc_hd__buf_1 _28665_ (.A(_22285_),
    .X(_22286_));
 sky130_vsdinv _28666_ (.A(_22286_),
    .Y(_22287_));
 sky130_fd_sc_hd__and4_4 _28667_ (.A(_22193_),
    .B(_22191_),
    .C(_22243_),
    .D(_22276_),
    .X(_22288_));
 sky130_fd_sc_hd__xor2_4 _28668_ (.A(_22287_),
    .B(_22288_),
    .X(_22289_));
 sky130_fd_sc_hd__buf_1 _28669_ (.A(_22100_),
    .X(_22290_));
 sky130_fd_sc_hd__buf_1 _28670_ (.A(_22102_),
    .X(_22291_));
 sky130_fd_sc_hd__nand3_4 _28671_ (.A(_22287_),
    .B(_22075_),
    .C(_22078_),
    .Y(_22292_));
 sky130_vsdinv _28672_ (.A(_22292_),
    .Y(_22293_));
 sky130_fd_sc_hd__a2111oi_4 _28673_ (.A1(_22289_),
    .A2(_22290_),
    .B1(_22291_),
    .C1(_22106_),
    .D1(_22293_),
    .Y(_22294_));
 sky130_fd_sc_hd__nand3_4 _28674_ (.A(_22231_),
    .B(_22233_),
    .C(_22258_),
    .Y(_22295_));
 sky130_vsdinv _28675_ (.A(_22295_),
    .Y(_22296_));
 sky130_fd_sc_hd__o21ai_4 _28676_ (.A1(_22234_),
    .A2(_22236_),
    .B1(_22296_),
    .Y(_22297_));
 sky130_fd_sc_hd__buf_1 _28677_ (.A(_22256_),
    .X(_22298_));
 sky130_fd_sc_hd__maj3_4 _28678_ (.A(_22298_),
    .B(_22231_),
    .C(_22262_),
    .X(_22299_));
 sky130_fd_sc_hd__xor2_4 _28679_ (.A(\decoded_imm_uj[10] ),
    .B(_22285_),
    .X(_22300_));
 sky130_fd_sc_hd__a21boi_4 _28680_ (.A1(_22297_),
    .A2(_22299_),
    .B1_N(_22300_),
    .Y(_22301_));
 sky130_fd_sc_hd__a21oi_4 _28681_ (.A1(_22298_),
    .A2(_22263_),
    .B1(_22232_),
    .Y(_22302_));
 sky130_fd_sc_hd__o21a_4 _28682_ (.A1(_22234_),
    .A2(_22236_),
    .B1(_22296_),
    .X(_22303_));
 sky130_fd_sc_hd__a2111oi_4 _28683_ (.A1(\decoded_imm_uj[9] ),
    .A2(_22276_),
    .B1(_22300_),
    .C1(_22302_),
    .D1(_22303_),
    .Y(_22304_));
 sky130_fd_sc_hd__or3_4 _28684_ (.A(_22260_),
    .B(_22301_),
    .C(_22304_),
    .X(_22305_));
 sky130_fd_sc_hd__buf_1 _28685_ (.A(_18774_),
    .X(_22306_));
 sky130_fd_sc_hd__or2_4 _28686_ (.A(_22306_),
    .B(_22289_),
    .X(_22307_));
 sky130_fd_sc_hd__buf_1 _28687_ (.A(_22066_),
    .X(_22308_));
 sky130_fd_sc_hd__buf_1 _28688_ (.A(_22308_),
    .X(_22309_));
 sky130_fd_sc_hd__a21oi_4 _28689_ (.A1(_22305_),
    .A2(_22307_),
    .B1(_22309_),
    .Y(_22310_));
 sky130_fd_sc_hd__buf_1 _28690_ (.A(_21948_),
    .X(_22311_));
 sky130_fd_sc_hd__o21ai_4 _28691_ (.A1(_22294_),
    .A2(_22310_),
    .B1(_22311_),
    .Y(_22312_));
 sky130_fd_sc_hd__a21oi_4 _28692_ (.A1(_22213_),
    .A2(_22286_),
    .B1(_22244_),
    .Y(_22313_));
 sky130_fd_sc_hd__buf_1 _28693_ (.A(_19114_),
    .X(_22314_));
 sky130_fd_sc_hd__buf_1 _28694_ (.A(_22314_),
    .X(_22315_));
 sky130_fd_sc_hd__o21ai_4 _28695_ (.A1(_22315_),
    .A2(\reg_next_pc[10] ),
    .B1(_22246_),
    .Y(_22316_));
 sky130_fd_sc_hd__a21oi_4 _28696_ (.A1(_22312_),
    .A2(_22313_),
    .B1(_22316_),
    .Y(_00499_));
 sky130_fd_sc_hd__or2_4 _28697_ (.A(_22248_),
    .B(\reg_out[11] ),
    .X(_22317_));
 sky130_fd_sc_hd__o21a_4 _28698_ (.A1(_22280_),
    .A2(\alu_out_q[11] ),
    .B1(_22317_),
    .X(_22318_));
 sky130_fd_sc_hd__nand2_4 _28699_ (.A(_22318_),
    .B(_21913_),
    .Y(_22319_));
 sky130_fd_sc_hd__buf_1 _28700_ (.A(_22188_),
    .X(_22320_));
 sky130_fd_sc_hd__nand3_4 _28701_ (.A(_22320_),
    .B(\reg_next_pc[11] ),
    .C(_22252_),
    .Y(_22321_));
 sky130_fd_sc_hd__nand2_4 _28702_ (.A(_22319_),
    .B(_22321_),
    .Y(_22322_));
 sky130_fd_sc_hd__nand4_4 _28703_ (.A(_22225_),
    .B(_22243_),
    .C(_22276_),
    .D(_22286_),
    .Y(_22323_));
 sky130_fd_sc_hd__xor2_4 _28704_ (.A(_22322_),
    .B(_22323_),
    .X(_22324_));
 sky130_fd_sc_hd__buf_1 _28705_ (.A(_22105_),
    .X(_22325_));
 sky130_fd_sc_hd__buf_1 _28706_ (.A(_22269_),
    .X(_22326_));
 sky130_fd_sc_hd__buf_1 _28707_ (.A(_22270_),
    .X(_22327_));
 sky130_vsdinv _28708_ (.A(_22322_),
    .Y(_22328_));
 sky130_fd_sc_hd__buf_1 _28709_ (.A(_22328_),
    .X(_22329_));
 sky130_fd_sc_hd__nand3_4 _28710_ (.A(_22326_),
    .B(_22327_),
    .C(_22329_),
    .Y(_22330_));
 sky130_vsdinv _28711_ (.A(_22330_),
    .Y(_22331_));
 sky130_fd_sc_hd__a2111oi_4 _28712_ (.A1(_22324_),
    .A2(_22290_),
    .B1(_22291_),
    .C1(_22325_),
    .D1(_22331_),
    .Y(_22332_));
 sky130_fd_sc_hd__xor2_4 _28713_ (.A(\decoded_imm_uj[11] ),
    .B(_22322_),
    .X(_22333_));
 sky130_fd_sc_hd__a211o_4 _28714_ (.A1(\decoded_imm_uj[10] ),
    .A2(_22286_),
    .B1(_22333_),
    .C1(_22301_),
    .X(_22334_));
 sky130_vsdinv _28715_ (.A(\decoded_imm_uj[10] ),
    .Y(_22335_));
 sky130_fd_sc_hd__a21oi_4 _28716_ (.A1(_22283_),
    .A2(_22284_),
    .B1(_22335_),
    .Y(_22336_));
 sky130_fd_sc_hd__o21ai_4 _28717_ (.A1(_22336_),
    .A2(_22301_),
    .B1(_22333_),
    .Y(_22337_));
 sky130_fd_sc_hd__nand3_4 _28718_ (.A(_22334_),
    .B(_18776_),
    .C(_22337_),
    .Y(_22338_));
 sky130_fd_sc_hd__or2_4 _28719_ (.A(_22306_),
    .B(_22324_),
    .X(_22339_));
 sky130_fd_sc_hd__a21oi_4 _28720_ (.A1(_22338_),
    .A2(_22339_),
    .B1(_22309_),
    .Y(_22340_));
 sky130_fd_sc_hd__o21ai_4 _28721_ (.A1(_22332_),
    .A2(_22340_),
    .B1(_22311_),
    .Y(_22341_));
 sky130_fd_sc_hd__buf_1 _28722_ (.A(_22084_),
    .X(_22342_));
 sky130_fd_sc_hd__a21oi_4 _28723_ (.A1(_22342_),
    .A2(_22322_),
    .B1(_22244_),
    .Y(_22343_));
 sky130_fd_sc_hd__o21ai_4 _28724_ (.A1(_22315_),
    .A2(\reg_next_pc[11] ),
    .B1(_22246_),
    .Y(_22344_));
 sky130_fd_sc_hd__a21oi_4 _28725_ (.A1(_22341_),
    .A2(_22343_),
    .B1(_22344_),
    .Y(_00500_));
 sky130_fd_sc_hd__or2_4 _28726_ (.A(_22248_),
    .B(\reg_out[12] ),
    .X(_22345_));
 sky130_fd_sc_hd__o21a_4 _28727_ (.A1(_22184_),
    .A2(\alu_out_q[12] ),
    .B1(_22345_),
    .X(_22346_));
 sky130_fd_sc_hd__o21a_4 _28728_ (.A1(_22216_),
    .A2(_22346_),
    .B1(_21967_),
    .X(_22347_));
 sky130_fd_sc_hd__o21ai_4 _28729_ (.A1(_21961_),
    .A2(_22347_),
    .B1(\reg_next_pc[12] ),
    .Y(_22348_));
 sky130_fd_sc_hd__buf_1 _28730_ (.A(_21968_),
    .X(_22349_));
 sky130_fd_sc_hd__nand3_4 _28731_ (.A(_22346_),
    .B(_22221_),
    .C(_22349_),
    .Y(_22350_));
 sky130_fd_sc_hd__and2_4 _28732_ (.A(_22348_),
    .B(_22350_),
    .X(_22351_));
 sky130_fd_sc_hd__buf_1 _28733_ (.A(_22351_),
    .X(_22352_));
 sky130_fd_sc_hd__buf_1 _28734_ (.A(_22352_),
    .X(_22353_));
 sky130_fd_sc_hd__nor2_4 _28735_ (.A(_22328_),
    .B(_22323_),
    .Y(_22354_));
 sky130_fd_sc_hd__xor2_4 _28736_ (.A(_22353_),
    .B(_22354_),
    .X(_22355_));
 sky130_fd_sc_hd__and3_4 _28737_ (.A(_22348_),
    .B(_22107_),
    .C(_22350_),
    .X(_22356_));
 sky130_fd_sc_hd__a2111oi_4 _28738_ (.A1(_22355_),
    .A2(_22290_),
    .B1(_22291_),
    .C1(_22325_),
    .D1(_22356_),
    .Y(_22357_));
 sky130_vsdinv _28739_ (.A(\decoded_imm_uj[11] ),
    .Y(_22358_));
 sky130_fd_sc_hd__a21oi_4 _28740_ (.A1(_22319_),
    .A2(_22321_),
    .B1(_22358_),
    .Y(_22359_));
 sky130_vsdinv _28741_ (.A(_22359_),
    .Y(_22360_));
 sky130_vsdinv _28742_ (.A(\decoded_imm_uj[12] ),
    .Y(_22361_));
 sky130_fd_sc_hd__xor2_4 _28743_ (.A(_22361_),
    .B(_22352_),
    .X(_22362_));
 sky130_vsdinv _28744_ (.A(_22362_),
    .Y(_22363_));
 sky130_fd_sc_hd__a21oi_4 _28745_ (.A1(_22337_),
    .A2(_22360_),
    .B1(_22363_),
    .Y(_22364_));
 sky130_fd_sc_hd__and3_4 _28746_ (.A(_22337_),
    .B(_22360_),
    .C(_22363_),
    .X(_22365_));
 sky130_fd_sc_hd__or3_4 _28747_ (.A(_22260_),
    .B(_22364_),
    .C(_22365_),
    .X(_22366_));
 sky130_fd_sc_hd__or2_4 _28748_ (.A(_22306_),
    .B(_22355_),
    .X(_22367_));
 sky130_fd_sc_hd__a21oi_4 _28749_ (.A1(_22366_),
    .A2(_22367_),
    .B1(_22309_),
    .Y(_22368_));
 sky130_fd_sc_hd__o21ai_4 _28750_ (.A1(_22357_),
    .A2(_22368_),
    .B1(_22311_),
    .Y(_22369_));
 sky130_vsdinv _28751_ (.A(_22353_),
    .Y(_22370_));
 sky130_fd_sc_hd__buf_1 _28752_ (.A(_19080_),
    .X(_22371_));
 sky130_fd_sc_hd__buf_1 _28753_ (.A(_22371_),
    .X(_22372_));
 sky130_fd_sc_hd__a21oi_4 _28754_ (.A1(_22342_),
    .A2(_22370_),
    .B1(_22372_),
    .Y(_22373_));
 sky130_fd_sc_hd__buf_1 _28755_ (.A(_18536_),
    .X(_22374_));
 sky130_fd_sc_hd__buf_1 _28756_ (.A(_22374_),
    .X(_22375_));
 sky130_fd_sc_hd__o21ai_4 _28757_ (.A1(_22315_),
    .A2(\reg_next_pc[12] ),
    .B1(_22375_),
    .Y(_22376_));
 sky130_fd_sc_hd__a21oi_4 _28758_ (.A1(_22369_),
    .A2(_22373_),
    .B1(_22376_),
    .Y(_00501_));
 sky130_fd_sc_hd__buf_1 _28759_ (.A(_22280_),
    .X(_22377_));
 sky130_fd_sc_hd__or2_4 _28760_ (.A(_22279_),
    .B(\reg_out[13] ),
    .X(_22378_));
 sky130_fd_sc_hd__o21a_4 _28761_ (.A1(_22377_),
    .A2(\alu_out_q[13] ),
    .B1(_22378_),
    .X(_22379_));
 sky130_fd_sc_hd__nand2_4 _28762_ (.A(_22379_),
    .B(_21913_),
    .Y(_22380_));
 sky130_fd_sc_hd__buf_1 _28763_ (.A(_22252_),
    .X(_22381_));
 sky130_fd_sc_hd__nand3_4 _28764_ (.A(_22320_),
    .B(\reg_next_pc[13] ),
    .C(_22381_),
    .Y(_22382_));
 sky130_fd_sc_hd__nand2_4 _28765_ (.A(_22380_),
    .B(_22382_),
    .Y(_22383_));
 sky130_fd_sc_hd__buf_1 _28766_ (.A(_22383_),
    .X(_22384_));
 sky130_vsdinv _28767_ (.A(_22384_),
    .Y(_22385_));
 sky130_fd_sc_hd__nor3_4 _28768_ (.A(_22329_),
    .B(_22353_),
    .C(_22323_),
    .Y(_22386_));
 sky130_fd_sc_hd__xor2_4 _28769_ (.A(_22385_),
    .B(_22386_),
    .X(_22387_));
 sky130_fd_sc_hd__nand3_4 _28770_ (.A(_22326_),
    .B(_22327_),
    .C(_22385_),
    .Y(_22388_));
 sky130_vsdinv _28771_ (.A(_22388_),
    .Y(_22389_));
 sky130_fd_sc_hd__a2111oi_4 _28772_ (.A1(_22387_),
    .A2(_22290_),
    .B1(_22291_),
    .C1(_22325_),
    .D1(_22389_),
    .Y(_22390_));
 sky130_fd_sc_hd__xor2_4 _28773_ (.A(\decoded_imm_uj[13] ),
    .B(_22383_),
    .X(_22391_));
 sky130_fd_sc_hd__a211o_4 _28774_ (.A1(\decoded_imm_uj[12] ),
    .A2(_22370_),
    .B1(_22391_),
    .C1(_22364_),
    .X(_22392_));
 sky130_fd_sc_hd__a21oi_4 _28775_ (.A1(_22348_),
    .A2(_22350_),
    .B1(_22361_),
    .Y(_22393_));
 sky130_fd_sc_hd__o21ai_4 _28776_ (.A1(_22393_),
    .A2(_22364_),
    .B1(_22391_),
    .Y(_22394_));
 sky130_fd_sc_hd__nand3_4 _28777_ (.A(_22392_),
    .B(_18776_),
    .C(_22394_),
    .Y(_22395_));
 sky130_fd_sc_hd__or2_4 _28778_ (.A(_22057_),
    .B(_22387_),
    .X(_22396_));
 sky130_fd_sc_hd__a21oi_4 _28779_ (.A1(_22395_),
    .A2(_22396_),
    .B1(_22309_),
    .Y(_22397_));
 sky130_fd_sc_hd__o21ai_4 _28780_ (.A1(_22390_),
    .A2(_22397_),
    .B1(_22311_),
    .Y(_22398_));
 sky130_fd_sc_hd__a21oi_4 _28781_ (.A1(_22342_),
    .A2(_22384_),
    .B1(_22372_),
    .Y(_22399_));
 sky130_fd_sc_hd__o21ai_4 _28782_ (.A1(_22315_),
    .A2(\reg_next_pc[13] ),
    .B1(_22375_),
    .Y(_22400_));
 sky130_fd_sc_hd__a21oi_4 _28783_ (.A1(_22398_),
    .A2(_22399_),
    .B1(_22400_),
    .Y(_00502_));
 sky130_fd_sc_hd__buf_1 _28784_ (.A(_21961_),
    .X(_22401_));
 sky130_fd_sc_hd__or2_4 _28785_ (.A(\alu_out_q[14] ),
    .B(_22280_),
    .X(_22402_));
 sky130_fd_sc_hd__o21a_4 _28786_ (.A1(_22279_),
    .A2(\reg_out[14] ),
    .B1(_22402_),
    .X(_22403_));
 sky130_fd_sc_hd__o21a_4 _28787_ (.A1(_22216_),
    .A2(_22403_),
    .B1(_22221_),
    .X(_22404_));
 sky130_fd_sc_hd__o21ai_4 _28788_ (.A1(_22401_),
    .A2(_22404_),
    .B1(\reg_next_pc[14] ),
    .Y(_22405_));
 sky130_fd_sc_hd__buf_1 _28789_ (.A(_22221_),
    .X(_22406_));
 sky130_fd_sc_hd__nand3_4 _28790_ (.A(_22403_),
    .B(_22406_),
    .C(_22349_),
    .Y(_22407_));
 sky130_fd_sc_hd__and2_4 _28791_ (.A(_22405_),
    .B(_22407_),
    .X(_22408_));
 sky130_fd_sc_hd__buf_1 _28792_ (.A(_22408_),
    .X(_22409_));
 sky130_fd_sc_hd__a2111oi_4 _28793_ (.A1(_22348_),
    .A2(_22350_),
    .B1(_22329_),
    .C1(_22385_),
    .D1(_22323_),
    .Y(_22410_));
 sky130_fd_sc_hd__xor2_4 _28794_ (.A(_22409_),
    .B(_22410_),
    .X(_22411_));
 sky130_fd_sc_hd__buf_1 _28795_ (.A(_22100_),
    .X(_22412_));
 sky130_fd_sc_hd__buf_1 _28796_ (.A(_22102_),
    .X(_22413_));
 sky130_fd_sc_hd__buf_1 _28797_ (.A(_22032_),
    .X(_22414_));
 sky130_fd_sc_hd__and3_4 _28798_ (.A(_22405_),
    .B(_22414_),
    .C(_22407_),
    .X(_22415_));
 sky130_fd_sc_hd__a2111oi_4 _28799_ (.A1(_22411_),
    .A2(_22412_),
    .B1(_22413_),
    .C1(_22325_),
    .D1(_22415_),
    .Y(_22416_));
 sky130_vsdinv _28800_ (.A(\decoded_imm_uj[14] ),
    .Y(_22417_));
 sky130_fd_sc_hd__xor2_4 _28801_ (.A(_22417_),
    .B(_22409_),
    .X(_22418_));
 sky130_fd_sc_hd__nand2_4 _28802_ (.A(_22384_),
    .B(\decoded_imm_uj[13] ),
    .Y(_22419_));
 sky130_fd_sc_hd__nand2_4 _28803_ (.A(_22394_),
    .B(_22419_),
    .Y(_22420_));
 sky130_fd_sc_hd__or2_4 _28804_ (.A(_22418_),
    .B(_22420_),
    .X(_22421_));
 sky130_fd_sc_hd__nand2_4 _28805_ (.A(_22420_),
    .B(_22418_),
    .Y(_22422_));
 sky130_fd_sc_hd__nand3_4 _28806_ (.A(_22421_),
    .B(_18776_),
    .C(_22422_),
    .Y(_22423_));
 sky130_fd_sc_hd__or2_4 _28807_ (.A(_22057_),
    .B(_22411_),
    .X(_22424_));
 sky130_fd_sc_hd__buf_1 _28808_ (.A(_22195_),
    .X(_22425_));
 sky130_fd_sc_hd__a21oi_4 _28809_ (.A1(_22423_),
    .A2(_22424_),
    .B1(_22425_),
    .Y(_22426_));
 sky130_fd_sc_hd__buf_1 _28810_ (.A(_21948_),
    .X(_22427_));
 sky130_fd_sc_hd__o21ai_4 _28811_ (.A1(_22416_),
    .A2(_22426_),
    .B1(_22427_),
    .Y(_22428_));
 sky130_vsdinv _28812_ (.A(_22409_),
    .Y(_22429_));
 sky130_fd_sc_hd__a21oi_4 _28813_ (.A1(_22342_),
    .A2(_22429_),
    .B1(_22372_),
    .Y(_22430_));
 sky130_fd_sc_hd__buf_1 _28814_ (.A(_22314_),
    .X(_22431_));
 sky130_fd_sc_hd__o21ai_4 _28815_ (.A1(_22431_),
    .A2(\reg_next_pc[14] ),
    .B1(_22375_),
    .Y(_22432_));
 sky130_fd_sc_hd__a21oi_4 _28816_ (.A1(_22428_),
    .A2(_22430_),
    .B1(_22432_),
    .Y(_00503_));
 sky130_fd_sc_hd__buf_1 _28817_ (.A(_22377_),
    .X(_22433_));
 sky130_fd_sc_hd__buf_1 _28818_ (.A(_22279_),
    .X(_22434_));
 sky130_fd_sc_hd__or2_4 _28819_ (.A(_22434_),
    .B(\reg_out[15] ),
    .X(_22435_));
 sky130_fd_sc_hd__o21a_4 _28820_ (.A1(_22433_),
    .A2(\alu_out_q[15] ),
    .B1(_22435_),
    .X(_22436_));
 sky130_fd_sc_hd__nand2_4 _28821_ (.A(_22436_),
    .B(_21914_),
    .Y(_22437_));
 sky130_fd_sc_hd__buf_1 _28822_ (.A(_22320_),
    .X(_22438_));
 sky130_fd_sc_hd__nand3_4 _28823_ (.A(_22438_),
    .B(\reg_next_pc[15] ),
    .C(_22381_),
    .Y(_22439_));
 sky130_fd_sc_hd__nand2_4 _28824_ (.A(_22437_),
    .B(_22439_),
    .Y(_22440_));
 sky130_fd_sc_hd__buf_1 _28825_ (.A(_22440_),
    .X(_22441_));
 sky130_fd_sc_hd__nand4_4 _28826_ (.A(_22354_),
    .B(_22370_),
    .C(_22384_),
    .D(_22429_),
    .Y(_22442_));
 sky130_fd_sc_hd__xor2_4 _28827_ (.A(_22441_),
    .B(_22442_),
    .X(_22443_));
 sky130_fd_sc_hd__a21oi_4 _28828_ (.A1(_22405_),
    .A2(_22407_),
    .B1(_22417_),
    .Y(_22444_));
 sky130_vsdinv _28829_ (.A(_22444_),
    .Y(_22445_));
 sky130_fd_sc_hd__buf_1 _28830_ (.A(\decoded_imm_uj[15] ),
    .X(_22446_));
 sky130_fd_sc_hd__xor2_4 _28831_ (.A(_22446_),
    .B(_22441_),
    .X(_22447_));
 sky130_fd_sc_hd__a21oi_4 _28832_ (.A1(_22422_),
    .A2(_22445_),
    .B1(_22447_),
    .Y(_22448_));
 sky130_fd_sc_hd__and3_4 _28833_ (.A(_22422_),
    .B(_22445_),
    .C(_22447_),
    .X(_22449_));
 sky130_fd_sc_hd__nor3_4 _28834_ (.A(_22197_),
    .B(_22448_),
    .C(_22449_),
    .Y(_22450_));
 sky130_fd_sc_hd__a211o_4 _28835_ (.A1(_22183_),
    .A2(_22443_),
    .B1(_22196_),
    .C1(_22450_),
    .X(_22451_));
 sky130_fd_sc_hd__buf_1 _28836_ (.A(_22070_),
    .X(_22452_));
 sky130_vsdinv _28837_ (.A(_22441_),
    .Y(_22453_));
 sky130_fd_sc_hd__buf_1 _28838_ (.A(_22453_),
    .X(_22454_));
 sky130_fd_sc_hd__nand3_4 _28839_ (.A(_22207_),
    .B(_22208_),
    .C(_22454_),
    .Y(_22455_));
 sky130_vsdinv _28840_ (.A(_22455_),
    .Y(_22456_));
 sky130_fd_sc_hd__a211o_4 _28841_ (.A1(_22443_),
    .A2(_22452_),
    .B1(_22206_),
    .C1(_22456_),
    .X(_22457_));
 sky130_fd_sc_hd__a21o_4 _28842_ (.A1(_22451_),
    .A2(_22457_),
    .B1(_22274_),
    .X(_22458_));
 sky130_fd_sc_hd__buf_1 _28843_ (.A(_22083_),
    .X(_22459_));
 sky130_fd_sc_hd__buf_1 _28844_ (.A(_22459_),
    .X(_22460_));
 sky130_fd_sc_hd__a21oi_4 _28845_ (.A1(_22460_),
    .A2(_22441_),
    .B1(_22372_),
    .Y(_22461_));
 sky130_fd_sc_hd__o21ai_4 _28846_ (.A1(_22431_),
    .A2(\reg_next_pc[15] ),
    .B1(_22375_),
    .Y(_22462_));
 sky130_fd_sc_hd__a21oi_4 _28847_ (.A1(_22458_),
    .A2(_22461_),
    .B1(_22462_),
    .Y(_00504_));
 sky130_fd_sc_hd__buf_1 _28848_ (.A(_22216_),
    .X(_22463_));
 sky130_fd_sc_hd__or2_4 _28849_ (.A(_22434_),
    .B(\reg_out[16] ),
    .X(_22464_));
 sky130_fd_sc_hd__o21a_4 _28850_ (.A1(_22377_),
    .A2(\alu_out_q[16] ),
    .B1(_22464_),
    .X(_22465_));
 sky130_fd_sc_hd__o21a_4 _28851_ (.A1(_22463_),
    .A2(_22465_),
    .B1(_22406_),
    .X(_22466_));
 sky130_fd_sc_hd__o21ai_4 _28852_ (.A1(_22401_),
    .A2(_22466_),
    .B1(\reg_next_pc[16] ),
    .Y(_22467_));
 sky130_fd_sc_hd__buf_1 _28853_ (.A(_22467_),
    .X(_22468_));
 sky130_fd_sc_hd__nand3_4 _28854_ (.A(_22465_),
    .B(_22406_),
    .C(_22349_),
    .Y(_22469_));
 sky130_fd_sc_hd__buf_1 _28855_ (.A(_22469_),
    .X(_22470_));
 sky130_fd_sc_hd__and2_4 _28856_ (.A(_22468_),
    .B(_22470_),
    .X(_22471_));
 sky130_fd_sc_hd__buf_1 _28857_ (.A(_22471_),
    .X(_22472_));
 sky130_fd_sc_hd__nor2_4 _28858_ (.A(_22453_),
    .B(_22442_),
    .Y(_22473_));
 sky130_fd_sc_hd__xor2_4 _28859_ (.A(_22472_),
    .B(_22473_),
    .X(_22474_));
 sky130_fd_sc_hd__buf_1 _28860_ (.A(_22105_),
    .X(_22475_));
 sky130_fd_sc_hd__and3_4 _28861_ (.A(_22468_),
    .B(_22414_),
    .C(_22470_),
    .X(_22476_));
 sky130_fd_sc_hd__a2111oi_4 _28862_ (.A1(_22474_),
    .A2(_22412_),
    .B1(_22413_),
    .C1(_22475_),
    .D1(_22476_),
    .Y(_22477_));
 sky130_fd_sc_hd__buf_1 _28863_ (.A(_22111_),
    .X(_22478_));
 sky130_fd_sc_hd__a21oi_4 _28864_ (.A1(\decoded_imm_uj[15] ),
    .A2(_22440_),
    .B1(_22444_),
    .Y(_22479_));
 sky130_fd_sc_hd__nand2_4 _28865_ (.A(_22422_),
    .B(_22479_),
    .Y(_22480_));
 sky130_vsdinv _28866_ (.A(_22439_),
    .Y(_22481_));
 sky130_fd_sc_hd__a211o_4 _28867_ (.A1(_22436_),
    .A2(_21915_),
    .B1(_22446_),
    .C1(_22481_),
    .X(_22482_));
 sky130_vsdinv _28868_ (.A(\decoded_imm_uj[16] ),
    .Y(_22483_));
 sky130_fd_sc_hd__a21o_4 _28869_ (.A1(_22467_),
    .A2(_22469_),
    .B1(_22483_),
    .X(_22484_));
 sky130_fd_sc_hd__buf_1 _28870_ (.A(_22484_),
    .X(_22485_));
 sky130_fd_sc_hd__nand3_4 _28871_ (.A(_22468_),
    .B(_22483_),
    .C(_22470_),
    .Y(_22486_));
 sky130_fd_sc_hd__and2_4 _28872_ (.A(_22485_),
    .B(_22486_),
    .X(_22487_));
 sky130_fd_sc_hd__a21o_4 _28873_ (.A1(_22480_),
    .A2(_22482_),
    .B1(_22487_),
    .X(_22488_));
 sky130_fd_sc_hd__nand3_4 _28874_ (.A(_22480_),
    .B(_22482_),
    .C(_22487_),
    .Y(_22489_));
 sky130_fd_sc_hd__a21oi_4 _28875_ (.A1(_22488_),
    .A2(_22489_),
    .B1(_22122_),
    .Y(_22490_));
 sky130_fd_sc_hd__a2111oi_4 _28876_ (.A1(_22478_),
    .A2(_22474_),
    .B1(_22229_),
    .C1(_22113_),
    .D1(_22490_),
    .Y(_22491_));
 sky130_fd_sc_hd__o21ai_4 _28877_ (.A1(_22477_),
    .A2(_22491_),
    .B1(_22427_),
    .Y(_22492_));
 sky130_vsdinv _28878_ (.A(_22472_),
    .Y(_22493_));
 sky130_fd_sc_hd__buf_1 _28879_ (.A(_22371_),
    .X(_22494_));
 sky130_fd_sc_hd__a21oi_4 _28880_ (.A1(_22460_),
    .A2(_22493_),
    .B1(_22494_),
    .Y(_22495_));
 sky130_fd_sc_hd__buf_1 _28881_ (.A(_22374_),
    .X(_22496_));
 sky130_fd_sc_hd__o21ai_4 _28882_ (.A1(_22431_),
    .A2(\reg_next_pc[16] ),
    .B1(_22496_),
    .Y(_22497_));
 sky130_fd_sc_hd__a21oi_4 _28883_ (.A1(_22492_),
    .A2(_22495_),
    .B1(_22497_),
    .Y(_00505_));
 sky130_fd_sc_hd__buf_1 _28884_ (.A(_22434_),
    .X(_22498_));
 sky130_fd_sc_hd__or2_4 _28885_ (.A(\alu_out_q[17] ),
    .B(_22377_),
    .X(_22499_));
 sky130_fd_sc_hd__o21a_4 _28886_ (.A1(_22498_),
    .A2(\reg_out[17] ),
    .B1(_22499_),
    .X(_22500_));
 sky130_fd_sc_hd__nand2_4 _28887_ (.A(_22500_),
    .B(_21913_),
    .Y(_22501_));
 sky130_fd_sc_hd__nand3_4 _28888_ (.A(_22320_),
    .B(\reg_next_pc[17] ),
    .C(_22381_),
    .Y(_22502_));
 sky130_fd_sc_hd__nand2_4 _28889_ (.A(_22501_),
    .B(_22502_),
    .Y(_22503_));
 sky130_fd_sc_hd__xor2_4 _28890_ (.A(\decoded_imm_uj[17] ),
    .B(_22503_),
    .X(_22504_));
 sky130_fd_sc_hd__a21oi_4 _28891_ (.A1(_22489_),
    .A2(_22485_),
    .B1(_22504_),
    .Y(_22505_));
 sky130_fd_sc_hd__nand3_4 _28892_ (.A(_22489_),
    .B(_22485_),
    .C(_22504_),
    .Y(_22506_));
 sky130_fd_sc_hd__buf_1 _28893_ (.A(_18775_),
    .X(_22507_));
 sky130_fd_sc_hd__nand2_4 _28894_ (.A(_22506_),
    .B(_22507_),
    .Y(_22508_));
 sky130_fd_sc_hd__buf_1 _28895_ (.A(_22503_),
    .X(_22509_));
 sky130_vsdinv _28896_ (.A(_22509_),
    .Y(_22510_));
 sky130_fd_sc_hd__buf_1 _28897_ (.A(_22510_),
    .X(_22511_));
 sky130_fd_sc_hd__nor3_4 _28898_ (.A(_22454_),
    .B(_22472_),
    .C(_22442_),
    .Y(_22512_));
 sky130_fd_sc_hd__xor2_4 _28899_ (.A(_22511_),
    .B(_22512_),
    .X(_22513_));
 sky130_fd_sc_hd__a21oi_4 _28900_ (.A1(_22513_),
    .A2(_22266_),
    .B1(_22067_),
    .Y(_22514_));
 sky130_fd_sc_hd__o21ai_4 _28901_ (.A1(_22505_),
    .A2(_22508_),
    .B1(_22514_),
    .Y(_22515_));
 sky130_fd_sc_hd__nand3_4 _28902_ (.A(_22511_),
    .B(_22269_),
    .C(_22270_),
    .Y(_22516_));
 sky130_vsdinv _28903_ (.A(_22516_),
    .Y(_22517_));
 sky130_fd_sc_hd__a211o_4 _28904_ (.A1(_22513_),
    .A2(_22452_),
    .B1(_22206_),
    .C1(_22517_),
    .X(_22518_));
 sky130_fd_sc_hd__a21o_4 _28905_ (.A1(_22515_),
    .A2(_22518_),
    .B1(_22274_),
    .X(_22519_));
 sky130_fd_sc_hd__a21oi_4 _28906_ (.A1(_22460_),
    .A2(_22509_),
    .B1(_22494_),
    .Y(_22520_));
 sky130_fd_sc_hd__o21ai_4 _28907_ (.A1(_22431_),
    .A2(\reg_next_pc[17] ),
    .B1(_22496_),
    .Y(_22521_));
 sky130_fd_sc_hd__a21oi_4 _28908_ (.A1(_22519_),
    .A2(_22520_),
    .B1(_22521_),
    .Y(_00506_));
 sky130_fd_sc_hd__buf_1 _28909_ (.A(_22433_),
    .X(_22522_));
 sky130_fd_sc_hd__or2_4 _28910_ (.A(_22498_),
    .B(\reg_out[18] ),
    .X(_22523_));
 sky130_fd_sc_hd__o21a_4 _28911_ (.A1(_22522_),
    .A2(\alu_out_q[18] ),
    .B1(_22523_),
    .X(_22524_));
 sky130_fd_sc_hd__nand2_4 _28912_ (.A(_22524_),
    .B(_21914_),
    .Y(_22525_));
 sky130_fd_sc_hd__buf_1 _28913_ (.A(_22381_),
    .X(_22526_));
 sky130_fd_sc_hd__nand3_4 _28914_ (.A(_22438_),
    .B(\reg_next_pc[18] ),
    .C(_22526_),
    .Y(_22527_));
 sky130_fd_sc_hd__nand2_4 _28915_ (.A(_22525_),
    .B(_22527_),
    .Y(_22528_));
 sky130_fd_sc_hd__buf_1 _28916_ (.A(_22528_),
    .X(_22529_));
 sky130_vsdinv _28917_ (.A(_22529_),
    .Y(_22530_));
 sky130_fd_sc_hd__a2111oi_4 _28918_ (.A1(_22468_),
    .A2(_22470_),
    .B1(_22454_),
    .C1(_22511_),
    .D1(_22442_),
    .Y(_22531_));
 sky130_fd_sc_hd__xor2_4 _28919_ (.A(_22530_),
    .B(_22531_),
    .X(_22532_));
 sky130_fd_sc_hd__nand3_4 _28920_ (.A(_22326_),
    .B(_22327_),
    .C(_22530_),
    .Y(_22533_));
 sky130_vsdinv _28921_ (.A(_22533_),
    .Y(_22534_));
 sky130_fd_sc_hd__a2111oi_4 _28922_ (.A1(_22532_),
    .A2(_22412_),
    .B1(_22413_),
    .C1(_22475_),
    .D1(_22534_),
    .Y(_22535_));
 sky130_fd_sc_hd__xor2_4 _28923_ (.A(\decoded_imm_uj[18] ),
    .B(_22528_),
    .X(_22536_));
 sky130_fd_sc_hd__nand3_4 _28924_ (.A(_22484_),
    .B(_22486_),
    .C(_22504_),
    .Y(_22537_));
 sky130_vsdinv _28925_ (.A(_22537_),
    .Y(_22538_));
 sky130_fd_sc_hd__nand3_4 _28926_ (.A(_22480_),
    .B(_22482_),
    .C(_22538_),
    .Y(_22539_));
 sky130_vsdinv _28927_ (.A(\decoded_imm_uj[17] ),
    .Y(_22540_));
 sky130_fd_sc_hd__maj3_4 _28928_ (.A(_22540_),
    .B(_22485_),
    .C(_22510_),
    .X(_22541_));
 sky130_fd_sc_hd__nand2_4 _28929_ (.A(_22539_),
    .B(_22541_),
    .Y(_22542_));
 sky130_fd_sc_hd__xnor2_4 _28930_ (.A(_22536_),
    .B(_22542_),
    .Y(_22543_));
 sky130_fd_sc_hd__buf_1 _28931_ (.A(_22306_),
    .X(_22544_));
 sky130_fd_sc_hd__a21o_4 _28932_ (.A1(_22532_),
    .A2(_22064_),
    .B1(_22308_),
    .X(_22545_));
 sky130_fd_sc_hd__a21oi_4 _28933_ (.A1(_22543_),
    .A2(_22544_),
    .B1(_22545_),
    .Y(_22546_));
 sky130_fd_sc_hd__o21ai_4 _28934_ (.A1(_22535_),
    .A2(_22546_),
    .B1(_22427_),
    .Y(_22547_));
 sky130_fd_sc_hd__a21oi_4 _28935_ (.A1(_22460_),
    .A2(_22529_),
    .B1(_22494_),
    .Y(_22548_));
 sky130_fd_sc_hd__buf_1 _28936_ (.A(_22314_),
    .X(_22549_));
 sky130_fd_sc_hd__o21ai_4 _28937_ (.A1(_22549_),
    .A2(\reg_next_pc[18] ),
    .B1(_22496_),
    .Y(_22550_));
 sky130_fd_sc_hd__a21oi_4 _28938_ (.A1(_22547_),
    .A2(_22548_),
    .B1(_22550_),
    .Y(_00507_));
 sky130_fd_sc_hd__or2_4 _28939_ (.A(_22498_),
    .B(\reg_out[19] ),
    .X(_22551_));
 sky130_fd_sc_hd__o21a_4 _28940_ (.A1(_22522_),
    .A2(\alu_out_q[19] ),
    .B1(_22551_),
    .X(_22552_));
 sky130_fd_sc_hd__nand2_4 _28941_ (.A(_22552_),
    .B(_21914_),
    .Y(_22553_));
 sky130_fd_sc_hd__nand3_4 _28942_ (.A(_22438_),
    .B(\reg_next_pc[19] ),
    .C(_22526_),
    .Y(_22554_));
 sky130_fd_sc_hd__nand2_4 _28943_ (.A(_22553_),
    .B(_22554_),
    .Y(_22555_));
 sky130_fd_sc_hd__buf_1 _28944_ (.A(_22555_),
    .X(_22556_));
 sky130_vsdinv _28945_ (.A(_22556_),
    .Y(_22557_));
 sky130_fd_sc_hd__and4_4 _28946_ (.A(_22473_),
    .B(_22493_),
    .C(_22509_),
    .D(_22528_),
    .X(_22558_));
 sky130_fd_sc_hd__xor2_4 _28947_ (.A(_22557_),
    .B(_22558_),
    .X(_22559_));
 sky130_fd_sc_hd__xor2_4 _28948_ (.A(\decoded_imm_uj[19] ),
    .B(_22555_),
    .X(_22560_));
 sky130_fd_sc_hd__a21boi_4 _28949_ (.A1(_22525_),
    .A2(_22527_),
    .B1_N(\decoded_imm_uj[18] ),
    .Y(_22561_));
 sky130_fd_sc_hd__a21oi_4 _28950_ (.A1(_22542_),
    .A2(_22536_),
    .B1(_22561_),
    .Y(_22562_));
 sky130_fd_sc_hd__a21oi_4 _28951_ (.A1(_22562_),
    .A2(_22560_),
    .B1(_22110_),
    .Y(_22563_));
 sky130_fd_sc_hd__o21a_4 _28952_ (.A1(_22560_),
    .A2(_22562_),
    .B1(_22563_),
    .X(_22564_));
 sky130_fd_sc_hd__a211o_4 _28953_ (.A1(_22183_),
    .A2(_22559_),
    .B1(_22196_),
    .C1(_22564_),
    .X(_22565_));
 sky130_fd_sc_hd__buf_1 _28954_ (.A(_18557_),
    .X(_22566_));
 sky130_fd_sc_hd__nand3_4 _28955_ (.A(_22207_),
    .B(_22208_),
    .C(_22557_),
    .Y(_22567_));
 sky130_vsdinv _28956_ (.A(_22567_),
    .Y(_22568_));
 sky130_fd_sc_hd__a211o_4 _28957_ (.A1(_22559_),
    .A2(_22452_),
    .B1(_22566_),
    .C1(_22568_),
    .X(_22569_));
 sky130_fd_sc_hd__a21o_4 _28958_ (.A1(_22565_),
    .A2(_22569_),
    .B1(_22274_),
    .X(_22570_));
 sky130_fd_sc_hd__buf_1 _28959_ (.A(_22459_),
    .X(_22571_));
 sky130_fd_sc_hd__a21oi_4 _28960_ (.A1(_22571_),
    .A2(_22556_),
    .B1(_22494_),
    .Y(_22572_));
 sky130_fd_sc_hd__o21ai_4 _28961_ (.A1(_22549_),
    .A2(\reg_next_pc[19] ),
    .B1(_22496_),
    .Y(_22573_));
 sky130_fd_sc_hd__a21oi_4 _28962_ (.A1(_22570_),
    .A2(_22572_),
    .B1(_22573_),
    .Y(_00508_));
 sky130_fd_sc_hd__or2_4 _28963_ (.A(_22434_),
    .B(\reg_out[20] ),
    .X(_22574_));
 sky130_fd_sc_hd__o21a_4 _28964_ (.A1(_22433_),
    .A2(\alu_out_q[20] ),
    .B1(_22574_),
    .X(_22575_));
 sky130_fd_sc_hd__buf_1 _28965_ (.A(_22406_),
    .X(_22576_));
 sky130_fd_sc_hd__o21a_4 _28966_ (.A1(_22463_),
    .A2(_22575_),
    .B1(_22576_),
    .X(_22577_));
 sky130_fd_sc_hd__o21ai_4 _28967_ (.A1(_22401_),
    .A2(_22577_),
    .B1(\reg_next_pc[20] ),
    .Y(_22578_));
 sky130_fd_sc_hd__buf_1 _28968_ (.A(_22349_),
    .X(_22579_));
 sky130_fd_sc_hd__nand3_4 _28969_ (.A(_22575_),
    .B(_22576_),
    .C(_22579_),
    .Y(_22580_));
 sky130_fd_sc_hd__and2_4 _28970_ (.A(_22578_),
    .B(_22580_),
    .X(_22581_));
 sky130_fd_sc_hd__buf_1 _28971_ (.A(_22581_),
    .X(_22582_));
 sky130_fd_sc_hd__and4_4 _28972_ (.A(_22512_),
    .B(_22509_),
    .C(_22529_),
    .D(_22555_),
    .X(_22583_));
 sky130_fd_sc_hd__xor2_4 _28973_ (.A(_22582_),
    .B(_22583_),
    .X(_22584_));
 sky130_fd_sc_hd__and3_4 _28974_ (.A(_22578_),
    .B(_22414_),
    .C(_22580_),
    .X(_22585_));
 sky130_fd_sc_hd__a2111oi_4 _28975_ (.A1(_22584_),
    .A2(_22412_),
    .B1(_22413_),
    .C1(_22475_),
    .D1(_22585_),
    .Y(_22586_));
 sky130_fd_sc_hd__and2_4 _28976_ (.A(_22536_),
    .B(_22560_),
    .X(_22587_));
 sky130_vsdinv _28977_ (.A(\decoded_imm_uj[20] ),
    .Y(_22588_));
 sky130_fd_sc_hd__a21o_4 _28978_ (.A1(_22578_),
    .A2(_22580_),
    .B1(_22588_),
    .X(_22589_));
 sky130_fd_sc_hd__buf_1 _28979_ (.A(_22589_),
    .X(_22590_));
 sky130_fd_sc_hd__nand3_4 _28980_ (.A(_22578_),
    .B(_22588_),
    .C(_22580_),
    .Y(_22591_));
 sky130_fd_sc_hd__and2_4 _28981_ (.A(_22590_),
    .B(_22591_),
    .X(_22592_));
 sky130_fd_sc_hd__maj3_4 _28982_ (.A(\decoded_imm_uj[19] ),
    .B(_22561_),
    .C(_22555_),
    .X(_22593_));
 sky130_fd_sc_hd__a211o_4 _28983_ (.A1(_22542_),
    .A2(_22587_),
    .B1(_22592_),
    .C1(_22593_),
    .X(_22594_));
 sky130_fd_sc_hd__nand2_4 _28984_ (.A(_22542_),
    .B(_22587_),
    .Y(_22595_));
 sky130_vsdinv _28985_ (.A(_22593_),
    .Y(_22596_));
 sky130_fd_sc_hd__nand2_4 _28986_ (.A(_22595_),
    .B(_22596_),
    .Y(_22597_));
 sky130_fd_sc_hd__nand2_4 _28987_ (.A(_22597_),
    .B(_22592_),
    .Y(_22598_));
 sky130_fd_sc_hd__a21oi_4 _28988_ (.A1(_22594_),
    .A2(_22598_),
    .B1(_22144_),
    .Y(_22599_));
 sky130_fd_sc_hd__a2111oi_4 _28989_ (.A1(_22478_),
    .A2(_22584_),
    .B1(_22229_),
    .C1(_21975_),
    .D1(_22599_),
    .Y(_22600_));
 sky130_fd_sc_hd__o21ai_4 _28990_ (.A1(_22586_),
    .A2(_22600_),
    .B1(_22427_),
    .Y(_22601_));
 sky130_vsdinv _28991_ (.A(_22582_),
    .Y(_22602_));
 sky130_fd_sc_hd__buf_1 _28992_ (.A(_22371_),
    .X(_22603_));
 sky130_fd_sc_hd__a21oi_4 _28993_ (.A1(_22571_),
    .A2(_22602_),
    .B1(_22603_),
    .Y(_22604_));
 sky130_fd_sc_hd__buf_1 _28994_ (.A(_22374_),
    .X(_22605_));
 sky130_fd_sc_hd__o21ai_4 _28995_ (.A1(_22549_),
    .A2(\reg_next_pc[20] ),
    .B1(_22605_),
    .Y(_22606_));
 sky130_fd_sc_hd__a21oi_4 _28996_ (.A1(_22601_),
    .A2(_22604_),
    .B1(_22606_),
    .Y(_00510_));
 sky130_fd_sc_hd__buf_1 _28997_ (.A(_22433_),
    .X(_22607_));
 sky130_fd_sc_hd__buf_1 _28998_ (.A(_22498_),
    .X(_22608_));
 sky130_fd_sc_hd__or2_4 _28999_ (.A(_22608_),
    .B(\reg_out[21] ),
    .X(_22609_));
 sky130_fd_sc_hd__o21a_4 _29000_ (.A1(_22607_),
    .A2(\alu_out_q[21] ),
    .B1(_22609_),
    .X(_22610_));
 sky130_fd_sc_hd__nand2_4 _29001_ (.A(_22610_),
    .B(_21915_),
    .Y(_22611_));
 sky130_fd_sc_hd__buf_1 _29002_ (.A(_22438_),
    .X(_22612_));
 sky130_fd_sc_hd__nand3_4 _29003_ (.A(_22612_),
    .B(\reg_next_pc[21] ),
    .C(_22526_),
    .Y(_22613_));
 sky130_fd_sc_hd__nand2_4 _29004_ (.A(_22611_),
    .B(_22613_),
    .Y(_22614_));
 sky130_fd_sc_hd__xor2_4 _29005_ (.A(\decoded_imm_uj[21] ),
    .B(_22614_),
    .X(_22615_));
 sky130_fd_sc_hd__a21oi_4 _29006_ (.A1(_22598_),
    .A2(_22590_),
    .B1(_22615_),
    .Y(_22616_));
 sky130_fd_sc_hd__nand3_4 _29007_ (.A(_22598_),
    .B(_22590_),
    .C(_22615_),
    .Y(_22617_));
 sky130_fd_sc_hd__buf_1 _29008_ (.A(_18774_),
    .X(_22618_));
 sky130_fd_sc_hd__buf_1 _29009_ (.A(_22618_),
    .X(_22619_));
 sky130_fd_sc_hd__nand2_4 _29010_ (.A(_22617_),
    .B(_22619_),
    .Y(_22620_));
 sky130_vsdinv _29011_ (.A(_22614_),
    .Y(_22621_));
 sky130_fd_sc_hd__and4_4 _29012_ (.A(_22531_),
    .B(_22529_),
    .C(_22556_),
    .D(_22602_),
    .X(_22622_));
 sky130_fd_sc_hd__xor2_4 _29013_ (.A(_22621_),
    .B(_22622_),
    .X(_22623_));
 sky130_fd_sc_hd__a21oi_4 _29014_ (.A1(_22623_),
    .A2(_22266_),
    .B1(_22067_),
    .Y(_22624_));
 sky130_fd_sc_hd__o21ai_4 _29015_ (.A1(_22616_),
    .A2(_22620_),
    .B1(_22624_),
    .Y(_22625_));
 sky130_fd_sc_hd__nand3_4 _29016_ (.A(_22207_),
    .B(_22208_),
    .C(_22621_),
    .Y(_22626_));
 sky130_vsdinv _29017_ (.A(_22626_),
    .Y(_22627_));
 sky130_fd_sc_hd__a211o_4 _29018_ (.A1(_22623_),
    .A2(_22452_),
    .B1(_22566_),
    .C1(_22627_),
    .X(_22628_));
 sky130_fd_sc_hd__buf_1 _29019_ (.A(_18547_),
    .X(_22629_));
 sky130_fd_sc_hd__a21o_4 _29020_ (.A1(_22625_),
    .A2(_22628_),
    .B1(_22629_),
    .X(_22630_));
 sky130_fd_sc_hd__buf_1 _29021_ (.A(_22614_),
    .X(_22631_));
 sky130_fd_sc_hd__a21oi_4 _29022_ (.A1(_22571_),
    .A2(_22631_),
    .B1(_22603_),
    .Y(_22632_));
 sky130_fd_sc_hd__o21ai_4 _29023_ (.A1(_22549_),
    .A2(\reg_next_pc[21] ),
    .B1(_22605_),
    .Y(_22633_));
 sky130_fd_sc_hd__a21oi_4 _29024_ (.A1(_22630_),
    .A2(_22632_),
    .B1(_22633_),
    .Y(_00511_));
 sky130_fd_sc_hd__buf_1 _29025_ (.A(_22401_),
    .X(_22634_));
 sky130_fd_sc_hd__or2_4 _29026_ (.A(_22608_),
    .B(\reg_out[22] ),
    .X(_22635_));
 sky130_fd_sc_hd__o21a_4 _29027_ (.A1(_22522_),
    .A2(\alu_out_q[22] ),
    .B1(_22635_),
    .X(_22636_));
 sky130_fd_sc_hd__o21a_4 _29028_ (.A1(_22463_),
    .A2(_22636_),
    .B1(_22576_),
    .X(_22637_));
 sky130_fd_sc_hd__o21ai_4 _29029_ (.A1(_22634_),
    .A2(_22637_),
    .B1(\reg_next_pc[22] ),
    .Y(_22638_));
 sky130_fd_sc_hd__buf_1 _29030_ (.A(_22576_),
    .X(_22639_));
 sky130_fd_sc_hd__nand3_4 _29031_ (.A(_22636_),
    .B(_22639_),
    .C(_22579_),
    .Y(_22640_));
 sky130_fd_sc_hd__and2_4 _29032_ (.A(_22638_),
    .B(_22640_),
    .X(_22641_));
 sky130_fd_sc_hd__buf_1 _29033_ (.A(_22641_),
    .X(_22642_));
 sky130_fd_sc_hd__and4_4 _29034_ (.A(_22558_),
    .B(_22556_),
    .C(_22602_),
    .D(_22631_),
    .X(_22643_));
 sky130_fd_sc_hd__xor2_4 _29035_ (.A(_22642_),
    .B(_22643_),
    .X(_22644_));
 sky130_fd_sc_hd__buf_1 _29036_ (.A(_22100_),
    .X(_22645_));
 sky130_fd_sc_hd__buf_1 _29037_ (.A(_22102_),
    .X(_22646_));
 sky130_fd_sc_hd__and3_4 _29038_ (.A(_22638_),
    .B(_22414_),
    .C(_22640_),
    .X(_22647_));
 sky130_fd_sc_hd__a2111oi_4 _29039_ (.A1(_22644_),
    .A2(_22645_),
    .B1(_22646_),
    .C1(_22475_),
    .D1(_22647_),
    .Y(_22648_));
 sky130_vsdinv _29040_ (.A(\decoded_imm_uj[22] ),
    .Y(_22649_));
 sky130_fd_sc_hd__a21o_4 _29041_ (.A1(_22638_),
    .A2(_22640_),
    .B1(_22649_),
    .X(_22650_));
 sky130_fd_sc_hd__buf_1 _29042_ (.A(_22650_),
    .X(_22651_));
 sky130_fd_sc_hd__nand3_4 _29043_ (.A(_22638_),
    .B(_22649_),
    .C(_22640_),
    .Y(_22652_));
 sky130_fd_sc_hd__and2_4 _29044_ (.A(_22651_),
    .B(_22652_),
    .X(_22653_));
 sky130_vsdinv _29045_ (.A(_22653_),
    .Y(_22654_));
 sky130_fd_sc_hd__nand3_4 _29046_ (.A(_22590_),
    .B(_22591_),
    .C(_22615_),
    .Y(_22655_));
 sky130_vsdinv _29047_ (.A(_22655_),
    .Y(_22656_));
 sky130_vsdinv _29048_ (.A(\decoded_imm_uj[21] ),
    .Y(_22657_));
 sky130_fd_sc_hd__maj3_4 _29049_ (.A(_22657_),
    .B(_22589_),
    .C(_22621_),
    .X(_22658_));
 sky130_fd_sc_hd__a21boi_4 _29050_ (.A1(_22597_),
    .A2(_22656_),
    .B1_N(_22658_),
    .Y(_22659_));
 sky130_fd_sc_hd__or2_4 _29051_ (.A(_22654_),
    .B(_22659_),
    .X(_22660_));
 sky130_fd_sc_hd__nand2_4 _29052_ (.A(_22659_),
    .B(_22654_),
    .Y(_22661_));
 sky130_fd_sc_hd__a21oi_4 _29053_ (.A1(_22660_),
    .A2(_22661_),
    .B1(_22144_),
    .Y(_22662_));
 sky130_fd_sc_hd__a2111oi_4 _29054_ (.A1(_22478_),
    .A2(_22644_),
    .B1(_22229_),
    .C1(_21975_),
    .D1(_22662_),
    .Y(_22663_));
 sky130_fd_sc_hd__buf_1 _29055_ (.A(_18485_),
    .X(_22664_));
 sky130_fd_sc_hd__o21ai_4 _29056_ (.A1(_22648_),
    .A2(_22663_),
    .B1(_22664_),
    .Y(_22665_));
 sky130_vsdinv _29057_ (.A(_22642_),
    .Y(_22666_));
 sky130_fd_sc_hd__a21oi_4 _29058_ (.A1(_22571_),
    .A2(_22666_),
    .B1(_22603_),
    .Y(_22667_));
 sky130_fd_sc_hd__buf_1 _29059_ (.A(_22314_),
    .X(_22668_));
 sky130_fd_sc_hd__o21ai_4 _29060_ (.A1(_22668_),
    .A2(\reg_next_pc[22] ),
    .B1(_22605_),
    .Y(_22669_));
 sky130_fd_sc_hd__a21oi_4 _29061_ (.A1(_22665_),
    .A2(_22667_),
    .B1(_22669_),
    .Y(_00512_));
 sky130_fd_sc_hd__buf_1 _29062_ (.A(_22608_),
    .X(_22670_));
 sky130_fd_sc_hd__or2_4 _29063_ (.A(_22670_),
    .B(\reg_out[23] ),
    .X(_22671_));
 sky130_fd_sc_hd__o21a_4 _29064_ (.A1(_22607_),
    .A2(\alu_out_q[23] ),
    .B1(_22671_),
    .X(_22672_));
 sky130_fd_sc_hd__nand2_4 _29065_ (.A(_22672_),
    .B(_21915_),
    .Y(_22673_));
 sky130_fd_sc_hd__buf_1 _29066_ (.A(_22526_),
    .X(_22674_));
 sky130_fd_sc_hd__nand3_4 _29067_ (.A(_22612_),
    .B(\reg_next_pc[23] ),
    .C(_22674_),
    .Y(_22675_));
 sky130_fd_sc_hd__nand2_4 _29068_ (.A(_22673_),
    .B(_22675_),
    .Y(_22676_));
 sky130_vsdinv _29069_ (.A(_22676_),
    .Y(_22677_));
 sky130_fd_sc_hd__and4_4 _29070_ (.A(_22583_),
    .B(_22602_),
    .C(_22631_),
    .D(_22666_),
    .X(_22678_));
 sky130_fd_sc_hd__buf_1 _29071_ (.A(_22678_),
    .X(_22679_));
 sky130_fd_sc_hd__xor2_4 _29072_ (.A(_22677_),
    .B(_22679_),
    .X(_22680_));
 sky130_fd_sc_hd__xor2_4 _29073_ (.A(\decoded_imm_uj[23] ),
    .B(_22676_),
    .X(_22681_));
 sky130_fd_sc_hd__a21oi_4 _29074_ (.A1(_22660_),
    .A2(_22651_),
    .B1(_22681_),
    .Y(_22682_));
 sky130_fd_sc_hd__and3_4 _29075_ (.A(_22660_),
    .B(_22651_),
    .C(_22681_),
    .X(_22683_));
 sky130_fd_sc_hd__nor3_4 _29076_ (.A(_22197_),
    .B(_22682_),
    .C(_22683_),
    .Y(_22684_));
 sky130_fd_sc_hd__a211o_4 _29077_ (.A1(_22183_),
    .A2(_22680_),
    .B1(_22145_),
    .C1(_22684_),
    .X(_22685_));
 sky130_fd_sc_hd__buf_1 _29078_ (.A(_22070_),
    .X(_22686_));
 sky130_fd_sc_hd__nand3_4 _29079_ (.A(_22148_),
    .B(_22149_),
    .C(_22677_),
    .Y(_22687_));
 sky130_vsdinv _29080_ (.A(_22687_),
    .Y(_22688_));
 sky130_fd_sc_hd__a211o_4 _29081_ (.A1(_22680_),
    .A2(_22686_),
    .B1(_22566_),
    .C1(_22688_),
    .X(_22689_));
 sky130_fd_sc_hd__a21o_4 _29082_ (.A1(_22685_),
    .A2(_22689_),
    .B1(_22629_),
    .X(_22690_));
 sky130_fd_sc_hd__buf_1 _29083_ (.A(_22459_),
    .X(_22691_));
 sky130_fd_sc_hd__buf_1 _29084_ (.A(_22676_),
    .X(_22692_));
 sky130_fd_sc_hd__a21oi_4 _29085_ (.A1(_22691_),
    .A2(_22692_),
    .B1(_22603_),
    .Y(_22693_));
 sky130_fd_sc_hd__o21ai_4 _29086_ (.A1(_22668_),
    .A2(\reg_next_pc[23] ),
    .B1(_22605_),
    .Y(_22694_));
 sky130_fd_sc_hd__a21oi_4 _29087_ (.A1(_22690_),
    .A2(_22693_),
    .B1(_22694_),
    .Y(_00513_));
 sky130_fd_sc_hd__buf_1 _29088_ (.A(_22463_),
    .X(_22695_));
 sky130_fd_sc_hd__or2_4 _29089_ (.A(\alu_out_q[24] ),
    .B(_22522_),
    .X(_22696_));
 sky130_fd_sc_hd__o21a_4 _29090_ (.A1(_22608_),
    .A2(\reg_out[24] ),
    .B1(_22696_),
    .X(_22697_));
 sky130_fd_sc_hd__o21a_4 _29091_ (.A1(_22695_),
    .A2(_22697_),
    .B1(_22639_),
    .X(_22698_));
 sky130_fd_sc_hd__o21ai_4 _29092_ (.A1(_22634_),
    .A2(_22698_),
    .B1(\reg_next_pc[24] ),
    .Y(_22699_));
 sky130_fd_sc_hd__nand3_4 _29093_ (.A(_22697_),
    .B(_22639_),
    .C(_22579_),
    .Y(_22700_));
 sky130_fd_sc_hd__and2_4 _29094_ (.A(_22699_),
    .B(_22700_),
    .X(_22701_));
 sky130_fd_sc_hd__buf_1 _29095_ (.A(_22701_),
    .X(_22702_));
 sky130_fd_sc_hd__and4_4 _29096_ (.A(_22622_),
    .B(_22631_),
    .C(_22666_),
    .D(_22692_),
    .X(_22703_));
 sky130_fd_sc_hd__xor2_4 _29097_ (.A(_22702_),
    .B(_22703_),
    .X(_22704_));
 sky130_fd_sc_hd__buf_1 _29098_ (.A(_22105_),
    .X(_22705_));
 sky130_fd_sc_hd__and3_4 _29099_ (.A(_22699_),
    .B(_22033_),
    .C(_22700_),
    .X(_22706_));
 sky130_fd_sc_hd__a2111oi_4 _29100_ (.A1(_22704_),
    .A2(_22645_),
    .B1(_22646_),
    .C1(_22705_),
    .D1(_22706_),
    .Y(_22707_));
 sky130_fd_sc_hd__buf_1 _29101_ (.A(_19135_),
    .X(_22708_));
 sky130_vsdinv _29102_ (.A(\decoded_imm_uj[24] ),
    .Y(_22709_));
 sky130_fd_sc_hd__xor2_4 _29103_ (.A(_22709_),
    .B(_22702_),
    .X(_22710_));
 sky130_fd_sc_hd__nand3_4 _29104_ (.A(_22651_),
    .B(_22652_),
    .C(_22681_),
    .Y(_22711_));
 sky130_vsdinv _29105_ (.A(\decoded_imm_uj[23] ),
    .Y(_22712_));
 sky130_fd_sc_hd__maj3_4 _29106_ (.A(_22712_),
    .B(_22650_),
    .C(_22677_),
    .X(_22713_));
 sky130_fd_sc_hd__o21ai_4 _29107_ (.A1(_22711_),
    .A2(_22659_),
    .B1(_22713_),
    .Y(_22714_));
 sky130_fd_sc_hd__or2_4 _29108_ (.A(_22710_),
    .B(_22714_),
    .X(_22715_));
 sky130_fd_sc_hd__nand2_4 _29109_ (.A(_22714_),
    .B(_22710_),
    .Y(_22716_));
 sky130_fd_sc_hd__a21oi_4 _29110_ (.A1(_22715_),
    .A2(_22716_),
    .B1(_22144_),
    .Y(_22717_));
 sky130_fd_sc_hd__a2111oi_4 _29111_ (.A1(_22478_),
    .A2(_22704_),
    .B1(_22708_),
    .C1(_21975_),
    .D1(_22717_),
    .Y(_22718_));
 sky130_fd_sc_hd__o21ai_4 _29112_ (.A1(_22707_),
    .A2(_22718_),
    .B1(_22664_),
    .Y(_22719_));
 sky130_vsdinv _29113_ (.A(_22702_),
    .Y(_22720_));
 sky130_fd_sc_hd__buf_1 _29114_ (.A(_22720_),
    .X(_22721_));
 sky130_fd_sc_hd__buf_1 _29115_ (.A(_22371_),
    .X(_22722_));
 sky130_fd_sc_hd__a21oi_4 _29116_ (.A1(_22691_),
    .A2(_22721_),
    .B1(_22722_),
    .Y(_22723_));
 sky130_fd_sc_hd__buf_1 _29117_ (.A(_22374_),
    .X(_22724_));
 sky130_fd_sc_hd__o21ai_4 _29118_ (.A1(_22668_),
    .A2(\reg_next_pc[24] ),
    .B1(_22724_),
    .Y(_22725_));
 sky130_fd_sc_hd__a21oi_4 _29119_ (.A1(_22719_),
    .A2(_22723_),
    .B1(_22725_),
    .Y(_00514_));
 sky130_fd_sc_hd__a21oi_4 _29120_ (.A1(_22699_),
    .A2(_22700_),
    .B1(_22709_),
    .Y(_22726_));
 sky130_vsdinv _29121_ (.A(_22726_),
    .Y(_22727_));
 sky130_fd_sc_hd__buf_1 _29122_ (.A(_22670_),
    .X(_22728_));
 sky130_fd_sc_hd__or2_4 _29123_ (.A(\alu_out_q[25] ),
    .B(_22607_),
    .X(_22729_));
 sky130_fd_sc_hd__o21a_4 _29124_ (.A1(_22728_),
    .A2(\reg_out[25] ),
    .B1(_22729_),
    .X(_22730_));
 sky130_fd_sc_hd__nand2_4 _29125_ (.A(_22730_),
    .B(_21916_),
    .Y(_22731_));
 sky130_fd_sc_hd__buf_1 _29126_ (.A(_22612_),
    .X(_22732_));
 sky130_fd_sc_hd__buf_1 _29127_ (.A(_22674_),
    .X(_22733_));
 sky130_fd_sc_hd__nand3_4 _29128_ (.A(_22732_),
    .B(\reg_next_pc[25] ),
    .C(_22733_),
    .Y(_22734_));
 sky130_fd_sc_hd__nand2_4 _29129_ (.A(_22731_),
    .B(_22734_),
    .Y(_22735_));
 sky130_fd_sc_hd__buf_1 _29130_ (.A(_22735_),
    .X(_22736_));
 sky130_fd_sc_hd__xor2_4 _29131_ (.A(\decoded_imm_uj[25] ),
    .B(_22736_),
    .X(_22737_));
 sky130_fd_sc_hd__a21oi_4 _29132_ (.A1(_22716_),
    .A2(_22727_),
    .B1(_22737_),
    .Y(_22738_));
 sky130_vsdinv _29133_ (.A(\decoded_imm_uj[25] ),
    .Y(_22739_));
 sky130_fd_sc_hd__a21oi_4 _29134_ (.A1(_22731_),
    .A2(_22734_),
    .B1(_22739_),
    .Y(_22740_));
 sky130_vsdinv _29135_ (.A(_22740_),
    .Y(_22741_));
 sky130_fd_sc_hd__nand3_4 _29136_ (.A(_22731_),
    .B(_22739_),
    .C(_22734_),
    .Y(_22742_));
 sky130_fd_sc_hd__buf_1 _29137_ (.A(_22742_),
    .X(_22743_));
 sky130_fd_sc_hd__a41o_4 _29138_ (.A1(_22716_),
    .A2(_22727_),
    .A3(_22741_),
    .A4(_22743_),
    .B1(_22260_),
    .X(_22744_));
 sky130_vsdinv _29139_ (.A(_22736_),
    .Y(_22745_));
 sky130_fd_sc_hd__and4_4 _29140_ (.A(_22643_),
    .B(_22666_),
    .C(_22676_),
    .D(_22720_),
    .X(_22746_));
 sky130_fd_sc_hd__xor2_4 _29141_ (.A(_22745_),
    .B(_22746_),
    .X(_22747_));
 sky130_fd_sc_hd__a21oi_4 _29142_ (.A1(_22747_),
    .A2(_22266_),
    .B1(_22067_),
    .Y(_22748_));
 sky130_fd_sc_hd__o21ai_4 _29143_ (.A1(_22738_),
    .A2(_22744_),
    .B1(_22748_),
    .Y(_22749_));
 sky130_fd_sc_hd__nand3_4 _29144_ (.A(_22745_),
    .B(_22269_),
    .C(_22270_),
    .Y(_22750_));
 sky130_vsdinv _29145_ (.A(_22750_),
    .Y(_22751_));
 sky130_fd_sc_hd__a211o_4 _29146_ (.A1(_22747_),
    .A2(_22686_),
    .B1(_22566_),
    .C1(_22751_),
    .X(_22752_));
 sky130_fd_sc_hd__a21o_4 _29147_ (.A1(_22749_),
    .A2(_22752_),
    .B1(_22629_),
    .X(_22753_));
 sky130_fd_sc_hd__a21oi_4 _29148_ (.A1(_22691_),
    .A2(_22736_),
    .B1(_22722_),
    .Y(_22754_));
 sky130_fd_sc_hd__o21ai_4 _29149_ (.A1(_22668_),
    .A2(\reg_next_pc[25] ),
    .B1(_22724_),
    .Y(_22755_));
 sky130_fd_sc_hd__a21oi_4 _29150_ (.A1(_22753_),
    .A2(_22754_),
    .B1(_22755_),
    .Y(_00515_));
 sky130_fd_sc_hd__buf_1 _29151_ (.A(_22607_),
    .X(_22756_));
 sky130_fd_sc_hd__or2_4 _29152_ (.A(_22670_),
    .B(\reg_out[26] ),
    .X(_22757_));
 sky130_fd_sc_hd__o21a_4 _29153_ (.A1(_22756_),
    .A2(\alu_out_q[26] ),
    .B1(_22757_),
    .X(_22758_));
 sky130_fd_sc_hd__nand2_4 _29154_ (.A(_22758_),
    .B(_21916_),
    .Y(_22759_));
 sky130_fd_sc_hd__nand3_4 _29155_ (.A(_22732_),
    .B(\reg_next_pc[26] ),
    .C(_22674_),
    .Y(_22760_));
 sky130_fd_sc_hd__nand2_4 _29156_ (.A(_22759_),
    .B(_22760_),
    .Y(_22761_));
 sky130_fd_sc_hd__buf_1 _29157_ (.A(_22761_),
    .X(_22762_));
 sky130_vsdinv _29158_ (.A(_22762_),
    .Y(_22763_));
 sky130_fd_sc_hd__nand3_4 _29159_ (.A(_22326_),
    .B(_22327_),
    .C(_22763_),
    .Y(_22764_));
 sky130_vsdinv _29160_ (.A(_22764_),
    .Y(_22765_));
 sky130_fd_sc_hd__and4_4 _29161_ (.A(_22703_),
    .B(_22721_),
    .C(_22735_),
    .D(_22761_),
    .X(_22766_));
 sky130_fd_sc_hd__buf_1 _29162_ (.A(_22766_),
    .X(_22767_));
 sky130_vsdinv _29163_ (.A(_22767_),
    .Y(_22768_));
 sky130_fd_sc_hd__a41o_4 _29164_ (.A1(_22679_),
    .A2(_22692_),
    .A3(_22721_),
    .A4(_22736_),
    .B1(_22762_),
    .X(_22769_));
 sky130_fd_sc_hd__a21oi_4 _29165_ (.A1(_22768_),
    .A2(_22769_),
    .B1(_22034_),
    .Y(_22770_));
 sky130_fd_sc_hd__nor3_4 _29166_ (.A(_22035_),
    .B(_22765_),
    .C(_22770_),
    .Y(_22771_));
 sky130_fd_sc_hd__xor2_4 _29167_ (.A(\decoded_imm_uj[26] ),
    .B(_22761_),
    .X(_22772_));
 sky130_fd_sc_hd__nand3_4 _29168_ (.A(_22714_),
    .B(_22710_),
    .C(_22743_),
    .Y(_22773_));
 sky130_vsdinv _29169_ (.A(_22773_),
    .Y(_22774_));
 sky130_fd_sc_hd__a2111o_4 _29170_ (.A1(_22726_),
    .A2(_22743_),
    .B1(_22740_),
    .C1(_22772_),
    .D1(_22774_),
    .X(_22775_));
 sky130_fd_sc_hd__a21oi_4 _29171_ (.A1(_22726_),
    .A2(_22743_),
    .B1(_22740_),
    .Y(_22776_));
 sky130_fd_sc_hd__a21bo_4 _29172_ (.A1(_22773_),
    .A2(_22776_),
    .B1_N(_22772_),
    .X(_22777_));
 sky130_fd_sc_hd__nand3_4 _29173_ (.A(_22775_),
    .B(_22507_),
    .C(_22777_),
    .Y(_22778_));
 sky130_fd_sc_hd__nand3_4 _29174_ (.A(_22768_),
    .B(_21923_),
    .C(_22769_),
    .Y(_22779_));
 sky130_fd_sc_hd__a21oi_4 _29175_ (.A1(_22778_),
    .A2(_22779_),
    .B1(_22425_),
    .Y(_22780_));
 sky130_fd_sc_hd__o21ai_4 _29176_ (.A1(_22771_),
    .A2(_22780_),
    .B1(_22664_),
    .Y(_22781_));
 sky130_fd_sc_hd__a21oi_4 _29177_ (.A1(_22691_),
    .A2(_22762_),
    .B1(_22722_),
    .Y(_22782_));
 sky130_fd_sc_hd__buf_1 _29178_ (.A(_19114_),
    .X(_22783_));
 sky130_fd_sc_hd__buf_1 _29179_ (.A(_22783_),
    .X(_22784_));
 sky130_fd_sc_hd__o21ai_4 _29180_ (.A1(_22784_),
    .A2(\reg_next_pc[26] ),
    .B1(_22724_),
    .Y(_22785_));
 sky130_fd_sc_hd__a21oi_4 _29181_ (.A1(_22781_),
    .A2(_22782_),
    .B1(_22785_),
    .Y(_00516_));
 sky130_fd_sc_hd__or2_4 _29182_ (.A(_22670_),
    .B(\reg_out[27] ),
    .X(_22786_));
 sky130_fd_sc_hd__o21a_4 _29183_ (.A1(_22756_),
    .A2(\alu_out_q[27] ),
    .B1(_22786_),
    .X(_22787_));
 sky130_fd_sc_hd__nand2_4 _29184_ (.A(_22787_),
    .B(_21916_),
    .Y(_22788_));
 sky130_fd_sc_hd__nand3_4 _29185_ (.A(_22612_),
    .B(\reg_next_pc[27] ),
    .C(_22674_),
    .Y(_22789_));
 sky130_fd_sc_hd__nand2_4 _29186_ (.A(_22788_),
    .B(_22789_),
    .Y(_22790_));
 sky130_vsdinv _29187_ (.A(_22790_),
    .Y(_22791_));
 sky130_fd_sc_hd__xor2_4 _29188_ (.A(_22791_),
    .B(_22767_),
    .X(_22792_));
 sky130_vsdinv _29189_ (.A(\decoded_imm_uj[26] ),
    .Y(_22793_));
 sky130_fd_sc_hd__a21oi_4 _29190_ (.A1(_22759_),
    .A2(_22760_),
    .B1(_22793_),
    .Y(_22794_));
 sky130_vsdinv _29191_ (.A(_22794_),
    .Y(_22795_));
 sky130_fd_sc_hd__xor2_4 _29192_ (.A(\decoded_imm_uj[27] ),
    .B(_22790_),
    .X(_22796_));
 sky130_fd_sc_hd__a21oi_4 _29193_ (.A1(_22777_),
    .A2(_22795_),
    .B1(_22796_),
    .Y(_22797_));
 sky130_fd_sc_hd__and3_4 _29194_ (.A(_22777_),
    .B(_22795_),
    .C(_22796_),
    .X(_22798_));
 sky130_fd_sc_hd__nor3_4 _29195_ (.A(_22197_),
    .B(_22797_),
    .C(_22798_),
    .Y(_22799_));
 sky130_fd_sc_hd__a211o_4 _29196_ (.A1(_22122_),
    .A2(_22792_),
    .B1(_22145_),
    .C1(_22799_),
    .X(_22800_));
 sky130_fd_sc_hd__nand3_4 _29197_ (.A(_22148_),
    .B(_22149_),
    .C(_22791_),
    .Y(_22801_));
 sky130_vsdinv _29198_ (.A(_22801_),
    .Y(_22802_));
 sky130_fd_sc_hd__a211o_4 _29199_ (.A1(_22792_),
    .A2(_22686_),
    .B1(_21953_),
    .C1(_22802_),
    .X(_22803_));
 sky130_fd_sc_hd__a21o_4 _29200_ (.A1(_22800_),
    .A2(_22803_),
    .B1(_22629_),
    .X(_22804_));
 sky130_fd_sc_hd__buf_1 _29201_ (.A(_22459_),
    .X(_22805_));
 sky130_fd_sc_hd__buf_1 _29202_ (.A(_22790_),
    .X(_22806_));
 sky130_fd_sc_hd__a21oi_4 _29203_ (.A1(_22805_),
    .A2(_22806_),
    .B1(_22722_),
    .Y(_22807_));
 sky130_fd_sc_hd__o21ai_4 _29204_ (.A1(_22784_),
    .A2(\reg_next_pc[27] ),
    .B1(_22724_),
    .Y(_22808_));
 sky130_fd_sc_hd__a21oi_4 _29205_ (.A1(_22804_),
    .A2(_22807_),
    .B1(_22808_),
    .Y(_00517_));
 sky130_fd_sc_hd__or2_4 _29206_ (.A(_22728_),
    .B(\reg_out[28] ),
    .X(_22809_));
 sky130_fd_sc_hd__o21a_4 _29207_ (.A1(_22756_),
    .A2(\alu_out_q[28] ),
    .B1(_22809_),
    .X(_22810_));
 sky130_fd_sc_hd__buf_1 _29208_ (.A(_22639_),
    .X(_22811_));
 sky130_fd_sc_hd__o21a_4 _29209_ (.A1(_22695_),
    .A2(_22810_),
    .B1(_22811_),
    .X(_22812_));
 sky130_fd_sc_hd__o21ai_4 _29210_ (.A1(_22634_),
    .A2(_22812_),
    .B1(\reg_next_pc[28] ),
    .Y(_22813_));
 sky130_fd_sc_hd__buf_1 _29211_ (.A(_22579_),
    .X(_22814_));
 sky130_fd_sc_hd__nand3_4 _29212_ (.A(_22810_),
    .B(_22811_),
    .C(_22814_),
    .Y(_22815_));
 sky130_fd_sc_hd__and2_4 _29213_ (.A(_22813_),
    .B(_22815_),
    .X(_22816_));
 sky130_fd_sc_hd__buf_1 _29214_ (.A(_22816_),
    .X(_22817_));
 sky130_fd_sc_hd__and4_4 _29215_ (.A(_22746_),
    .B(_22735_),
    .C(_22761_),
    .D(_22806_),
    .X(_22818_));
 sky130_fd_sc_hd__buf_1 _29216_ (.A(_22818_),
    .X(_22819_));
 sky130_fd_sc_hd__xor2_4 _29217_ (.A(_22817_),
    .B(_22819_),
    .X(_22820_));
 sky130_fd_sc_hd__and3_4 _29218_ (.A(_22813_),
    .B(_22033_),
    .C(_22815_),
    .X(_22821_));
 sky130_fd_sc_hd__a2111oi_4 _29219_ (.A1(_22820_),
    .A2(_22645_),
    .B1(_22646_),
    .C1(_22705_),
    .D1(_22821_),
    .Y(_22822_));
 sky130_vsdinv _29220_ (.A(\decoded_imm_uj[28] ),
    .Y(_22823_));
 sky130_fd_sc_hd__a21oi_4 _29221_ (.A1(_22813_),
    .A2(_22815_),
    .B1(_22823_),
    .Y(_22824_));
 sky130_fd_sc_hd__and3_4 _29222_ (.A(_22813_),
    .B(_22823_),
    .C(_22815_),
    .X(_22825_));
 sky130_fd_sc_hd__nor2_4 _29223_ (.A(_22824_),
    .B(_22825_),
    .Y(_22826_));
 sky130_fd_sc_hd__and4_4 _29224_ (.A(_22772_),
    .B(_22796_),
    .C(_22741_),
    .D(_22742_),
    .X(_22827_));
 sky130_fd_sc_hd__nand3_4 _29225_ (.A(_22714_),
    .B(_22710_),
    .C(_22827_),
    .Y(_22828_));
 sky130_fd_sc_hd__nand2_4 _29226_ (.A(_22772_),
    .B(_22796_),
    .Y(_22829_));
 sky130_vsdinv _29227_ (.A(\decoded_imm_uj[27] ),
    .Y(_22830_));
 sky130_fd_sc_hd__maj3_4 _29228_ (.A(_22830_),
    .B(_22795_),
    .C(_22791_),
    .X(_22831_));
 sky130_fd_sc_hd__o21a_4 _29229_ (.A1(_22829_),
    .A2(_22776_),
    .B1(_22831_),
    .X(_22832_));
 sky130_fd_sc_hd__nand2_4 _29230_ (.A(_22828_),
    .B(_22832_),
    .Y(_22833_));
 sky130_fd_sc_hd__xor2_4 _29231_ (.A(_22826_),
    .B(_22833_),
    .X(_22834_));
 sky130_fd_sc_hd__a21oi_4 _29232_ (.A1(_22820_),
    .A2(_22064_),
    .B1(_22308_),
    .Y(_22835_));
 sky130_fd_sc_hd__o21a_4 _29233_ (.A1(_22112_),
    .A2(_22834_),
    .B1(_22835_),
    .X(_22836_));
 sky130_fd_sc_hd__o21ai_4 _29234_ (.A1(_22822_),
    .A2(_22836_),
    .B1(_22664_),
    .Y(_22837_));
 sky130_vsdinv _29235_ (.A(_22817_),
    .Y(_22838_));
 sky130_fd_sc_hd__buf_1 _29236_ (.A(_19091_),
    .X(_22839_));
 sky130_fd_sc_hd__a21oi_4 _29237_ (.A1(_22805_),
    .A2(_22838_),
    .B1(_22839_),
    .Y(_22840_));
 sky130_fd_sc_hd__buf_1 _29238_ (.A(_18536_),
    .X(_22841_));
 sky130_fd_sc_hd__buf_1 _29239_ (.A(_22841_),
    .X(_22842_));
 sky130_fd_sc_hd__o21ai_4 _29240_ (.A1(_22784_),
    .A2(\reg_next_pc[28] ),
    .B1(_22842_),
    .Y(_22843_));
 sky130_fd_sc_hd__a21oi_4 _29241_ (.A1(_22837_),
    .A2(_22840_),
    .B1(_22843_),
    .Y(_00518_));
 sky130_fd_sc_hd__buf_1 _29242_ (.A(_22756_),
    .X(_22844_));
 sky130_fd_sc_hd__buf_1 _29243_ (.A(_22728_),
    .X(_22845_));
 sky130_fd_sc_hd__or2_4 _29244_ (.A(_22845_),
    .B(\reg_out[29] ),
    .X(_22846_));
 sky130_fd_sc_hd__o21a_4 _29245_ (.A1(_22844_),
    .A2(\alu_out_q[29] ),
    .B1(_22846_),
    .X(_22847_));
 sky130_fd_sc_hd__nand2_4 _29246_ (.A(_22847_),
    .B(_21917_),
    .Y(_22848_));
 sky130_fd_sc_hd__nand3_4 _29247_ (.A(_22732_),
    .B(\reg_next_pc[29] ),
    .C(_22733_),
    .Y(_22849_));
 sky130_fd_sc_hd__nand2_4 _29248_ (.A(_22848_),
    .B(_22849_),
    .Y(_22850_));
 sky130_fd_sc_hd__buf_1 _29249_ (.A(_22850_),
    .X(_22851_));
 sky130_vsdinv _29250_ (.A(_22851_),
    .Y(_22852_));
 sky130_fd_sc_hd__and4_4 _29251_ (.A(_22679_),
    .B(_22692_),
    .C(_22721_),
    .D(_22735_),
    .X(_22853_));
 sky130_fd_sc_hd__and4_4 _29252_ (.A(_22853_),
    .B(_22762_),
    .C(_22806_),
    .D(_22838_),
    .X(_22854_));
 sky130_fd_sc_hd__xor2_4 _29253_ (.A(_22852_),
    .B(_22854_),
    .X(_22855_));
 sky130_fd_sc_hd__nand3_4 _29254_ (.A(_22075_),
    .B(_22078_),
    .C(_22852_),
    .Y(_22856_));
 sky130_vsdinv _29255_ (.A(_22856_),
    .Y(_22857_));
 sky130_fd_sc_hd__a2111oi_4 _29256_ (.A1(_22855_),
    .A2(_22645_),
    .B1(_22646_),
    .C1(_22705_),
    .D1(_22857_),
    .Y(_22858_));
 sky130_fd_sc_hd__nand2_4 _29257_ (.A(_22850_),
    .B(\decoded_imm_uj[29] ),
    .Y(_22859_));
 sky130_vsdinv _29258_ (.A(\decoded_imm_uj[29] ),
    .Y(_22860_));
 sky130_fd_sc_hd__nand3_4 _29259_ (.A(_22848_),
    .B(_22860_),
    .C(_22849_),
    .Y(_22861_));
 sky130_fd_sc_hd__and2_4 _29260_ (.A(_22859_),
    .B(_22861_),
    .X(_22862_));
 sky130_vsdinv _29261_ (.A(_22825_),
    .Y(_22863_));
 sky130_fd_sc_hd__a21oi_4 _29262_ (.A1(_22833_),
    .A2(_22863_),
    .B1(_22824_),
    .Y(_22864_));
 sky130_fd_sc_hd__xor2_4 _29263_ (.A(_22862_),
    .B(_22864_),
    .X(_22865_));
 sky130_fd_sc_hd__a21o_4 _29264_ (.A1(_22855_),
    .A2(_22111_),
    .B1(_22195_),
    .X(_22866_));
 sky130_fd_sc_hd__a21oi_4 _29265_ (.A1(_22865_),
    .A2(_22544_),
    .B1(_22866_),
    .Y(_22867_));
 sky130_fd_sc_hd__o21ai_4 _29266_ (.A1(_22858_),
    .A2(_22867_),
    .B1(_21990_),
    .Y(_22868_));
 sky130_fd_sc_hd__a21oi_4 _29267_ (.A1(_22805_),
    .A2(_22851_),
    .B1(_22839_),
    .Y(_22869_));
 sky130_fd_sc_hd__o21ai_4 _29268_ (.A1(_22784_),
    .A2(\reg_next_pc[29] ),
    .B1(_22842_),
    .Y(_22870_));
 sky130_fd_sc_hd__a21oi_4 _29269_ (.A1(_22868_),
    .A2(_22869_),
    .B1(_22870_),
    .Y(_00519_));
 sky130_fd_sc_hd__or2_4 _29270_ (.A(_22728_),
    .B(\reg_out[30] ),
    .X(_22871_));
 sky130_fd_sc_hd__o21a_4 _29271_ (.A1(_22844_),
    .A2(\alu_out_q[30] ),
    .B1(_22871_),
    .X(_22872_));
 sky130_fd_sc_hd__o21a_4 _29272_ (.A1(_22695_),
    .A2(_22872_),
    .B1(_22811_),
    .X(_22873_));
 sky130_fd_sc_hd__o21ai_4 _29273_ (.A1(_22634_),
    .A2(_22873_),
    .B1(\reg_next_pc[30] ),
    .Y(_22874_));
 sky130_fd_sc_hd__buf_1 _29274_ (.A(_22811_),
    .X(_22875_));
 sky130_fd_sc_hd__nand3_4 _29275_ (.A(_22872_),
    .B(_22875_),
    .C(_22814_),
    .Y(_22876_));
 sky130_fd_sc_hd__and3_4 _29276_ (.A(_22874_),
    .B(_22107_),
    .C(_22876_),
    .X(_22877_));
 sky130_fd_sc_hd__nand4_4 _29277_ (.A(_22767_),
    .B(_22806_),
    .C(_22838_),
    .D(_22851_),
    .Y(_22878_));
 sky130_fd_sc_hd__and2_4 _29278_ (.A(_22874_),
    .B(_22876_),
    .X(_22879_));
 sky130_fd_sc_hd__nand2_4 _29279_ (.A(_22878_),
    .B(_22879_),
    .Y(_22880_));
 sky130_vsdinv _29280_ (.A(_22879_),
    .Y(_22881_));
 sky130_fd_sc_hd__nand4_4 _29281_ (.A(_22819_),
    .B(_22838_),
    .C(_22851_),
    .D(_22881_),
    .Y(_22882_));
 sky130_fd_sc_hd__a21oi_4 _29282_ (.A1(_22880_),
    .A2(_22882_),
    .B1(_22034_),
    .Y(_22883_));
 sky130_fd_sc_hd__nor3_4 _29283_ (.A(_22035_),
    .B(_22877_),
    .C(_22883_),
    .Y(_22884_));
 sky130_vsdinv _29284_ (.A(\decoded_imm_uj[30] ),
    .Y(_22885_));
 sky130_fd_sc_hd__a21oi_4 _29285_ (.A1(_22874_),
    .A2(_22876_),
    .B1(_22885_),
    .Y(_22886_));
 sky130_fd_sc_hd__and3_4 _29286_ (.A(_22874_),
    .B(_22885_),
    .C(_22876_),
    .X(_22887_));
 sky130_fd_sc_hd__nor2_4 _29287_ (.A(_22886_),
    .B(_22887_),
    .Y(_22888_));
 sky130_vsdinv _29288_ (.A(_22861_),
    .Y(_22889_));
 sky130_fd_sc_hd__o21ai_4 _29289_ (.A1(_22889_),
    .A2(_22864_),
    .B1(_22859_),
    .Y(_22890_));
 sky130_fd_sc_hd__o21a_4 _29290_ (.A1(_22888_),
    .A2(_22890_),
    .B1(_22057_),
    .X(_22891_));
 sky130_fd_sc_hd__nand2_4 _29291_ (.A(_22890_),
    .B(_22888_),
    .Y(_22892_));
 sky130_fd_sc_hd__nand2_4 _29292_ (.A(_22891_),
    .B(_22892_),
    .Y(_22893_));
 sky130_fd_sc_hd__nand3_4 _29293_ (.A(_22880_),
    .B(_21923_),
    .C(_22882_),
    .Y(_22894_));
 sky130_fd_sc_hd__a21oi_4 _29294_ (.A1(_22893_),
    .A2(_22894_),
    .B1(_22425_),
    .Y(_22895_));
 sky130_fd_sc_hd__o21ai_4 _29295_ (.A1(_22884_),
    .A2(_22895_),
    .B1(_21990_),
    .Y(_22896_));
 sky130_fd_sc_hd__a21oi_4 _29296_ (.A1(_22805_),
    .A2(_22881_),
    .B1(_22839_),
    .Y(_22897_));
 sky130_fd_sc_hd__buf_1 _29297_ (.A(_22783_),
    .X(_22898_));
 sky130_fd_sc_hd__o21ai_4 _29298_ (.A1(_22898_),
    .A2(\reg_next_pc[30] ),
    .B1(_22842_),
    .Y(_22899_));
 sky130_fd_sc_hd__a21oi_4 _29299_ (.A1(_22896_),
    .A2(_22897_),
    .B1(_22899_),
    .Y(_00521_));
 sky130_vsdinv _29300_ (.A(_22886_),
    .Y(_22900_));
 sky130_fd_sc_hd__or2_4 _29301_ (.A(_22845_),
    .B(\reg_out[31] ),
    .X(_22901_));
 sky130_fd_sc_hd__o21a_4 _29302_ (.A1(_22844_),
    .A2(\alu_out_q[31] ),
    .B1(_22901_),
    .X(_22902_));
 sky130_fd_sc_hd__nand2_4 _29303_ (.A(_22902_),
    .B(_21917_),
    .Y(_22903_));
 sky130_fd_sc_hd__nand3_4 _29304_ (.A(_22732_),
    .B(\reg_next_pc[31] ),
    .C(_22733_),
    .Y(_22904_));
 sky130_fd_sc_hd__nand2_4 _29305_ (.A(_22903_),
    .B(_22904_),
    .Y(_22905_));
 sky130_fd_sc_hd__xor2_4 _29306_ (.A(\decoded_imm_uj[31] ),
    .B(_22905_),
    .X(_22906_));
 sky130_fd_sc_hd__a21oi_4 _29307_ (.A1(_22892_),
    .A2(_22900_),
    .B1(_22906_),
    .Y(_22907_));
 sky130_fd_sc_hd__nand3_4 _29308_ (.A(_22892_),
    .B(_22900_),
    .C(_22906_),
    .Y(_22908_));
 sky130_fd_sc_hd__nand2_4 _29309_ (.A(_22908_),
    .B(_21949_),
    .Y(_22909_));
 sky130_fd_sc_hd__xor2_4 _29310_ (.A(_22905_),
    .B(_22882_),
    .X(_22910_));
 sky130_fd_sc_hd__a21oi_4 _29311_ (.A1(_22910_),
    .A2(_22064_),
    .B1(_22308_),
    .Y(_22911_));
 sky130_fd_sc_hd__o21ai_4 _29312_ (.A1(_22907_),
    .A2(_22909_),
    .B1(_22911_),
    .Y(_22912_));
 sky130_vsdinv _29313_ (.A(_22905_),
    .Y(_22913_));
 sky130_fd_sc_hd__nand3_4 _29314_ (.A(_22148_),
    .B(_22149_),
    .C(_22913_),
    .Y(_22914_));
 sky130_vsdinv _29315_ (.A(_22914_),
    .Y(_22915_));
 sky130_fd_sc_hd__a211o_4 _29316_ (.A1(_22910_),
    .A2(_22686_),
    .B1(_21953_),
    .C1(_22915_),
    .X(_22916_));
 sky130_fd_sc_hd__nand2_4 _29317_ (.A(_22912_),
    .B(_22916_),
    .Y(_22917_));
 sky130_fd_sc_hd__nand2_4 _29318_ (.A(_22917_),
    .B(_22125_),
    .Y(_22918_));
 sky130_fd_sc_hd__a21oi_4 _29319_ (.A1(_22084_),
    .A2(_22905_),
    .B1(_22839_),
    .Y(_22919_));
 sky130_fd_sc_hd__o21ai_4 _29320_ (.A1(_22898_),
    .A2(\reg_next_pc[31] ),
    .B1(_22842_),
    .Y(_22920_));
 sky130_fd_sc_hd__a21oi_4 _29321_ (.A1(_22918_),
    .A2(_22919_),
    .B1(_22920_),
    .Y(_00522_));
 sky130_fd_sc_hd__buf_1 _29322_ (.A(_22841_),
    .X(_22921_));
 sky130_fd_sc_hd__o21ai_4 _29323_ (.A1(_22898_),
    .A2(_21361_),
    .B1(_22921_),
    .Y(_22922_));
 sky130_fd_sc_hd__a21oi_4 _29324_ (.A1(_21920_),
    .A2(_19123_),
    .B1(_22922_),
    .Y(_00594_));
 sky130_fd_sc_hd__buf_1 _29325_ (.A(_18850_),
    .X(_22923_));
 sky130_fd_sc_hd__buf_1 _29326_ (.A(_22923_),
    .X(_22924_));
 sky130_fd_sc_hd__buf_1 _29327_ (.A(_18850_),
    .X(_22925_));
 sky130_fd_sc_hd__buf_1 _29328_ (.A(_22925_),
    .X(_22926_));
 sky130_fd_sc_hd__nor2_4 _29329_ (.A(_22926_),
    .B(_18304_),
    .Y(_22927_));
 sky130_fd_sc_hd__a211o_4 _29330_ (.A1(_21955_),
    .A2(_22924_),
    .B1(_18894_),
    .C1(_22927_),
    .X(_22928_));
 sky130_vsdinv _29331_ (.A(_22928_),
    .Y(_00605_));
 sky130_fd_sc_hd__buf_1 _29332_ (.A(_18234_),
    .X(_22929_));
 sky130_fd_sc_hd__o21a_4 _29333_ (.A1(_22924_),
    .A2(_21404_),
    .B1(_22929_),
    .X(_22930_));
 sky130_fd_sc_hd__o21a_4 _29334_ (.A1(_19082_),
    .A2(_21972_),
    .B1(_22930_),
    .X(_00616_));
 sky130_fd_sc_hd__nor2_4 _29335_ (.A(_22926_),
    .B(_21418_),
    .Y(_22931_));
 sky130_fd_sc_hd__a211o_4 _29336_ (.A1(_22062_),
    .A2(_22924_),
    .B1(_18894_),
    .C1(_22931_),
    .X(_22932_));
 sky130_vsdinv _29337_ (.A(_22932_),
    .Y(_00619_));
 sky130_fd_sc_hd__o21ai_4 _29338_ (.A1(_22898_),
    .A2(_21441_),
    .B1(_22921_),
    .Y(_22933_));
 sky130_fd_sc_hd__a21oi_4 _29339_ (.A1(_22095_),
    .A2(_19123_),
    .B1(_22933_),
    .Y(_00620_));
 sky130_fd_sc_hd__buf_1 _29340_ (.A(_18574_),
    .X(_22934_));
 sky130_fd_sc_hd__nor2_4 _29341_ (.A(_22926_),
    .B(_21458_),
    .Y(_22935_));
 sky130_fd_sc_hd__a211o_4 _29342_ (.A1(_22142_),
    .A2(_22924_),
    .B1(_22934_),
    .C1(_22935_),
    .X(_22936_));
 sky130_vsdinv _29343_ (.A(_22936_),
    .Y(_00621_));
 sky130_fd_sc_hd__buf_1 _29344_ (.A(_18851_),
    .X(_22937_));
 sky130_fd_sc_hd__nor2_4 _29345_ (.A(_22926_),
    .B(_21476_),
    .Y(_22938_));
 sky130_fd_sc_hd__a211o_4 _29346_ (.A1(_22164_),
    .A2(_22937_),
    .B1(_22934_),
    .C1(_22938_),
    .X(_22939_));
 sky130_vsdinv _29347_ (.A(_22939_),
    .Y(_00622_));
 sky130_fd_sc_hd__buf_1 _29348_ (.A(_22925_),
    .X(_22940_));
 sky130_fd_sc_hd__nor2_4 _29349_ (.A(_22940_),
    .B(_21490_),
    .Y(_22941_));
 sky130_fd_sc_hd__a211o_4 _29350_ (.A1(_22192_),
    .A2(_22937_),
    .B1(_22934_),
    .C1(_22941_),
    .X(_22942_));
 sky130_vsdinv _29351_ (.A(_22942_),
    .Y(_00623_));
 sky130_fd_sc_hd__buf_1 _29352_ (.A(_22783_),
    .X(_22943_));
 sky130_fd_sc_hd__o21ai_4 _29353_ (.A1(_22943_),
    .A2(_21523_),
    .B1(_22921_),
    .Y(_22944_));
 sky130_fd_sc_hd__a21oi_4 _29354_ (.A1(_22224_),
    .A2(_19123_),
    .B1(_22944_),
    .Y(_00624_));
 sky130_fd_sc_hd__nor2_4 _29355_ (.A(_22940_),
    .B(_21541_),
    .Y(_22945_));
 sky130_fd_sc_hd__a211o_4 _29356_ (.A1(_22263_),
    .A2(_22937_),
    .B1(_22934_),
    .C1(_22945_),
    .X(_22946_));
 sky130_vsdinv _29357_ (.A(_22946_),
    .Y(_00625_));
 sky130_fd_sc_hd__buf_1 _29358_ (.A(_18574_),
    .X(_22947_));
 sky130_fd_sc_hd__nor2_4 _29359_ (.A(_22940_),
    .B(_21559_),
    .Y(_22948_));
 sky130_fd_sc_hd__a211o_4 _29360_ (.A1(_22287_),
    .A2(_22937_),
    .B1(_22947_),
    .C1(_22948_),
    .X(_22949_));
 sky130_vsdinv _29361_ (.A(_22949_),
    .Y(_00595_));
 sky130_fd_sc_hd__buf_1 _29362_ (.A(_22923_),
    .X(_22950_));
 sky130_fd_sc_hd__nor2_4 _29363_ (.A(_22940_),
    .B(_21574_),
    .Y(_22951_));
 sky130_fd_sc_hd__a211o_4 _29364_ (.A1(_22329_),
    .A2(_22950_),
    .B1(_22947_),
    .C1(_22951_),
    .X(_22952_));
 sky130_vsdinv _29365_ (.A(_22952_),
    .Y(_00596_));
 sky130_fd_sc_hd__buf_1 _29366_ (.A(_19122_),
    .X(_22953_));
 sky130_fd_sc_hd__o21ai_4 _29367_ (.A1(_22943_),
    .A2(_21587_),
    .B1(_22921_),
    .Y(_22954_));
 sky130_fd_sc_hd__a21oi_4 _29368_ (.A1(_22353_),
    .A2(_22953_),
    .B1(_22954_),
    .Y(_00597_));
 sky130_fd_sc_hd__buf_1 _29369_ (.A(_22925_),
    .X(_22955_));
 sky130_fd_sc_hd__nor2_4 _29370_ (.A(_22955_),
    .B(_21617_),
    .Y(_22956_));
 sky130_fd_sc_hd__a211o_4 _29371_ (.A1(_22385_),
    .A2(_22950_),
    .B1(_22947_),
    .C1(_22956_),
    .X(_22957_));
 sky130_vsdinv _29372_ (.A(_22957_),
    .Y(_00598_));
 sky130_fd_sc_hd__buf_1 _29373_ (.A(_22841_),
    .X(_22958_));
 sky130_fd_sc_hd__o21ai_4 _29374_ (.A1(_22943_),
    .A2(_21635_),
    .B1(_22958_),
    .Y(_22959_));
 sky130_fd_sc_hd__a21oi_4 _29375_ (.A1(_22409_),
    .A2(_22953_),
    .B1(_22959_),
    .Y(_00599_));
 sky130_fd_sc_hd__nor2_4 _29376_ (.A(_22955_),
    .B(_21650_),
    .Y(_22960_));
 sky130_fd_sc_hd__a211o_4 _29377_ (.A1(_22454_),
    .A2(_22950_),
    .B1(_22947_),
    .C1(_22960_),
    .X(_22961_));
 sky130_vsdinv _29378_ (.A(_22961_),
    .Y(_00600_));
 sky130_fd_sc_hd__o21ai_4 _29379_ (.A1(_22943_),
    .A2(_21665_),
    .B1(_22958_),
    .Y(_22962_));
 sky130_fd_sc_hd__a21oi_4 _29380_ (.A1(_22472_),
    .A2(_22953_),
    .B1(_22962_),
    .Y(_00601_));
 sky130_fd_sc_hd__buf_1 _29381_ (.A(_18284_),
    .X(_22963_));
 sky130_fd_sc_hd__nor2_4 _29382_ (.A(_22955_),
    .B(_21674_),
    .Y(_22964_));
 sky130_fd_sc_hd__a211o_4 _29383_ (.A1(_22511_),
    .A2(_22950_),
    .B1(_22963_),
    .C1(_22964_),
    .X(_22965_));
 sky130_vsdinv _29384_ (.A(_22965_),
    .Y(_00602_));
 sky130_fd_sc_hd__buf_1 _29385_ (.A(_22923_),
    .X(_22966_));
 sky130_fd_sc_hd__nor2_4 _29386_ (.A(_22955_),
    .B(_21701_),
    .Y(_22967_));
 sky130_fd_sc_hd__a211o_4 _29387_ (.A1(_22530_),
    .A2(_22966_),
    .B1(_22963_),
    .C1(_22967_),
    .X(_22968_));
 sky130_vsdinv _29388_ (.A(_22968_),
    .Y(_00603_));
 sky130_fd_sc_hd__buf_1 _29389_ (.A(_22925_),
    .X(_22969_));
 sky130_fd_sc_hd__nor2_4 _29390_ (.A(_22969_),
    .B(_21717_),
    .Y(_22970_));
 sky130_fd_sc_hd__a211o_4 _29391_ (.A1(_22557_),
    .A2(_22966_),
    .B1(_22963_),
    .C1(_22970_),
    .X(_22971_));
 sky130_vsdinv _29392_ (.A(_22971_),
    .Y(_00604_));
 sky130_fd_sc_hd__buf_1 _29393_ (.A(_22783_),
    .X(_22972_));
 sky130_fd_sc_hd__o21ai_4 _29394_ (.A1(_22972_),
    .A2(_21735_),
    .B1(_22958_),
    .Y(_22973_));
 sky130_fd_sc_hd__a21oi_4 _29395_ (.A1(_22582_),
    .A2(_22953_),
    .B1(_22973_),
    .Y(_00606_));
 sky130_fd_sc_hd__nor2_4 _29396_ (.A(_22969_),
    .B(_21743_),
    .Y(_22974_));
 sky130_fd_sc_hd__a211o_4 _29397_ (.A1(_22621_),
    .A2(_22966_),
    .B1(_22963_),
    .C1(_22974_),
    .X(_22975_));
 sky130_vsdinv _29398_ (.A(_22975_),
    .Y(_00607_));
 sky130_fd_sc_hd__buf_1 _29399_ (.A(_19122_),
    .X(_22976_));
 sky130_fd_sc_hd__o21ai_4 _29400_ (.A1(_22972_),
    .A2(_21762_),
    .B1(_22958_),
    .Y(_22977_));
 sky130_fd_sc_hd__a21oi_4 _29401_ (.A1(_22642_),
    .A2(_22976_),
    .B1(_22977_),
    .Y(_00608_));
 sky130_fd_sc_hd__buf_1 _29402_ (.A(_18284_),
    .X(_22978_));
 sky130_fd_sc_hd__nor2_4 _29403_ (.A(_22969_),
    .B(_21772_),
    .Y(_22979_));
 sky130_fd_sc_hd__a211o_4 _29404_ (.A1(_22677_),
    .A2(_22966_),
    .B1(_22978_),
    .C1(_22979_),
    .X(_22980_));
 sky130_vsdinv _29405_ (.A(_22980_),
    .Y(_00609_));
 sky130_fd_sc_hd__buf_1 _29406_ (.A(_22841_),
    .X(_22981_));
 sky130_fd_sc_hd__o21ai_4 _29407_ (.A1(_22972_),
    .A2(_21788_),
    .B1(_22981_),
    .Y(_22982_));
 sky130_fd_sc_hd__a21oi_4 _29408_ (.A1(_22702_),
    .A2(_22976_),
    .B1(_22982_),
    .Y(_00610_));
 sky130_fd_sc_hd__buf_1 _29409_ (.A(_22923_),
    .X(_22983_));
 sky130_fd_sc_hd__nor2_4 _29410_ (.A(_22969_),
    .B(_21796_),
    .Y(_22984_));
 sky130_fd_sc_hd__a211o_4 _29411_ (.A1(_22745_),
    .A2(_22983_),
    .B1(_22978_),
    .C1(_22984_),
    .X(_22985_));
 sky130_vsdinv _29412_ (.A(_22985_),
    .Y(_00611_));
 sky130_fd_sc_hd__buf_1 _29413_ (.A(_19100_),
    .X(_22986_));
 sky130_fd_sc_hd__nor2_4 _29414_ (.A(_22986_),
    .B(_21817_),
    .Y(_22987_));
 sky130_fd_sc_hd__a211o_4 _29415_ (.A1(_22763_),
    .A2(_22983_),
    .B1(_22978_),
    .C1(_22987_),
    .X(_22988_));
 sky130_vsdinv _29416_ (.A(_22988_),
    .Y(_00612_));
 sky130_fd_sc_hd__nor2_4 _29417_ (.A(_22986_),
    .B(_21829_),
    .Y(_22989_));
 sky130_fd_sc_hd__a211o_4 _29418_ (.A1(_22791_),
    .A2(_22983_),
    .B1(_22978_),
    .C1(_22989_),
    .X(_22990_));
 sky130_vsdinv _29419_ (.A(_22990_),
    .Y(_00613_));
 sky130_fd_sc_hd__o21ai_4 _29420_ (.A1(_22972_),
    .A2(_21850_),
    .B1(_22981_),
    .Y(_22991_));
 sky130_fd_sc_hd__a21oi_4 _29421_ (.A1(_22817_),
    .A2(_22976_),
    .B1(_22991_),
    .Y(_00614_));
 sky130_fd_sc_hd__buf_1 _29422_ (.A(_18284_),
    .X(_22992_));
 sky130_fd_sc_hd__nor2_4 _29423_ (.A(_22986_),
    .B(_21865_),
    .Y(_22993_));
 sky130_fd_sc_hd__a211o_4 _29424_ (.A1(_22852_),
    .A2(_22983_),
    .B1(_22992_),
    .C1(_22993_),
    .X(_22994_));
 sky130_vsdinv _29425_ (.A(_22994_),
    .Y(_00615_));
 sky130_fd_sc_hd__o21ai_4 _29426_ (.A1(_19102_),
    .A2(_21887_),
    .B1(_22981_),
    .Y(_22995_));
 sky130_fd_sc_hd__a21oi_4 _29427_ (.A1(_22879_),
    .A2(_22976_),
    .B1(_22995_),
    .Y(_00617_));
 sky130_fd_sc_hd__buf_1 _29428_ (.A(_19114_),
    .X(_22996_));
 sky130_fd_sc_hd__nor2_4 _29429_ (.A(_22986_),
    .B(_21900_),
    .Y(_22997_));
 sky130_fd_sc_hd__a211o_4 _29430_ (.A1(_22913_),
    .A2(_22996_),
    .B1(_22992_),
    .C1(_22997_),
    .X(_22998_));
 sky130_vsdinv _29431_ (.A(_22998_),
    .Y(_00618_));
 sky130_fd_sc_hd__buf_1 _29432_ (.A(\count_instr[0] ),
    .X(_22999_));
 sky130_vsdinv _29433_ (.A(_22999_),
    .Y(_23000_));
 sky130_fd_sc_hd__nor3_4 _29434_ (.A(_19133_),
    .B(_18404_),
    .C(_19137_),
    .Y(_23001_));
 sky130_vsdinv _29435_ (.A(_23001_),
    .Y(_23002_));
 sky130_fd_sc_hd__buf_1 _29436_ (.A(_23002_),
    .X(_23003_));
 sky130_fd_sc_hd__buf_1 _29437_ (.A(_22999_),
    .X(_23004_));
 sky130_fd_sc_hd__buf_1 _29438_ (.A(_23001_),
    .X(_23005_));
 sky130_fd_sc_hd__buf_1 _29439_ (.A(_23005_),
    .X(_23006_));
 sky130_fd_sc_hd__buf_1 _29440_ (.A(_18506_),
    .X(_23007_));
 sky130_fd_sc_hd__o21a_4 _29441_ (.A1(_23004_),
    .A2(_23006_),
    .B1(_23007_),
    .X(_23008_));
 sky130_fd_sc_hd__o21ai_4 _29442_ (.A1(_23000_),
    .A2(_23003_),
    .B1(_23008_),
    .Y(_23009_));
 sky130_vsdinv _29443_ (.A(_23009_),
    .Y(_00068_));
 sky130_fd_sc_hd__buf_1 _29444_ (.A(\count_instr[1] ),
    .X(_23010_));
 sky130_fd_sc_hd__buf_1 _29445_ (.A(_19135_),
    .X(_23011_));
 sky130_fd_sc_hd__buf_1 _29446_ (.A(_19138_),
    .X(_23012_));
 sky130_fd_sc_hd__nor4_4 _29447_ (.A(_23011_),
    .B(_23000_),
    .C(_21926_),
    .D(_23012_),
    .Y(_23013_));
 sky130_fd_sc_hd__o21a_4 _29448_ (.A1(_23010_),
    .A2(_23013_),
    .B1(_19012_),
    .X(_23014_));
 sky130_fd_sc_hd__and4_4 _29449_ (.A(_18465_),
    .B(_18849_),
    .C(_18405_),
    .D(_18468_),
    .X(_23015_));
 sky130_fd_sc_hd__buf_1 _29450_ (.A(_23015_),
    .X(_23016_));
 sky130_fd_sc_hd__buf_1 _29451_ (.A(_18542_),
    .X(_23017_));
 sky130_fd_sc_hd__and4_4 _29452_ (.A(_23016_),
    .B(_23017_),
    .C(_22999_),
    .D(\count_instr[1] ),
    .X(_23018_));
 sky130_vsdinv _29453_ (.A(_23018_),
    .Y(_23019_));
 sky130_fd_sc_hd__nand2_4 _29454_ (.A(_23014_),
    .B(_23019_),
    .Y(_23020_));
 sky130_vsdinv _29455_ (.A(_23020_),
    .Y(_00079_));
 sky130_fd_sc_hd__buf_1 _29456_ (.A(_23015_),
    .X(_23021_));
 sky130_fd_sc_hd__buf_1 _29457_ (.A(_21985_),
    .X(_23022_));
 sky130_fd_sc_hd__buf_1 _29458_ (.A(\count_instr[2] ),
    .X(_23023_));
 sky130_fd_sc_hd__a41o_4 _29459_ (.A1(_23021_),
    .A2(_23022_),
    .A3(_23004_),
    .A4(_23010_),
    .B1(_23023_),
    .X(_23024_));
 sky130_fd_sc_hd__buf_1 _29460_ (.A(_23001_),
    .X(_23025_));
 sky130_fd_sc_hd__buf_1 _29461_ (.A(_23025_),
    .X(_23026_));
 sky130_fd_sc_hd__buf_1 _29462_ (.A(_23026_),
    .X(_23027_));
 sky130_fd_sc_hd__nand4_4 _29463_ (.A(_23004_),
    .B(_23027_),
    .C(_23010_),
    .D(_23023_),
    .Y(_23028_));
 sky130_fd_sc_hd__and3_4 _29464_ (.A(_23024_),
    .B(_19034_),
    .C(_23028_),
    .X(_00090_));
 sky130_fd_sc_hd__nand2_4 _29465_ (.A(_23028_),
    .B(\count_instr[3] ),
    .Y(_23029_));
 sky130_fd_sc_hd__buf_1 _29466_ (.A(_23021_),
    .X(_23030_));
 sky130_fd_sc_hd__buf_1 _29467_ (.A(_23022_),
    .X(_23031_));
 sky130_vsdinv _29468_ (.A(\count_instr[3] ),
    .Y(_23032_));
 sky130_fd_sc_hd__and4_4 _29469_ (.A(_23032_),
    .B(_23004_),
    .C(_23010_),
    .D(_23023_),
    .X(_23033_));
 sky130_fd_sc_hd__nand3_4 _29470_ (.A(_23030_),
    .B(_23031_),
    .C(_23033_),
    .Y(_23034_));
 sky130_fd_sc_hd__buf_1 _29471_ (.A(_19494_),
    .X(_23035_));
 sky130_fd_sc_hd__buf_1 _29472_ (.A(_23035_),
    .X(_23036_));
 sky130_fd_sc_hd__a21oi_4 _29473_ (.A1(_23029_),
    .A2(_23034_),
    .B1(_23036_),
    .Y(_00101_));
 sky130_fd_sc_hd__buf_1 _29474_ (.A(\count_instr[4] ),
    .X(_23037_));
 sky130_vsdinv _29475_ (.A(_19138_),
    .Y(_23038_));
 sky130_fd_sc_hd__and4_4 _29476_ (.A(\count_instr[0] ),
    .B(\count_instr[1] ),
    .C(\count_instr[2] ),
    .D(\count_instr[3] ),
    .X(_23039_));
 sky130_fd_sc_hd__buf_1 _29477_ (.A(_23039_),
    .X(_23040_));
 sky130_fd_sc_hd__buf_1 _29478_ (.A(_23040_),
    .X(_23041_));
 sky130_fd_sc_hd__and4_4 _29479_ (.A(_23038_),
    .B(_21927_),
    .C(_18407_),
    .D(_23041_),
    .X(_23042_));
 sky130_fd_sc_hd__buf_1 _29480_ (.A(_18536_),
    .X(_23043_));
 sky130_fd_sc_hd__o21a_4 _29481_ (.A1(_23037_),
    .A2(_23042_),
    .B1(_23043_),
    .X(_23044_));
 sky130_fd_sc_hd__buf_1 _29482_ (.A(_23015_),
    .X(_23045_));
 sky130_fd_sc_hd__buf_1 _29483_ (.A(_23041_),
    .X(_23046_));
 sky130_fd_sc_hd__and4_4 _29484_ (.A(_23045_),
    .B(_21951_),
    .C(_23037_),
    .D(_23046_),
    .X(_23047_));
 sky130_vsdinv _29485_ (.A(_23047_),
    .Y(_23048_));
 sky130_fd_sc_hd__nand2_4 _29486_ (.A(_23044_),
    .B(_23048_),
    .Y(_23049_));
 sky130_vsdinv _29487_ (.A(_23049_),
    .Y(_00112_));
 sky130_fd_sc_hd__buf_1 _29488_ (.A(_21927_),
    .X(_23050_));
 sky130_fd_sc_hd__buf_1 _29489_ (.A(_23050_),
    .X(_23051_));
 sky130_fd_sc_hd__buf_1 _29490_ (.A(_23016_),
    .X(_23052_));
 sky130_fd_sc_hd__buf_1 _29491_ (.A(_23046_),
    .X(_23053_));
 sky130_fd_sc_hd__nand2_4 _29492_ (.A(\count_instr[4] ),
    .B(\count_instr[5] ),
    .Y(_23054_));
 sky130_vsdinv _29493_ (.A(_23054_),
    .Y(_23055_));
 sky130_fd_sc_hd__buf_1 _29494_ (.A(_23055_),
    .X(_23056_));
 sky130_fd_sc_hd__a41oi_4 _29495_ (.A1(_23051_),
    .A2(_23052_),
    .A3(_23053_),
    .A4(_23056_),
    .B1(_19426_),
    .Y(_23057_));
 sky130_fd_sc_hd__o21a_4 _29496_ (.A1(\count_instr[5] ),
    .A2(_23047_),
    .B1(_23057_),
    .X(_00123_));
 sky130_fd_sc_hd__buf_1 _29497_ (.A(_23026_),
    .X(_23058_));
 sky130_fd_sc_hd__buf_1 _29498_ (.A(\count_instr[6] ),
    .X(_23059_));
 sky130_fd_sc_hd__and4_4 _29499_ (.A(_23058_),
    .B(_23059_),
    .C(_23053_),
    .D(_23056_),
    .X(_23060_));
 sky130_fd_sc_hd__buf_1 _29500_ (.A(_23041_),
    .X(_23061_));
 sky130_fd_sc_hd__and4_4 _29501_ (.A(_18780_),
    .B(_19101_),
    .C(_23061_),
    .D(_23056_),
    .X(_23062_));
 sky130_fd_sc_hd__buf_1 _29502_ (.A(_21128_),
    .X(_23063_));
 sky130_fd_sc_hd__o21ai_4 _29503_ (.A1(_23059_),
    .A2(_23062_),
    .B1(_23063_),
    .Y(_23064_));
 sky130_fd_sc_hd__nor2_4 _29504_ (.A(_23060_),
    .B(_23064_),
    .Y(_00128_));
 sky130_fd_sc_hd__buf_1 _29505_ (.A(_23001_),
    .X(_23065_));
 sky130_fd_sc_hd__buf_1 _29506_ (.A(_23065_),
    .X(_23066_));
 sky130_vsdinv _29507_ (.A(\count_instr[7] ),
    .Y(_23067_));
 sky130_fd_sc_hd__a41o_4 _29508_ (.A1(_23066_),
    .A2(_23059_),
    .A3(_23061_),
    .A4(_23056_),
    .B1(_23067_),
    .X(_23068_));
 sky130_fd_sc_hd__buf_1 _29509_ (.A(_23022_),
    .X(_23069_));
 sky130_fd_sc_hd__o21a_4 _29510_ (.A1(_18562_),
    .A2(_22104_),
    .B1(_19120_),
    .X(_23070_));
 sky130_fd_sc_hd__and4_4 _29511_ (.A(_23046_),
    .B(_23059_),
    .C(_23067_),
    .D(_23055_),
    .X(_23071_));
 sky130_fd_sc_hd__nand4_4 _29512_ (.A(_23069_),
    .B(_21990_),
    .C(_23070_),
    .D(_23071_),
    .Y(_23072_));
 sky130_fd_sc_hd__a21oi_4 _29513_ (.A1(_23068_),
    .A2(_23072_),
    .B1(_23036_),
    .Y(_00129_));
 sky130_fd_sc_hd__buf_1 _29514_ (.A(\count_instr[8] ),
    .X(_23073_));
 sky130_fd_sc_hd__and4_4 _29515_ (.A(_23037_),
    .B(\count_instr[5] ),
    .C(\count_instr[6] ),
    .D(\count_instr[7] ),
    .X(_23074_));
 sky130_fd_sc_hd__and4_4 _29516_ (.A(_23021_),
    .B(_21952_),
    .C(_23061_),
    .D(_23074_),
    .X(_23075_));
 sky130_fd_sc_hd__and4_4 _29517_ (.A(_23055_),
    .B(\count_instr[6] ),
    .C(\count_instr[7] ),
    .D(\count_instr[8] ),
    .X(_23076_));
 sky130_fd_sc_hd__buf_1 _29518_ (.A(_23076_),
    .X(_23077_));
 sky130_fd_sc_hd__buf_1 _29519_ (.A(_19425_),
    .X(_23078_));
 sky130_fd_sc_hd__a41oi_4 _29520_ (.A1(_23051_),
    .A2(_23052_),
    .A3(_23053_),
    .A4(_23077_),
    .B1(_23078_),
    .Y(_23079_));
 sky130_fd_sc_hd__o21a_4 _29521_ (.A1(_23073_),
    .A2(_23075_),
    .B1(_23079_),
    .X(_00130_));
 sky130_fd_sc_hd__buf_1 _29522_ (.A(\count_instr[9] ),
    .X(_23080_));
 sky130_fd_sc_hd__buf_1 _29523_ (.A(_23080_),
    .X(_23081_));
 sky130_fd_sc_hd__and3_4 _29524_ (.A(_23040_),
    .B(_23074_),
    .C(_23073_),
    .X(_23082_));
 sky130_fd_sc_hd__and4_4 _29525_ (.A(_23038_),
    .B(_23017_),
    .C(_18553_),
    .D(_23082_),
    .X(_23083_));
 sky130_fd_sc_hd__o21a_4 _29526_ (.A1(_23081_),
    .A2(_23083_),
    .B1(_19111_),
    .X(_23084_));
 sky130_fd_sc_hd__buf_1 _29527_ (.A(_23025_),
    .X(_23085_));
 sky130_fd_sc_hd__and4_4 _29528_ (.A(_23085_),
    .B(_23080_),
    .C(_23046_),
    .D(_23077_),
    .X(_23086_));
 sky130_vsdinv _29529_ (.A(_23086_),
    .Y(_23087_));
 sky130_fd_sc_hd__and2_4 _29530_ (.A(_23084_),
    .B(_23087_),
    .X(_00131_));
 sky130_fd_sc_hd__buf_1 _29531_ (.A(\count_instr[10] ),
    .X(_23088_));
 sky130_vsdinv _29532_ (.A(_23088_),
    .Y(_23089_));
 sky130_fd_sc_hd__a41o_4 _29533_ (.A1(_23066_),
    .A2(_23081_),
    .A3(_23061_),
    .A4(_23077_),
    .B1(_23089_),
    .X(_23090_));
 sky130_fd_sc_hd__buf_1 _29534_ (.A(_18780_),
    .X(_23091_));
 sky130_fd_sc_hd__and4_4 _29535_ (.A(_23089_),
    .B(_19121_),
    .C(_23073_),
    .D(_23080_),
    .X(_23092_));
 sky130_fd_sc_hd__nand4_4 _29536_ (.A(_23091_),
    .B(_23053_),
    .C(_23074_),
    .D(_23092_),
    .Y(_23093_));
 sky130_fd_sc_hd__a21oi_4 _29537_ (.A1(_23090_),
    .A2(_23093_),
    .B1(_23036_),
    .Y(_00069_));
 sky130_fd_sc_hd__buf_1 _29538_ (.A(\count_instr[11] ),
    .X(_23094_));
 sky130_fd_sc_hd__a41o_4 _29539_ (.A1(_23042_),
    .A2(_23080_),
    .A3(_23088_),
    .A4(_23077_),
    .B1(_23094_),
    .X(_23095_));
 sky130_fd_sc_hd__buf_1 _29540_ (.A(_18233_),
    .X(_23096_));
 sky130_fd_sc_hd__buf_1 _29541_ (.A(_23096_),
    .X(_23097_));
 sky130_fd_sc_hd__and4_4 _29542_ (.A(_23015_),
    .B(_21985_),
    .C(_23041_),
    .D(_23076_),
    .X(_23098_));
 sky130_fd_sc_hd__nand4_4 _29543_ (.A(_23081_),
    .B(_23098_),
    .C(_23088_),
    .D(_23094_),
    .Y(_23099_));
 sky130_fd_sc_hd__nand3_4 _29544_ (.A(_23095_),
    .B(_23097_),
    .C(_23099_),
    .Y(_23100_));
 sky130_vsdinv _29545_ (.A(_23100_),
    .Y(_00070_));
 sky130_fd_sc_hd__buf_1 _29546_ (.A(\count_instr[12] ),
    .X(_23101_));
 sky130_fd_sc_hd__and4_4 _29547_ (.A(_23098_),
    .B(_23081_),
    .C(_23088_),
    .D(_23094_),
    .X(_23102_));
 sky130_fd_sc_hd__buf_1 _29548_ (.A(_23038_),
    .X(_23103_));
 sky130_fd_sc_hd__buf_1 _29549_ (.A(_22072_),
    .X(_23104_));
 sky130_fd_sc_hd__nand3_4 _29550_ (.A(\count_instr[9] ),
    .B(\count_instr[10] ),
    .C(\count_instr[11] ),
    .Y(_23105_));
 sky130_vsdinv _29551_ (.A(_23105_),
    .Y(_23106_));
 sky130_fd_sc_hd__and4_4 _29552_ (.A(_23076_),
    .B(\count_instr[12] ),
    .C(_23040_),
    .D(_23106_),
    .X(_23107_));
 sky130_fd_sc_hd__buf_1 _29553_ (.A(_23107_),
    .X(_23108_));
 sky130_fd_sc_hd__a41oi_4 _29554_ (.A1(_23051_),
    .A2(_23103_),
    .A3(_23104_),
    .A4(_23108_),
    .B1(_23078_),
    .Y(_23109_));
 sky130_fd_sc_hd__o21a_4 _29555_ (.A1(_23101_),
    .A2(_23102_),
    .B1(_23109_),
    .X(_00071_));
 sky130_fd_sc_hd__buf_1 _29556_ (.A(\count_instr[13] ),
    .X(_23110_));
 sky130_fd_sc_hd__buf_1 _29557_ (.A(_23017_),
    .X(_23111_));
 sky130_fd_sc_hd__and4_4 _29558_ (.A(_23103_),
    .B(_23111_),
    .C(_22035_),
    .D(_23108_),
    .X(_23112_));
 sky130_fd_sc_hd__buf_1 _29559_ (.A(_23050_),
    .X(_23113_));
 sky130_fd_sc_hd__a41oi_4 _29560_ (.A1(_23113_),
    .A2(_23052_),
    .A3(_23110_),
    .A4(_23108_),
    .B1(_23078_),
    .Y(_23114_));
 sky130_fd_sc_hd__o21a_4 _29561_ (.A1(_23110_),
    .A2(_23112_),
    .B1(_23114_),
    .X(_00072_));
 sky130_fd_sc_hd__and4_4 _29562_ (.A(_23016_),
    .B(_23050_),
    .C(_23110_),
    .D(_23108_),
    .X(_23115_));
 sky130_fd_sc_hd__buf_1 _29563_ (.A(\count_instr[14] ),
    .X(_23116_));
 sky130_fd_sc_hd__and4_4 _29564_ (.A(_23040_),
    .B(_23074_),
    .C(\count_instr[8] ),
    .D(_23106_),
    .X(_23117_));
 sky130_fd_sc_hd__buf_1 _29565_ (.A(_23117_),
    .X(_23118_));
 sky130_fd_sc_hd__nand2_4 _29566_ (.A(_18266_),
    .B(_18481_),
    .Y(_23119_));
 sky130_vsdinv _29567_ (.A(_23119_),
    .Y(_23120_));
 sky130_fd_sc_hd__and4_4 _29568_ (.A(_23118_),
    .B(_23101_),
    .C(\count_instr[13] ),
    .D(_23120_),
    .X(_23121_));
 sky130_fd_sc_hd__and4_4 _29569_ (.A(_19103_),
    .B(_18553_),
    .C(_21928_),
    .D(_23121_),
    .X(_23122_));
 sky130_fd_sc_hd__o21a_4 _29570_ (.A1(_23116_),
    .A2(_23122_),
    .B1(_19111_),
    .X(_23123_));
 sky130_fd_sc_hd__a21boi_4 _29571_ (.A1(_23115_),
    .A2(_23116_),
    .B1_N(_23123_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand3_4 _29572_ (.A(_23101_),
    .B(\count_instr[13] ),
    .C(\count_instr[14] ),
    .Y(_23124_));
 sky130_fd_sc_hd__nor4_4 _29573_ (.A(_18268_),
    .B(\count_instr[15] ),
    .C(_23124_),
    .D(_19136_),
    .Y(_23125_));
 sky130_fd_sc_hd__and2_4 _29574_ (.A(_23118_),
    .B(_23125_),
    .X(_23126_));
 sky130_fd_sc_hd__and4_4 _29575_ (.A(_19104_),
    .B(_23111_),
    .C(_19106_),
    .D(_23126_),
    .X(_23127_));
 sky130_fd_sc_hd__a21boi_4 _29576_ (.A1(_23115_),
    .A2(_23116_),
    .B1_N(\count_instr[15] ),
    .Y(_23128_));
 sky130_fd_sc_hd__buf_1 _29577_ (.A(_22929_),
    .X(_23129_));
 sky130_fd_sc_hd__o21a_4 _29578_ (.A1(_23127_),
    .A2(_23128_),
    .B1(_23129_),
    .X(_00074_));
 sky130_fd_sc_hd__buf_1 _29579_ (.A(\count_instr[16] ),
    .X(_23130_));
 sky130_fd_sc_hd__buf_1 _29580_ (.A(_23130_),
    .X(_23131_));
 sky130_fd_sc_hd__buf_1 _29581_ (.A(_21973_),
    .X(_23132_));
 sky130_fd_sc_hd__nand4_4 _29582_ (.A(\count_instr[12] ),
    .B(\count_instr[13] ),
    .C(\count_instr[14] ),
    .D(\count_instr[15] ),
    .Y(_23133_));
 sky130_vsdinv _29583_ (.A(_23133_),
    .Y(_23134_));
 sky130_fd_sc_hd__and4_4 _29584_ (.A(_23076_),
    .B(_23039_),
    .C(_23106_),
    .D(_23134_),
    .X(_23135_));
 sky130_fd_sc_hd__buf_1 _29585_ (.A(_23135_),
    .X(_23136_));
 sky130_fd_sc_hd__buf_1 _29586_ (.A(_23136_),
    .X(_23137_));
 sky130_vsdinv _29587_ (.A(_23137_),
    .Y(_23138_));
 sky130_fd_sc_hd__buf_1 _29588_ (.A(_19138_),
    .X(_23139_));
 sky130_fd_sc_hd__nor4_4 _29589_ (.A(_21958_),
    .B(_23132_),
    .C(_23138_),
    .D(_23139_),
    .Y(_23140_));
 sky130_fd_sc_hd__o21a_4 _29590_ (.A1(_23131_),
    .A2(_23140_),
    .B1(_23043_),
    .X(_23141_));
 sky130_fd_sc_hd__buf_1 _29591_ (.A(_23016_),
    .X(_23142_));
 sky130_fd_sc_hd__buf_1 _29592_ (.A(_23137_),
    .X(_23143_));
 sky130_fd_sc_hd__nand4_4 _29593_ (.A(_23113_),
    .B(_23142_),
    .C(_23131_),
    .D(_23143_),
    .Y(_23144_));
 sky130_fd_sc_hd__nand2_4 _29594_ (.A(_23141_),
    .B(_23144_),
    .Y(_23145_));
 sky130_vsdinv _29595_ (.A(_23145_),
    .Y(_00075_));
 sky130_fd_sc_hd__buf_1 _29596_ (.A(\count_instr[17] ),
    .X(_23146_));
 sky130_fd_sc_hd__and4_4 _29597_ (.A(_23065_),
    .B(_23131_),
    .C(_23146_),
    .D(_23143_),
    .X(_23147_));
 sky130_fd_sc_hd__buf_1 _29598_ (.A(_23134_),
    .X(_23148_));
 sky130_fd_sc_hd__nand3_4 _29599_ (.A(_23118_),
    .B(_23130_),
    .C(_23148_),
    .Y(_23149_));
 sky130_fd_sc_hd__nor4_4 _29600_ (.A(_19135_),
    .B(_21974_),
    .C(_23149_),
    .D(_23139_),
    .Y(_23150_));
 sky130_fd_sc_hd__o21ai_4 _29601_ (.A1(_23146_),
    .A2(_23150_),
    .B1(_23096_),
    .Y(_23151_));
 sky130_fd_sc_hd__or2_4 _29602_ (.A(_23147_),
    .B(_23151_),
    .X(_23152_));
 sky130_vsdinv _29603_ (.A(_23152_),
    .Y(_00076_));
 sky130_fd_sc_hd__nand3_4 _29604_ (.A(_23130_),
    .B(_23146_),
    .C(\count_instr[18] ),
    .Y(_23153_));
 sky130_vsdinv _29605_ (.A(_23140_),
    .Y(_23154_));
 sky130_fd_sc_hd__buf_1 _29606_ (.A(_23120_),
    .X(_23155_));
 sky130_fd_sc_hd__and4_4 _29607_ (.A(_23136_),
    .B(_23130_),
    .C(\count_instr[17] ),
    .D(_23155_),
    .X(_23156_));
 sky130_fd_sc_hd__and4_4 _29608_ (.A(_19103_),
    .B(_21953_),
    .C(_21928_),
    .D(_23156_),
    .X(_23157_));
 sky130_fd_sc_hd__o21a_4 _29609_ (.A1(\count_instr[18] ),
    .A2(_23157_),
    .B1(_19111_),
    .X(_23158_));
 sky130_fd_sc_hd__o21a_4 _29610_ (.A1(_23153_),
    .A2(_23154_),
    .B1(_23158_),
    .X(_00077_));
 sky130_fd_sc_hd__buf_1 _29611_ (.A(_23050_),
    .X(_23159_));
 sky130_vsdinv _29612_ (.A(_23153_),
    .Y(_23160_));
 sky130_vsdinv _29613_ (.A(\count_instr[19] ),
    .Y(_23161_));
 sky130_fd_sc_hd__a41o_4 _29614_ (.A1(_23052_),
    .A2(_23159_),
    .A3(_23143_),
    .A4(_23160_),
    .B1(_23161_),
    .X(_23162_));
 sky130_fd_sc_hd__and4_4 _29615_ (.A(_23143_),
    .B(_23161_),
    .C(_23070_),
    .D(_23160_),
    .X(_23163_));
 sky130_fd_sc_hd__nand4_4 _29616_ (.A(_23069_),
    .B(_19113_),
    .C(_19107_),
    .D(_23163_),
    .Y(_23164_));
 sky130_fd_sc_hd__a21oi_4 _29617_ (.A1(_23162_),
    .A2(_23164_),
    .B1(_23036_),
    .Y(_00078_));
 sky130_fd_sc_hd__buf_1 _29618_ (.A(_23026_),
    .X(_23165_));
 sky130_fd_sc_hd__nand4_4 _29619_ (.A(\count_instr[16] ),
    .B(\count_instr[17] ),
    .C(\count_instr[18] ),
    .D(\count_instr[19] ),
    .Y(_23166_));
 sky130_vsdinv _29620_ (.A(_23166_),
    .Y(_23167_));
 sky130_fd_sc_hd__buf_1 _29621_ (.A(_23167_),
    .X(_23168_));
 sky130_fd_sc_hd__and4_4 _29622_ (.A(_23117_),
    .B(\count_instr[20] ),
    .C(_23148_),
    .D(_23168_),
    .X(_23169_));
 sky130_fd_sc_hd__buf_1 _29623_ (.A(\count_instr[20] ),
    .X(_23170_));
 sky130_fd_sc_hd__buf_1 _29624_ (.A(_23167_),
    .X(_23171_));
 sky130_fd_sc_hd__and4_4 _29625_ (.A(_23117_),
    .B(_18849_),
    .C(_23148_),
    .D(_23171_),
    .X(_23172_));
 sky130_vsdinv _29626_ (.A(_23172_),
    .Y(_23173_));
 sky130_fd_sc_hd__nor3_4 _29627_ (.A(_23132_),
    .B(_23173_),
    .C(_21929_),
    .Y(_23174_));
 sky130_fd_sc_hd__buf_1 _29628_ (.A(_18506_),
    .X(_23175_));
 sky130_fd_sc_hd__o21ai_4 _29629_ (.A1(_23170_),
    .A2(_23174_),
    .B1(_23175_),
    .Y(_23176_));
 sky130_fd_sc_hd__a21o_4 _29630_ (.A1(_23165_),
    .A2(_23169_),
    .B1(_23176_),
    .X(_23177_));
 sky130_vsdinv _29631_ (.A(_23177_),
    .Y(_00080_));
 sky130_fd_sc_hd__buf_1 _29632_ (.A(\count_instr[21] ),
    .X(_23178_));
 sky130_vsdinv _29633_ (.A(_23169_),
    .Y(_23179_));
 sky130_fd_sc_hd__nor4_4 _29634_ (.A(_23011_),
    .B(_21926_),
    .C(_23179_),
    .D(_23012_),
    .Y(_23180_));
 sky130_fd_sc_hd__o21a_4 _29635_ (.A1(_23178_),
    .A2(_23180_),
    .B1(_23043_),
    .X(_23181_));
 sky130_fd_sc_hd__and4_4 _29636_ (.A(_23045_),
    .B(_21951_),
    .C(_23178_),
    .D(_23169_),
    .X(_23182_));
 sky130_vsdinv _29637_ (.A(_23182_),
    .Y(_23183_));
 sky130_fd_sc_hd__nand2_4 _29638_ (.A(_23181_),
    .B(_23183_),
    .Y(_23184_));
 sky130_vsdinv _29639_ (.A(_23184_),
    .Y(_00081_));
 sky130_fd_sc_hd__buf_1 _29640_ (.A(\count_instr[22] ),
    .X(_23185_));
 sky130_fd_sc_hd__and4_4 _29641_ (.A(_23058_),
    .B(_23178_),
    .C(_23185_),
    .D(_23169_),
    .X(_23186_));
 sky130_fd_sc_hd__and4_4 _29642_ (.A(_18779_),
    .B(_23170_),
    .C(_23178_),
    .D(_23172_),
    .X(_23187_));
 sky130_fd_sc_hd__o21ai_4 _29643_ (.A1(_23185_),
    .A2(_23187_),
    .B1(_18862_),
    .Y(_23188_));
 sky130_fd_sc_hd__nor2_4 _29644_ (.A(_23186_),
    .B(_23188_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand3_4 _29645_ (.A(_23170_),
    .B(\count_instr[21] ),
    .C(\count_instr[22] ),
    .Y(_23189_));
 sky130_fd_sc_hd__nor4_4 _29646_ (.A(_18267_),
    .B(\count_instr[23] ),
    .C(_23189_),
    .D(_19136_),
    .Y(_23190_));
 sky130_fd_sc_hd__and3_4 _29647_ (.A(_23137_),
    .B(_23168_),
    .C(_23190_),
    .X(_23191_));
 sky130_fd_sc_hd__and4_4 _29648_ (.A(_19104_),
    .B(_23111_),
    .C(_19106_),
    .D(_23191_),
    .X(_23192_));
 sky130_fd_sc_hd__a21boi_4 _29649_ (.A1(_23182_),
    .A2(_23185_),
    .B1_N(\count_instr[23] ),
    .Y(_23193_));
 sky130_fd_sc_hd__o21a_4 _29650_ (.A1(_23192_),
    .A2(_23193_),
    .B1(_23129_),
    .X(_00083_));
 sky130_fd_sc_hd__nand4_4 _29651_ (.A(\count_instr[20] ),
    .B(\count_instr[21] ),
    .C(\count_instr[22] ),
    .D(\count_instr[23] ),
    .Y(_23194_));
 sky130_vsdinv _29652_ (.A(_23194_),
    .Y(_23195_));
 sky130_fd_sc_hd__and4_4 _29653_ (.A(_23136_),
    .B(\count_instr[24] ),
    .C(_23171_),
    .D(_23195_),
    .X(_23196_));
 sky130_fd_sc_hd__buf_1 _29654_ (.A(_23196_),
    .X(_23197_));
 sky130_fd_sc_hd__buf_1 _29655_ (.A(\count_instr[24] ),
    .X(_23198_));
 sky130_fd_sc_hd__buf_1 _29656_ (.A(_23195_),
    .X(_23199_));
 sky130_fd_sc_hd__and4_4 _29657_ (.A(_23136_),
    .B(_18541_),
    .C(_23171_),
    .D(_23199_),
    .X(_23200_));
 sky130_vsdinv _29658_ (.A(_23200_),
    .Y(_23201_));
 sky130_fd_sc_hd__nor3_4 _29659_ (.A(_23132_),
    .B(_23201_),
    .C(_23139_),
    .Y(_23202_));
 sky130_fd_sc_hd__o21ai_4 _29660_ (.A1(_23198_),
    .A2(_23202_),
    .B1(_23175_),
    .Y(_23203_));
 sky130_fd_sc_hd__a21o_4 _29661_ (.A1(_23165_),
    .A2(_23197_),
    .B1(_23203_),
    .X(_23204_));
 sky130_vsdinv _29662_ (.A(_23204_),
    .Y(_00084_));
 sky130_fd_sc_hd__buf_1 _29663_ (.A(\count_instr[25] ),
    .X(_23205_));
 sky130_fd_sc_hd__buf_1 _29664_ (.A(_23205_),
    .X(_23206_));
 sky130_vsdinv _29665_ (.A(_23196_),
    .Y(_23207_));
 sky130_fd_sc_hd__nor4_4 _29666_ (.A(_23011_),
    .B(_23132_),
    .C(_23207_),
    .D(_23139_),
    .Y(_23208_));
 sky130_fd_sc_hd__o21a_4 _29667_ (.A1(_23206_),
    .A2(_23208_),
    .B1(_23043_),
    .X(_23209_));
 sky130_fd_sc_hd__and4_4 _29668_ (.A(_23045_),
    .B(_21951_),
    .C(_23205_),
    .D(_23197_),
    .X(_23210_));
 sky130_vsdinv _29669_ (.A(_23210_),
    .Y(_23211_));
 sky130_fd_sc_hd__nand2_4 _29670_ (.A(_23209_),
    .B(_23211_),
    .Y(_23212_));
 sky130_vsdinv _29671_ (.A(_23212_),
    .Y(_00085_));
 sky130_fd_sc_hd__buf_1 _29672_ (.A(\count_instr[26] ),
    .X(_23213_));
 sky130_vsdinv _29673_ (.A(_23213_),
    .Y(_23214_));
 sky130_fd_sc_hd__a41o_4 _29674_ (.A1(_23142_),
    .A2(_23159_),
    .A3(_23206_),
    .A4(_23197_),
    .B1(_23214_),
    .X(_23215_));
 sky130_fd_sc_hd__and4_4 _29675_ (.A(_23214_),
    .B(_19121_),
    .C(_23198_),
    .D(_23206_),
    .X(_23216_));
 sky130_fd_sc_hd__nand4_4 _29676_ (.A(_23104_),
    .B(_19075_),
    .C(_23200_),
    .D(_23216_),
    .Y(_23217_));
 sky130_fd_sc_hd__buf_1 _29677_ (.A(_23035_),
    .X(_23218_));
 sky130_fd_sc_hd__a21oi_4 _29678_ (.A1(_23215_),
    .A2(_23217_),
    .B1(_23218_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand4_4 _29679_ (.A(_23206_),
    .B(_23027_),
    .C(_23213_),
    .D(_23197_),
    .Y(_23219_));
 sky130_fd_sc_hd__nand2_4 _29680_ (.A(_23219_),
    .B(\count_instr[27] ),
    .Y(_23220_));
 sky130_fd_sc_hd__and4_4 _29681_ (.A(_23118_),
    .B(_23148_),
    .C(_23168_),
    .D(_23199_),
    .X(_23221_));
 sky130_fd_sc_hd__nand3_4 _29682_ (.A(_23198_),
    .B(_23205_),
    .C(_23213_),
    .Y(_23222_));
 sky130_fd_sc_hd__nor4_4 _29683_ (.A(_18479_),
    .B(\count_instr[27] ),
    .C(_23222_),
    .D(_21974_),
    .Y(_23223_));
 sky130_fd_sc_hd__and2_4 _29684_ (.A(_23221_),
    .B(_23223_),
    .X(_23224_));
 sky130_fd_sc_hd__nand4_4 _29685_ (.A(_23069_),
    .B(_19113_),
    .C(_23224_),
    .D(_19107_),
    .Y(_23225_));
 sky130_fd_sc_hd__a21oi_4 _29686_ (.A1(_23220_),
    .A2(_23225_),
    .B1(_23218_),
    .Y(_00087_));
 sky130_fd_sc_hd__and4_4 _29687_ (.A(_23082_),
    .B(_23106_),
    .C(_23134_),
    .D(_23171_),
    .X(_23226_));
 sky130_fd_sc_hd__nand4_4 _29688_ (.A(\count_instr[24] ),
    .B(\count_instr[25] ),
    .C(\count_instr[26] ),
    .D(\count_instr[27] ),
    .Y(_23227_));
 sky130_vsdinv _29689_ (.A(_23227_),
    .Y(_23228_));
 sky130_fd_sc_hd__and4_4 _29690_ (.A(_23226_),
    .B(_21927_),
    .C(_23199_),
    .D(_23228_),
    .X(_23229_));
 sky130_fd_sc_hd__nand4_4 _29691_ (.A(_19101_),
    .B(_18576_),
    .C(_22072_),
    .D(_23229_),
    .Y(_23230_));
 sky130_vsdinv _29692_ (.A(\count_instr[28] ),
    .Y(_23231_));
 sky130_fd_sc_hd__nand4_4 _29693_ (.A(_23135_),
    .B(_23167_),
    .C(_23195_),
    .D(_23228_),
    .Y(_23232_));
 sky130_fd_sc_hd__nor2_4 _29694_ (.A(_23231_),
    .B(_23232_),
    .Y(_23233_));
 sky130_vsdinv _29695_ (.A(_23233_),
    .Y(_23234_));
 sky130_fd_sc_hd__nor4_4 _29696_ (.A(_22708_),
    .B(_21926_),
    .C(_23234_),
    .D(_23012_),
    .Y(_23235_));
 sky130_fd_sc_hd__a211o_4 _29697_ (.A1(_23230_),
    .A2(_23231_),
    .B1(_22992_),
    .C1(_23235_),
    .X(_23236_));
 sky130_vsdinv _29698_ (.A(_23236_),
    .Y(_00088_));
 sky130_vsdinv _29699_ (.A(_23235_),
    .Y(_23237_));
 sky130_vsdinv _29700_ (.A(\count_instr[29] ),
    .Y(_23238_));
 sky130_fd_sc_hd__nor3_4 _29701_ (.A(_23231_),
    .B(_23238_),
    .C(_23232_),
    .Y(_23239_));
 sky130_fd_sc_hd__a41o_4 _29702_ (.A1(_23103_),
    .A2(_23159_),
    .A3(_21954_),
    .A4(_23239_),
    .B1(_18783_),
    .X(_23240_));
 sky130_fd_sc_hd__a21oi_4 _29703_ (.A1(_23237_),
    .A2(_23238_),
    .B1(_23240_),
    .Y(_00089_));
 sky130_vsdinv _29704_ (.A(\count_instr[30] ),
    .Y(_23241_));
 sky130_fd_sc_hd__a41o_4 _29705_ (.A1(_23103_),
    .A2(_21952_),
    .A3(_21954_),
    .A4(_23239_),
    .B1(_23241_),
    .X(_23242_));
 sky130_fd_sc_hd__and4_4 _29706_ (.A(_23241_),
    .B(_18851_),
    .C(\count_instr[28] ),
    .D(\count_instr[29] ),
    .X(_23243_));
 sky130_fd_sc_hd__nand4_4 _29707_ (.A(_23104_),
    .B(_19075_),
    .C(_23229_),
    .D(_23243_),
    .Y(_23244_));
 sky130_fd_sc_hd__a21oi_4 _29708_ (.A1(_23242_),
    .A2(_23244_),
    .B1(_23218_),
    .Y(_00091_));
 sky130_fd_sc_hd__nand4_4 _29709_ (.A(_23113_),
    .B(_23142_),
    .C(\count_instr[30] ),
    .D(_23239_),
    .Y(_23245_));
 sky130_fd_sc_hd__nand2_4 _29710_ (.A(_23245_),
    .B(\count_instr[31] ),
    .Y(_23246_));
 sky130_fd_sc_hd__and4_4 _29711_ (.A(_23137_),
    .B(_23168_),
    .C(_23199_),
    .D(_23228_),
    .X(_23247_));
 sky130_fd_sc_hd__nor3_4 _29712_ (.A(\count_instr[31] ),
    .B(_18550_),
    .C(_23241_),
    .Y(_23248_));
 sky130_fd_sc_hd__and4_4 _29713_ (.A(_23247_),
    .B(\count_instr[28] ),
    .C(\count_instr[29] ),
    .D(_23248_),
    .X(_23249_));
 sky130_fd_sc_hd__nand2_4 _29714_ (.A(_23091_),
    .B(_23249_),
    .Y(_23250_));
 sky130_fd_sc_hd__a21oi_4 _29715_ (.A1(_23246_),
    .A2(_23250_),
    .B1(_23218_),
    .Y(_00092_));
 sky130_fd_sc_hd__buf_1 _29716_ (.A(\count_instr[32] ),
    .X(_23251_));
 sky130_fd_sc_hd__nand2_4 _29717_ (.A(\count_instr[30] ),
    .B(\count_instr[31] ),
    .Y(_23252_));
 sky130_fd_sc_hd__nor4_4 _29718_ (.A(_23231_),
    .B(_23238_),
    .C(_23252_),
    .D(_23232_),
    .Y(_23253_));
 sky130_fd_sc_hd__buf_1 _29719_ (.A(_23253_),
    .X(_23254_));
 sky130_fd_sc_hd__and2_4 _29720_ (.A(_23254_),
    .B(_23017_),
    .X(_23255_));
 sky130_fd_sc_hd__and2_4 _29721_ (.A(_23255_),
    .B(_23142_),
    .X(_23256_));
 sky130_fd_sc_hd__buf_1 _29722_ (.A(_23026_),
    .X(_23257_));
 sky130_fd_sc_hd__and2_4 _29723_ (.A(_23254_),
    .B(_23251_),
    .X(_23258_));
 sky130_fd_sc_hd__a21oi_4 _29724_ (.A1(_23257_),
    .A2(_23258_),
    .B1(_20430_),
    .Y(_23259_));
 sky130_fd_sc_hd__o21a_4 _29725_ (.A1(_23251_),
    .A2(_23256_),
    .B1(_23259_),
    .X(_00093_));
 sky130_fd_sc_hd__buf_1 _29726_ (.A(\count_instr[33] ),
    .X(_23260_));
 sky130_fd_sc_hd__and3_4 _29727_ (.A(_23258_),
    .B(_23045_),
    .C(_21985_),
    .X(_23261_));
 sky130_fd_sc_hd__buf_1 _29728_ (.A(_18375_),
    .X(_23262_));
 sky130_fd_sc_hd__buf_1 _29729_ (.A(_23262_),
    .X(_23263_));
 sky130_fd_sc_hd__o21a_4 _29730_ (.A1(_23260_),
    .A2(_23261_),
    .B1(_23263_),
    .X(_23264_));
 sky130_fd_sc_hd__and3_4 _29731_ (.A(_23253_),
    .B(\count_instr[32] ),
    .C(_23260_),
    .X(_23265_));
 sky130_fd_sc_hd__buf_1 _29732_ (.A(_23265_),
    .X(_23266_));
 sky130_fd_sc_hd__and2_4 _29733_ (.A(_23065_),
    .B(_23266_),
    .X(_23267_));
 sky130_vsdinv _29734_ (.A(_23267_),
    .Y(_23268_));
 sky130_fd_sc_hd__nand2_4 _29735_ (.A(_23264_),
    .B(_23268_),
    .Y(_23269_));
 sky130_vsdinv _29736_ (.A(_23269_),
    .Y(_00094_));
 sky130_fd_sc_hd__buf_1 _29737_ (.A(\count_instr[34] ),
    .X(_23270_));
 sky130_vsdinv _29738_ (.A(_23270_),
    .Y(_23271_));
 sky130_fd_sc_hd__a21o_4 _29739_ (.A1(_23257_),
    .A2(_23266_),
    .B1(_23271_),
    .X(_23272_));
 sky130_fd_sc_hd__buf_1 _29740_ (.A(_18545_),
    .X(_23273_));
 sky130_vsdinv _29741_ (.A(_23273_),
    .Y(_23274_));
 sky130_fd_sc_hd__buf_1 _29742_ (.A(_23274_),
    .X(_23275_));
 sky130_fd_sc_hd__nand2_4 _29743_ (.A(_23251_),
    .B(_23260_),
    .Y(_23276_));
 sky130_fd_sc_hd__nor3_4 _29744_ (.A(_23270_),
    .B(_18551_),
    .C(_23276_),
    .Y(_23277_));
 sky130_fd_sc_hd__nand4_4 _29745_ (.A(_23069_),
    .B(_23275_),
    .C(_23254_),
    .D(_23277_),
    .Y(_23278_));
 sky130_fd_sc_hd__buf_1 _29746_ (.A(_23035_),
    .X(_23279_));
 sky130_fd_sc_hd__a21oi_4 _29747_ (.A1(_23272_),
    .A2(_23278_),
    .B1(_23279_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand3_4 _29748_ (.A(_23257_),
    .B(_23266_),
    .C(_23270_),
    .Y(_23280_));
 sky130_fd_sc_hd__nand2_4 _29749_ (.A(_23280_),
    .B(\count_instr[35] ),
    .Y(_23281_));
 sky130_fd_sc_hd__nor4_4 _29750_ (.A(_19091_),
    .B(_23271_),
    .C(\count_instr[35] ),
    .D(_23276_),
    .Y(_23282_));
 sky130_fd_sc_hd__nand3_4 _29751_ (.A(_23091_),
    .B(_23254_),
    .C(_23282_),
    .Y(_23283_));
 sky130_fd_sc_hd__a21oi_4 _29752_ (.A1(_23281_),
    .A2(_23283_),
    .B1(_23279_),
    .Y(_00096_));
 sky130_fd_sc_hd__nand2_4 _29753_ (.A(\count_instr[34] ),
    .B(\count_instr[35] ),
    .Y(_23284_));
 sky130_vsdinv _29754_ (.A(_23284_),
    .Y(_23285_));
 sky130_fd_sc_hd__and4_4 _29755_ (.A(_23253_),
    .B(\count_instr[32] ),
    .C(\count_instr[33] ),
    .D(_23285_),
    .X(_23286_));
 sky130_fd_sc_hd__buf_1 _29756_ (.A(\count_instr[36] ),
    .X(_23287_));
 sky130_fd_sc_hd__and3_4 _29757_ (.A(_23286_),
    .B(_23025_),
    .C(_23287_),
    .X(_23288_));
 sky130_fd_sc_hd__buf_1 _29758_ (.A(\count_instr[36] ),
    .X(_23289_));
 sky130_fd_sc_hd__a41oi_4 _29759_ (.A1(_23051_),
    .A2(_23266_),
    .A3(_23030_),
    .A4(_23285_),
    .B1(_23289_),
    .Y(_23290_));
 sky130_fd_sc_hd__nor3_4 _29760_ (.A(_18934_),
    .B(_23288_),
    .C(_23290_),
    .Y(_00097_));
 sky130_fd_sc_hd__buf_1 _29761_ (.A(\count_instr[37] ),
    .X(_23291_));
 sky130_fd_sc_hd__buf_1 _29762_ (.A(_23291_),
    .X(_23292_));
 sky130_fd_sc_hd__o21a_4 _29763_ (.A1(_23292_),
    .A2(_23288_),
    .B1(_23263_),
    .X(_23293_));
 sky130_fd_sc_hd__buf_1 _29764_ (.A(_23286_),
    .X(_23294_));
 sky130_fd_sc_hd__and4_4 _29765_ (.A(_23294_),
    .B(_23005_),
    .C(_23287_),
    .D(_23291_),
    .X(_23295_));
 sky130_vsdinv _29766_ (.A(_23295_),
    .Y(_23296_));
 sky130_fd_sc_hd__nand2_4 _29767_ (.A(_23293_),
    .B(_23296_),
    .Y(_23297_));
 sky130_vsdinv _29768_ (.A(_23297_),
    .Y(_00098_));
 sky130_vsdinv _29769_ (.A(\count_instr[38] ),
    .Y(_23298_));
 sky130_fd_sc_hd__a41o_4 _29770_ (.A1(_23294_),
    .A2(_23027_),
    .A3(_23289_),
    .A4(_23292_),
    .B1(_23298_),
    .X(_23299_));
 sky130_fd_sc_hd__and4_4 _29771_ (.A(_23298_),
    .B(_18851_),
    .C(_23287_),
    .D(_23291_),
    .X(_23300_));
 sky130_fd_sc_hd__nand4_4 _29772_ (.A(_23031_),
    .B(_23294_),
    .C(_23275_),
    .D(_23300_),
    .Y(_23301_));
 sky130_fd_sc_hd__a21oi_4 _29773_ (.A1(_23299_),
    .A2(_23301_),
    .B1(_23279_),
    .Y(_00099_));
 sky130_fd_sc_hd__and3_4 _29774_ (.A(_23286_),
    .B(_23287_),
    .C(_23291_),
    .X(_23302_));
 sky130_fd_sc_hd__nand3_4 _29775_ (.A(_23302_),
    .B(\count_instr[38] ),
    .C(_23058_),
    .Y(_23303_));
 sky130_fd_sc_hd__nand2_4 _29776_ (.A(_23303_),
    .B(\count_instr[39] ),
    .Y(_23304_));
 sky130_fd_sc_hd__nor3_4 _29777_ (.A(\count_instr[39] ),
    .B(_18550_),
    .C(_23298_),
    .Y(_23305_));
 sky130_fd_sc_hd__and3_4 _29778_ (.A(_23305_),
    .B(_23289_),
    .C(_23292_),
    .X(_23306_));
 sky130_fd_sc_hd__nand3_4 _29779_ (.A(_23294_),
    .B(_23091_),
    .C(_23306_),
    .Y(_23307_));
 sky130_fd_sc_hd__a21oi_4 _29780_ (.A1(_23304_),
    .A2(_23307_),
    .B1(_23279_),
    .Y(_00100_));
 sky130_fd_sc_hd__buf_1 _29781_ (.A(\count_instr[40] ),
    .X(_23308_));
 sky130_fd_sc_hd__buf_1 _29782_ (.A(_23308_),
    .X(_23309_));
 sky130_vsdinv _29783_ (.A(_23309_),
    .Y(_23310_));
 sky130_fd_sc_hd__nand2_4 _29784_ (.A(\count_instr[38] ),
    .B(\count_instr[39] ),
    .Y(_23311_));
 sky130_vsdinv _29785_ (.A(_23311_),
    .Y(_23312_));
 sky130_fd_sc_hd__and4_4 _29786_ (.A(_23286_),
    .B(\count_instr[36] ),
    .C(\count_instr[37] ),
    .D(_23312_),
    .X(_23313_));
 sky130_fd_sc_hd__buf_1 _29787_ (.A(_23313_),
    .X(_23314_));
 sky130_fd_sc_hd__nand3_4 _29788_ (.A(_23314_),
    .B(_23031_),
    .C(_23030_),
    .Y(_23315_));
 sky130_fd_sc_hd__a41o_4 _29789_ (.A1(_23302_),
    .A2(_23309_),
    .A3(_23066_),
    .A4(_23312_),
    .B1(_18530_),
    .X(_23316_));
 sky130_fd_sc_hd__a21oi_4 _29790_ (.A1(_23310_),
    .A2(_23315_),
    .B1(_23316_),
    .Y(_00102_));
 sky130_fd_sc_hd__buf_1 _29791_ (.A(\count_instr[41] ),
    .X(_23317_));
 sky130_fd_sc_hd__buf_1 _29792_ (.A(_23317_),
    .X(_23318_));
 sky130_fd_sc_hd__and3_4 _29793_ (.A(_23313_),
    .B(\count_instr[40] ),
    .C(_23005_),
    .X(_23319_));
 sky130_fd_sc_hd__o21a_4 _29794_ (.A1(_23318_),
    .A2(_23319_),
    .B1(_23263_),
    .X(_23320_));
 sky130_fd_sc_hd__and4_4 _29795_ (.A(_23314_),
    .B(_23308_),
    .C(_23317_),
    .D(_23005_),
    .X(_23321_));
 sky130_vsdinv _29796_ (.A(_23321_),
    .Y(_23322_));
 sky130_fd_sc_hd__nand2_4 _29797_ (.A(_23320_),
    .B(_23322_),
    .Y(_23323_));
 sky130_vsdinv _29798_ (.A(_23323_),
    .Y(_00103_));
 sky130_fd_sc_hd__buf_1 _29799_ (.A(\count_instr[42] ),
    .X(_23324_));
 sky130_vsdinv _29800_ (.A(_23324_),
    .Y(_23325_));
 sky130_fd_sc_hd__nand4_4 _29801_ (.A(_19115_),
    .B(_23325_),
    .C(_23309_),
    .D(_23318_),
    .Y(_23326_));
 sky130_fd_sc_hd__nand3_4 _29802_ (.A(_23302_),
    .B(_21952_),
    .C(_23312_),
    .Y(_23327_));
 sky130_fd_sc_hd__nor3_4 _29803_ (.A(_23273_),
    .B(_23326_),
    .C(_23327_),
    .Y(_23328_));
 sky130_fd_sc_hd__a41oi_4 _29804_ (.A1(_23309_),
    .A2(_23314_),
    .A3(_23318_),
    .A4(_23058_),
    .B1(_23325_),
    .Y(_23329_));
 sky130_fd_sc_hd__o21a_4 _29805_ (.A1(_23328_),
    .A2(_23329_),
    .B1(_23129_),
    .X(_00104_));
 sky130_vsdinv _29806_ (.A(\count_instr[43] ),
    .Y(_23330_));
 sky130_fd_sc_hd__a21o_4 _29807_ (.A1(_23321_),
    .A2(_23324_),
    .B1(_23330_),
    .X(_23331_));
 sky130_fd_sc_hd__and3_4 _29808_ (.A(_23330_),
    .B(_19120_),
    .C(\count_instr[42] ),
    .X(_23332_));
 sky130_fd_sc_hd__and3_4 _29809_ (.A(_23332_),
    .B(_23308_),
    .C(_23318_),
    .X(_23333_));
 sky130_fd_sc_hd__nand3_4 _29810_ (.A(_23314_),
    .B(_18781_),
    .C(_23333_),
    .Y(_23334_));
 sky130_fd_sc_hd__buf_1 _29811_ (.A(_23035_),
    .X(_23335_));
 sky130_fd_sc_hd__a21oi_4 _29812_ (.A1(_23331_),
    .A2(_23334_),
    .B1(_23335_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand3_4 _29813_ (.A(_23321_),
    .B(_23324_),
    .C(\count_instr[43] ),
    .Y(_23336_));
 sky130_fd_sc_hd__buf_1 _29814_ (.A(\count_instr[44] ),
    .X(_23337_));
 sky130_vsdinv _29815_ (.A(_23337_),
    .Y(_23338_));
 sky130_fd_sc_hd__nand2_4 _29816_ (.A(\count_instr[42] ),
    .B(\count_instr[43] ),
    .Y(_23339_));
 sky130_vsdinv _29817_ (.A(_23339_),
    .Y(_23340_));
 sky130_fd_sc_hd__and4_4 _29818_ (.A(_23313_),
    .B(\count_instr[40] ),
    .C(\count_instr[41] ),
    .D(_23340_),
    .X(_23341_));
 sky130_fd_sc_hd__nor4_4 _29819_ (.A(_19134_),
    .B(_23338_),
    .C(_21973_),
    .D(_19137_),
    .Y(_23342_));
 sky130_fd_sc_hd__a21o_4 _29820_ (.A1(_23341_),
    .A2(_23342_),
    .B1(_19977_),
    .X(_23343_));
 sky130_fd_sc_hd__a21oi_4 _29821_ (.A1(_23336_),
    .A2(_23338_),
    .B1(_23343_),
    .Y(_00106_));
 sky130_fd_sc_hd__buf_1 _29822_ (.A(\count_instr[45] ),
    .X(_23344_));
 sky130_fd_sc_hd__and2_4 _29823_ (.A(_23341_),
    .B(_23342_),
    .X(_23345_));
 sky130_fd_sc_hd__o21ai_4 _29824_ (.A1(_23344_),
    .A2(_23345_),
    .B1(_23175_),
    .Y(_23346_));
 sky130_fd_sc_hd__a21o_4 _29825_ (.A1(_23344_),
    .A2(_23345_),
    .B1(_23346_),
    .X(_23347_));
 sky130_vsdinv _29826_ (.A(_23347_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3_4 _29827_ (.A(_23313_),
    .B(_23308_),
    .C(_23317_),
    .X(_23348_));
 sky130_vsdinv _29828_ (.A(\count_instr[46] ),
    .Y(_23349_));
 sky130_fd_sc_hd__and4_4 _29829_ (.A(_23155_),
    .B(_23337_),
    .C(_23344_),
    .D(_23349_),
    .X(_23350_));
 sky130_fd_sc_hd__and4_4 _29830_ (.A(_23348_),
    .B(_23274_),
    .C(_23340_),
    .D(_23350_),
    .X(_23351_));
 sky130_fd_sc_hd__a41oi_4 _29831_ (.A1(_23344_),
    .A2(_23348_),
    .A3(_23340_),
    .A4(_23342_),
    .B1(_23349_),
    .Y(_23352_));
 sky130_fd_sc_hd__o21a_4 _29832_ (.A1(_23351_),
    .A2(_23352_),
    .B1(_23129_),
    .X(_00108_));
 sky130_fd_sc_hd__and4_4 _29833_ (.A(_23341_),
    .B(\count_instr[44] ),
    .C(\count_instr[45] ),
    .D(\count_instr[46] ),
    .X(_23353_));
 sky130_fd_sc_hd__buf_1 _29834_ (.A(\count_instr[47] ),
    .X(_23354_));
 sky130_fd_sc_hd__and3_4 _29835_ (.A(_23353_),
    .B(_23354_),
    .C(_23065_),
    .X(_23355_));
 sky130_vsdinv _29836_ (.A(_23355_),
    .Y(_23356_));
 sky130_fd_sc_hd__nand4_4 _29837_ (.A(_23337_),
    .B(_23341_),
    .C(\count_instr[45] ),
    .D(\count_instr[46] ),
    .Y(_23357_));
 sky130_fd_sc_hd__nor2_4 _29838_ (.A(_23002_),
    .B(_23357_),
    .Y(_23358_));
 sky130_fd_sc_hd__o21a_4 _29839_ (.A1(_23354_),
    .A2(_23358_),
    .B1(_23007_),
    .X(_23359_));
 sky130_fd_sc_hd__nand2_4 _29840_ (.A(_23356_),
    .B(_23359_),
    .Y(_23360_));
 sky130_vsdinv _29841_ (.A(_23360_),
    .Y(_00109_));
 sky130_fd_sc_hd__buf_1 _29842_ (.A(\count_instr[48] ),
    .X(_23361_));
 sky130_fd_sc_hd__buf_1 _29843_ (.A(_23353_),
    .X(_23362_));
 sky130_fd_sc_hd__buf_1 _29844_ (.A(_23354_),
    .X(_23363_));
 sky130_fd_sc_hd__and4_4 _29845_ (.A(_23362_),
    .B(_23111_),
    .C(_23363_),
    .D(_23021_),
    .X(_23364_));
 sky130_fd_sc_hd__buf_1 _29846_ (.A(_23354_),
    .X(_23365_));
 sky130_fd_sc_hd__buf_1 _29847_ (.A(_23362_),
    .X(_23366_));
 sky130_fd_sc_hd__a41oi_4 _29848_ (.A1(_23365_),
    .A2(_23366_),
    .A3(_23361_),
    .A4(_23165_),
    .B1(_23078_),
    .Y(_23367_));
 sky130_fd_sc_hd__o21a_4 _29849_ (.A1(_23361_),
    .A2(_23364_),
    .B1(_23367_),
    .X(_00110_));
 sky130_fd_sc_hd__and4_4 _29850_ (.A(_23362_),
    .B(_23363_),
    .C(_23361_),
    .D(_23006_),
    .X(_23368_));
 sky130_fd_sc_hd__nand2_4 _29851_ (.A(\count_instr[48] ),
    .B(\count_instr[49] ),
    .Y(_23369_));
 sky130_vsdinv _29852_ (.A(_23369_),
    .Y(_23370_));
 sky130_fd_sc_hd__buf_1 _29853_ (.A(_18786_),
    .X(_23371_));
 sky130_fd_sc_hd__buf_1 _29854_ (.A(_23371_),
    .X(_23372_));
 sky130_fd_sc_hd__a41oi_4 _29855_ (.A1(_23365_),
    .A2(_23366_),
    .A3(_23165_),
    .A4(_23370_),
    .B1(_23372_),
    .Y(_23373_));
 sky130_fd_sc_hd__o21a_4 _29856_ (.A1(\count_instr[49] ),
    .A2(_23368_),
    .B1(_23373_),
    .X(_00111_));
 sky130_fd_sc_hd__buf_1 _29857_ (.A(\count_instr[50] ),
    .X(_23374_));
 sky130_fd_sc_hd__nor4_4 _29858_ (.A(_19080_),
    .B(_23374_),
    .C(_23369_),
    .D(_23273_),
    .Y(_23375_));
 sky130_fd_sc_hd__and4_4 _29859_ (.A(_23362_),
    .B(_23022_),
    .C(_23363_),
    .D(_23375_),
    .X(_23376_));
 sky130_vsdinv _29860_ (.A(_23374_),
    .Y(_23377_));
 sky130_fd_sc_hd__a41oi_4 _29861_ (.A1(_23365_),
    .A2(_23366_),
    .A3(_23066_),
    .A4(_23370_),
    .B1(_23377_),
    .Y(_23378_));
 sky130_fd_sc_hd__buf_1 _29862_ (.A(_22929_),
    .X(_23379_));
 sky130_fd_sc_hd__o21a_4 _29863_ (.A1(_23376_),
    .A2(_23378_),
    .B1(_23379_),
    .X(_00113_));
 sky130_fd_sc_hd__nand4_4 _29864_ (.A(_23363_),
    .B(_23358_),
    .C(_23374_),
    .D(_23370_),
    .Y(_23380_));
 sky130_fd_sc_hd__nand2_4 _29865_ (.A(_23380_),
    .B(\count_instr[51] ),
    .Y(_23381_));
 sky130_fd_sc_hd__nor4_4 _29866_ (.A(_19091_),
    .B(_23377_),
    .C(\count_instr[51] ),
    .D(_23369_),
    .Y(_23382_));
 sky130_fd_sc_hd__nand4_4 _29867_ (.A(_23365_),
    .B(_23366_),
    .C(_18781_),
    .D(_23382_),
    .Y(_23383_));
 sky130_fd_sc_hd__a21oi_4 _29868_ (.A1(_23381_),
    .A2(_23383_),
    .B1(_23335_),
    .Y(_00114_));
 sky130_fd_sc_hd__buf_1 _29869_ (.A(\count_instr[52] ),
    .X(_23384_));
 sky130_fd_sc_hd__nand3_4 _29870_ (.A(\count_instr[49] ),
    .B(\count_instr[50] ),
    .C(\count_instr[51] ),
    .Y(_23385_));
 sky130_fd_sc_hd__nand3_4 _29871_ (.A(_23353_),
    .B(\count_instr[47] ),
    .C(\count_instr[48] ),
    .Y(_23386_));
 sky130_fd_sc_hd__nor3_4 _29872_ (.A(_23002_),
    .B(_23385_),
    .C(_23386_),
    .Y(_23387_));
 sky130_fd_sc_hd__o21a_4 _29873_ (.A1(_23384_),
    .A2(_23387_),
    .B1(_23263_),
    .X(_23388_));
 sky130_fd_sc_hd__nor2_4 _29874_ (.A(_23385_),
    .B(_23386_),
    .Y(_23389_));
 sky130_fd_sc_hd__buf_1 _29875_ (.A(_23389_),
    .X(_23390_));
 sky130_fd_sc_hd__buf_1 _29876_ (.A(_23390_),
    .X(_23391_));
 sky130_fd_sc_hd__nand3_4 _29877_ (.A(_23391_),
    .B(_23384_),
    .C(_23027_),
    .Y(_23392_));
 sky130_fd_sc_hd__nand2_4 _29878_ (.A(_23388_),
    .B(_23392_),
    .Y(_23393_));
 sky130_vsdinv _29879_ (.A(_23393_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand3_4 _29880_ (.A(_23390_),
    .B(_23384_),
    .C(_23085_),
    .Y(_23394_));
 sky130_vsdinv _29881_ (.A(\count_instr[53] ),
    .Y(_23395_));
 sky130_fd_sc_hd__nand2_4 _29882_ (.A(\count_instr[52] ),
    .B(\count_instr[53] ),
    .Y(_23396_));
 sky130_fd_sc_hd__nor4_4 _29883_ (.A(_23003_),
    .B(_23385_),
    .C(_23396_),
    .D(_23386_),
    .Y(_23397_));
 sky130_fd_sc_hd__a211o_4 _29884_ (.A1(_23394_),
    .A2(_23395_),
    .B1(_22992_),
    .C1(_23397_),
    .X(_23398_));
 sky130_vsdinv _29885_ (.A(_23398_),
    .Y(_00116_));
 sky130_fd_sc_hd__buf_1 _29886_ (.A(\count_instr[54] ),
    .X(_23399_));
 sky130_fd_sc_hd__o41ai_4 _29887_ (.A1(_23003_),
    .A2(_23385_),
    .A3(_23396_),
    .A4(_23386_),
    .B1(_23399_),
    .Y(_23400_));
 sky130_fd_sc_hd__nor4_4 _29888_ (.A(_23399_),
    .B(_23119_),
    .C(_23396_),
    .D(_23273_),
    .Y(_23401_));
 sky130_fd_sc_hd__nand2_4 _29889_ (.A(_23391_),
    .B(_23401_),
    .Y(_23402_));
 sky130_fd_sc_hd__a21oi_4 _29890_ (.A1(_23400_),
    .A2(_23402_),
    .B1(_23335_),
    .Y(_00117_));
 sky130_vsdinv _29891_ (.A(_23396_),
    .Y(_23403_));
 sky130_fd_sc_hd__a41o_4 _29892_ (.A1(_23391_),
    .A2(_23399_),
    .A3(_23085_),
    .A4(_23403_),
    .B1(\count_instr[55] ),
    .X(_23404_));
 sky130_fd_sc_hd__nand4_4 _29893_ (.A(_23399_),
    .B(_23387_),
    .C(\count_instr[55] ),
    .D(_23403_),
    .Y(_23405_));
 sky130_fd_sc_hd__and3_4 _29894_ (.A(_23404_),
    .B(_23405_),
    .C(_20932_),
    .X(_00118_));
 sky130_fd_sc_hd__buf_1 _29895_ (.A(\count_instr[56] ),
    .X(_23406_));
 sky130_fd_sc_hd__and4_4 _29896_ (.A(\count_instr[52] ),
    .B(\count_instr[53] ),
    .C(\count_instr[54] ),
    .D(\count_instr[55] ),
    .X(_23407_));
 sky130_fd_sc_hd__buf_1 _29897_ (.A(_23407_),
    .X(_23408_));
 sky130_fd_sc_hd__and3_4 _29898_ (.A(_23389_),
    .B(_23025_),
    .C(_23408_),
    .X(_23409_));
 sky130_fd_sc_hd__buf_1 _29899_ (.A(_23262_),
    .X(_23410_));
 sky130_fd_sc_hd__o21a_4 _29900_ (.A1(_23406_),
    .A2(_23409_),
    .B1(_23410_),
    .X(_23411_));
 sky130_fd_sc_hd__nand4_4 _29901_ (.A(_23406_),
    .B(_23390_),
    .C(_23085_),
    .D(_23408_),
    .Y(_23412_));
 sky130_fd_sc_hd__nand2_4 _29902_ (.A(_23411_),
    .B(_23412_),
    .Y(_23413_));
 sky130_vsdinv _29903_ (.A(_23413_),
    .Y(_00119_));
 sky130_fd_sc_hd__and3_4 _29904_ (.A(_23390_),
    .B(_23406_),
    .C(_23408_),
    .X(_23414_));
 sky130_fd_sc_hd__buf_1 _29905_ (.A(\count_instr[57] ),
    .X(_23415_));
 sky130_vsdinv _29906_ (.A(_23415_),
    .Y(_23416_));
 sky130_fd_sc_hd__nand3_4 _29907_ (.A(_23414_),
    .B(_23416_),
    .C(_23257_),
    .Y(_23417_));
 sky130_fd_sc_hd__nand2_4 _29908_ (.A(_23412_),
    .B(_23415_),
    .Y(_23418_));
 sky130_fd_sc_hd__a21oi_4 _29909_ (.A1(_23417_),
    .A2(_23418_),
    .B1(_23335_),
    .Y(_00120_));
 sky130_fd_sc_hd__buf_1 _29910_ (.A(\count_instr[58] ),
    .X(_23419_));
 sky130_fd_sc_hd__o21ai_4 _29911_ (.A1(_23416_),
    .A2(_23412_),
    .B1(_23419_),
    .Y(_23420_));
 sky130_vsdinv _29912_ (.A(_23419_),
    .Y(_23421_));
 sky130_fd_sc_hd__and4_4 _29913_ (.A(_23155_),
    .B(_23406_),
    .C(_23415_),
    .D(_23421_),
    .X(_23422_));
 sky130_fd_sc_hd__nand4_4 _29914_ (.A(_23275_),
    .B(_23391_),
    .C(_23408_),
    .D(_23422_),
    .Y(_23423_));
 sky130_fd_sc_hd__buf_1 _29915_ (.A(_19494_),
    .X(_23424_));
 sky130_fd_sc_hd__buf_1 _29916_ (.A(_23424_),
    .X(_23425_));
 sky130_fd_sc_hd__a21oi_4 _29917_ (.A1(_23420_),
    .A2(_23423_),
    .B1(_23425_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand3_4 _29918_ (.A(_23389_),
    .B(\count_instr[56] ),
    .C(_23407_),
    .Y(_23426_));
 sky130_fd_sc_hd__nor4_4 _29919_ (.A(_23416_),
    .B(_23421_),
    .C(_23003_),
    .D(_23426_),
    .Y(_23427_));
 sky130_fd_sc_hd__o21a_4 _29920_ (.A1(\count_instr[59] ),
    .A2(_23427_),
    .B1(_23410_),
    .X(_23428_));
 sky130_fd_sc_hd__and4_4 _29921_ (.A(_23389_),
    .B(\count_instr[56] ),
    .C(\count_instr[57] ),
    .D(_23407_),
    .X(_23429_));
 sky130_fd_sc_hd__buf_1 _29922_ (.A(_23429_),
    .X(_23430_));
 sky130_fd_sc_hd__nand4_4 _29923_ (.A(_23419_),
    .B(_23430_),
    .C(\count_instr[59] ),
    .D(_23006_),
    .Y(_23431_));
 sky130_fd_sc_hd__nand2_4 _29924_ (.A(_23428_),
    .B(_23431_),
    .Y(_23432_));
 sky130_vsdinv _29925_ (.A(_23432_),
    .Y(_00122_));
 sky130_vsdinv _29926_ (.A(\count_instr[60] ),
    .Y(_23433_));
 sky130_fd_sc_hd__buf_1 _29927_ (.A(\count_instr[60] ),
    .X(_23434_));
 sky130_fd_sc_hd__nand2_4 _29928_ (.A(\count_instr[58] ),
    .B(\count_instr[59] ),
    .Y(_23435_));
 sky130_vsdinv _29929_ (.A(_23435_),
    .Y(_23436_));
 sky130_fd_sc_hd__nand4_4 _29930_ (.A(_23434_),
    .B(_23430_),
    .C(_23006_),
    .D(_23436_),
    .Y(_23437_));
 sky130_fd_sc_hd__nand2_4 _29931_ (.A(_23437_),
    .B(_19126_),
    .Y(_23438_));
 sky130_fd_sc_hd__a21oi_4 _29932_ (.A1(_23431_),
    .A2(_23433_),
    .B1(_23438_),
    .Y(_00124_));
 sky130_fd_sc_hd__buf_1 _29933_ (.A(\count_instr[61] ),
    .X(_23439_));
 sky130_fd_sc_hd__nand3_4 _29934_ (.A(_23429_),
    .B(_23434_),
    .C(_23436_),
    .Y(_23440_));
 sky130_fd_sc_hd__or4_4 _29935_ (.A(_23439_),
    .B(_22425_),
    .C(_23012_),
    .D(_23440_),
    .X(_23441_));
 sky130_fd_sc_hd__nand2_4 _29936_ (.A(_23437_),
    .B(_23439_),
    .Y(_23442_));
 sky130_fd_sc_hd__a21oi_4 _29937_ (.A1(_23441_),
    .A2(_23442_),
    .B1(_23425_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand4_4 _29938_ (.A(_19120_),
    .B(_18778_),
    .C(\count_instr[61] ),
    .D(_21928_),
    .Y(_23443_));
 sky130_fd_sc_hd__nor2_4 _29939_ (.A(_22195_),
    .B(_23443_),
    .Y(_23444_));
 sky130_fd_sc_hd__nand4_4 _29940_ (.A(_23434_),
    .B(_23430_),
    .C(_23436_),
    .D(_23444_),
    .Y(_23445_));
 sky130_fd_sc_hd__nand2_4 _29941_ (.A(_23445_),
    .B(\count_instr[62] ),
    .Y(_23446_));
 sky130_vsdinv _29942_ (.A(\count_instr[62] ),
    .Y(_23447_));
 sky130_fd_sc_hd__and4_4 _29943_ (.A(_23155_),
    .B(_23434_),
    .C(_23439_),
    .D(_23447_),
    .X(_23448_));
 sky130_fd_sc_hd__nand4_4 _29944_ (.A(_23275_),
    .B(_23430_),
    .C(_23436_),
    .D(_23448_),
    .Y(_23449_));
 sky130_fd_sc_hd__a21oi_4 _29945_ (.A1(_23446_),
    .A2(_23449_),
    .B1(_23425_),
    .Y(_00126_));
 sky130_fd_sc_hd__nor4_4 _29946_ (.A(_23447_),
    .B(_22196_),
    .C(_23443_),
    .D(_23440_),
    .Y(_23450_));
 sky130_fd_sc_hd__nor4_4 _29947_ (.A(_23416_),
    .B(_23433_),
    .C(_23435_),
    .D(_23426_),
    .Y(_23451_));
 sky130_fd_sc_hd__a41oi_4 _29948_ (.A1(\count_instr[62] ),
    .A2(_23451_),
    .A3(\count_instr[63] ),
    .A4(_23444_),
    .B1(_18285_),
    .Y(_23452_));
 sky130_fd_sc_hd__o21ai_4 _29949_ (.A1(\count_instr[63] ),
    .A2(_23450_),
    .B1(_23452_),
    .Y(_23453_));
 sky130_vsdinv _29950_ (.A(_23453_),
    .Y(_00127_));
 sky130_fd_sc_hd__buf_1 _29951_ (.A(\irq_state[1] ),
    .X(_23454_));
 sky130_fd_sc_hd__nand3_4 _29952_ (.A(_18413_),
    .B(_18907_),
    .C(_23454_),
    .Y(_23455_));
 sky130_fd_sc_hd__nand2_4 _29953_ (.A(_19129_),
    .B(eoi[0]),
    .Y(_23456_));
 sky130_fd_sc_hd__a21o_4 _29954_ (.A1(_23455_),
    .A2(_23456_),
    .B1(_18579_),
    .X(_23457_));
 sky130_fd_sc_hd__nand2_4 _29955_ (.A(_21214_),
    .B(_19100_),
    .Y(_23458_));
 sky130_fd_sc_hd__buf_1 _29956_ (.A(_23458_),
    .X(_23459_));
 sky130_fd_sc_hd__buf_1 _29957_ (.A(_23459_),
    .X(_23460_));
 sky130_fd_sc_hd__nand2_4 _29958_ (.A(_19141_),
    .B(_20230_),
    .Y(_23461_));
 sky130_fd_sc_hd__buf_1 _29959_ (.A(_23461_),
    .X(_23462_));
 sky130_fd_sc_hd__buf_1 _29960_ (.A(_23462_),
    .X(_23463_));
 sky130_fd_sc_hd__nand3_4 _29961_ (.A(_23460_),
    .B(eoi[0]),
    .C(_23463_),
    .Y(_23464_));
 sky130_fd_sc_hd__a21oi_4 _29962_ (.A1(_23457_),
    .A2(_23464_),
    .B1(_23425_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand3_4 _29963_ (.A(_18410_),
    .B(_18935_),
    .C(_18903_),
    .Y(_23465_));
 sky130_fd_sc_hd__nand2_4 _29964_ (.A(_19129_),
    .B(eoi[1]),
    .Y(_23466_));
 sky130_fd_sc_hd__buf_1 _29965_ (.A(_18480_),
    .X(_23467_));
 sky130_fd_sc_hd__a21o_4 _29966_ (.A1(_23465_),
    .A2(_23466_),
    .B1(_23467_),
    .X(_23468_));
 sky130_fd_sc_hd__nand3_4 _29967_ (.A(_23460_),
    .B(eoi[1]),
    .C(_23463_),
    .Y(_23469_));
 sky130_fd_sc_hd__buf_1 _29968_ (.A(_23424_),
    .X(_23470_));
 sky130_fd_sc_hd__a21oi_4 _29969_ (.A1(_23468_),
    .A2(_23469_),
    .B1(_23470_),
    .Y(_00225_));
 sky130_fd_sc_hd__buf_1 _29970_ (.A(_23454_),
    .X(_23471_));
 sky130_fd_sc_hd__nand3_4 _29971_ (.A(_18416_),
    .B(_21991_),
    .C(_23471_),
    .Y(_23472_));
 sky130_fd_sc_hd__buf_1 _29972_ (.A(_23472_),
    .X(_23473_));
 sky130_fd_sc_hd__nand2_4 _29973_ (.A(_19129_),
    .B(eoi[2]),
    .Y(_23474_));
 sky130_fd_sc_hd__a21o_4 _29974_ (.A1(_23473_),
    .A2(_23474_),
    .B1(_23467_),
    .X(_23475_));
 sky130_fd_sc_hd__nand3_4 _29975_ (.A(_23460_),
    .B(eoi[2]),
    .C(_23463_),
    .Y(_23476_));
 sky130_fd_sc_hd__a21oi_4 _29976_ (.A1(_23475_),
    .A2(_23476_),
    .B1(_23470_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand3_4 _29977_ (.A(_18429_),
    .B(_18946_),
    .C(_18904_),
    .Y(_23477_));
 sky130_fd_sc_hd__buf_1 _29978_ (.A(_23477_),
    .X(_23478_));
 sky130_fd_sc_hd__buf_1 _29979_ (.A(_19128_),
    .X(_23479_));
 sky130_fd_sc_hd__buf_1 _29980_ (.A(_23479_),
    .X(_23480_));
 sky130_fd_sc_hd__nand2_4 _29981_ (.A(_23480_),
    .B(eoi[3]),
    .Y(_23481_));
 sky130_fd_sc_hd__a21o_4 _29982_ (.A1(_23478_),
    .A2(_23481_),
    .B1(_23467_),
    .X(_23482_));
 sky130_fd_sc_hd__buf_1 _29983_ (.A(_23462_),
    .X(_23483_));
 sky130_fd_sc_hd__nand3_4 _29984_ (.A(_23460_),
    .B(eoi[3]),
    .C(_23483_),
    .Y(_23484_));
 sky130_fd_sc_hd__a21oi_4 _29985_ (.A1(_23482_),
    .A2(_23484_),
    .B1(_23470_),
    .Y(_00239_));
 sky130_fd_sc_hd__buf_1 _29986_ (.A(_18903_),
    .X(_23485_));
 sky130_fd_sc_hd__nand3_4 _29987_ (.A(_18419_),
    .B(\irq_pending[4] ),
    .C(_23485_),
    .Y(_23486_));
 sky130_fd_sc_hd__buf_1 _29988_ (.A(_23486_),
    .X(_23487_));
 sky130_fd_sc_hd__buf_1 _29989_ (.A(_23487_),
    .X(_23488_));
 sky130_fd_sc_hd__nand2_4 _29990_ (.A(_23480_),
    .B(eoi[4]),
    .Y(_23489_));
 sky130_fd_sc_hd__a21o_4 _29991_ (.A1(_23488_),
    .A2(_23489_),
    .B1(_23467_),
    .X(_23490_));
 sky130_fd_sc_hd__buf_1 _29992_ (.A(_23459_),
    .X(_23491_));
 sky130_fd_sc_hd__nand3_4 _29993_ (.A(_23491_),
    .B(eoi[4]),
    .C(_23483_),
    .Y(_23492_));
 sky130_fd_sc_hd__a21oi_4 _29994_ (.A1(_23490_),
    .A2(_23492_),
    .B1(_23470_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand3_4 _29995_ (.A(_18432_),
    .B(\irq_pending[5] ),
    .C(_23485_),
    .Y(_23493_));
 sky130_fd_sc_hd__buf_1 _29996_ (.A(_23493_),
    .X(_23494_));
 sky130_fd_sc_hd__buf_1 _29997_ (.A(_23494_),
    .X(_23495_));
 sky130_fd_sc_hd__nand2_4 _29998_ (.A(_23480_),
    .B(eoi[5]),
    .Y(_23496_));
 sky130_fd_sc_hd__buf_1 _29999_ (.A(_18480_),
    .X(_23497_));
 sky130_fd_sc_hd__a21o_4 _30000_ (.A1(_23495_),
    .A2(_23496_),
    .B1(_23497_),
    .X(_23498_));
 sky130_fd_sc_hd__nand3_4 _30001_ (.A(_23491_),
    .B(eoi[5]),
    .C(_23483_),
    .Y(_23499_));
 sky130_fd_sc_hd__buf_1 _30002_ (.A(_23424_),
    .X(_23500_));
 sky130_fd_sc_hd__a21oi_4 _30003_ (.A1(_23498_),
    .A2(_23499_),
    .B1(_23500_),
    .Y(_00241_));
 sky130_fd_sc_hd__buf_1 _30004_ (.A(_23454_),
    .X(_23501_));
 sky130_fd_sc_hd__buf_1 _30005_ (.A(_23501_),
    .X(_23502_));
 sky130_fd_sc_hd__nand3_4 _30006_ (.A(_18414_),
    .B(\irq_pending[6] ),
    .C(_23502_),
    .Y(_23503_));
 sky130_fd_sc_hd__buf_1 _30007_ (.A(_23503_),
    .X(_23504_));
 sky130_fd_sc_hd__buf_1 _30008_ (.A(_23504_),
    .X(_23505_));
 sky130_fd_sc_hd__nand2_4 _30009_ (.A(_23480_),
    .B(eoi[6]),
    .Y(_23506_));
 sky130_fd_sc_hd__a21o_4 _30010_ (.A1(_23505_),
    .A2(_23506_),
    .B1(_23497_),
    .X(_23507_));
 sky130_fd_sc_hd__nand3_4 _30011_ (.A(_23491_),
    .B(eoi[6]),
    .C(_23483_),
    .Y(_23508_));
 sky130_fd_sc_hd__a21oi_4 _30012_ (.A1(_23507_),
    .A2(_23508_),
    .B1(_23500_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand3_4 _30013_ (.A(_18430_),
    .B(\irq_pending[7] ),
    .C(_23502_),
    .Y(_23509_));
 sky130_fd_sc_hd__buf_1 _30014_ (.A(_23509_),
    .X(_23510_));
 sky130_fd_sc_hd__buf_1 _30015_ (.A(_23510_),
    .X(_23511_));
 sky130_fd_sc_hd__buf_1 _30016_ (.A(_23479_),
    .X(_23512_));
 sky130_fd_sc_hd__nand2_4 _30017_ (.A(_23512_),
    .B(eoi[7]),
    .Y(_23513_));
 sky130_fd_sc_hd__a21o_4 _30018_ (.A1(_23511_),
    .A2(_23513_),
    .B1(_23497_),
    .X(_23514_));
 sky130_fd_sc_hd__buf_1 _30019_ (.A(_23461_),
    .X(_23515_));
 sky130_fd_sc_hd__buf_1 _30020_ (.A(_23515_),
    .X(_23516_));
 sky130_fd_sc_hd__nand3_4 _30021_ (.A(_23491_),
    .B(eoi[7]),
    .C(_23516_),
    .Y(_23517_));
 sky130_fd_sc_hd__a21oi_4 _30022_ (.A1(_23514_),
    .A2(_23517_),
    .B1(_23500_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand3_4 _30023_ (.A(_18436_),
    .B(\irq_pending[8] ),
    .C(_23502_),
    .Y(_23518_));
 sky130_fd_sc_hd__buf_1 _30024_ (.A(_23518_),
    .X(_23519_));
 sky130_fd_sc_hd__buf_1 _30025_ (.A(_23519_),
    .X(_23520_));
 sky130_fd_sc_hd__nand2_4 _30026_ (.A(_23512_),
    .B(eoi[8]),
    .Y(_23521_));
 sky130_fd_sc_hd__a21o_4 _30027_ (.A1(_23520_),
    .A2(_23521_),
    .B1(_23497_),
    .X(_23522_));
 sky130_fd_sc_hd__buf_1 _30028_ (.A(_23459_),
    .X(_23523_));
 sky130_fd_sc_hd__nand3_4 _30029_ (.A(_23523_),
    .B(eoi[8]),
    .C(_23516_),
    .Y(_23524_));
 sky130_fd_sc_hd__a21oi_4 _30030_ (.A1(_23522_),
    .A2(_23524_),
    .B1(_23500_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand3_4 _30031_ (.A(_18411_),
    .B(\irq_pending[9] ),
    .C(_23502_),
    .Y(_23525_));
 sky130_fd_sc_hd__buf_1 _30032_ (.A(_23525_),
    .X(_23526_));
 sky130_fd_sc_hd__buf_1 _30033_ (.A(_23526_),
    .X(_23527_));
 sky130_fd_sc_hd__nand2_4 _30034_ (.A(_23512_),
    .B(eoi[9]),
    .Y(_23528_));
 sky130_fd_sc_hd__buf_1 _30035_ (.A(_18479_),
    .X(_23529_));
 sky130_fd_sc_hd__buf_1 _30036_ (.A(_23529_),
    .X(_23530_));
 sky130_fd_sc_hd__a21o_4 _30037_ (.A1(_23527_),
    .A2(_23528_),
    .B1(_23530_),
    .X(_23531_));
 sky130_fd_sc_hd__nand3_4 _30038_ (.A(_23523_),
    .B(eoi[9]),
    .C(_23516_),
    .Y(_23532_));
 sky130_fd_sc_hd__buf_1 _30039_ (.A(_23424_),
    .X(_23533_));
 sky130_fd_sc_hd__a21oi_4 _30040_ (.A1(_23531_),
    .A2(_23532_),
    .B1(_23533_),
    .Y(_00245_));
 sky130_fd_sc_hd__buf_1 _30041_ (.A(_23501_),
    .X(_23534_));
 sky130_fd_sc_hd__nand3_4 _30042_ (.A(_18417_),
    .B(\irq_pending[10] ),
    .C(_23534_),
    .Y(_23535_));
 sky130_fd_sc_hd__buf_1 _30043_ (.A(_23535_),
    .X(_23536_));
 sky130_fd_sc_hd__buf_1 _30044_ (.A(_23536_),
    .X(_23537_));
 sky130_fd_sc_hd__nand2_4 _30045_ (.A(_23512_),
    .B(eoi[10]),
    .Y(_23538_));
 sky130_fd_sc_hd__a21o_4 _30046_ (.A1(_23537_),
    .A2(_23538_),
    .B1(_23530_),
    .X(_23539_));
 sky130_fd_sc_hd__nand3_4 _30047_ (.A(_23523_),
    .B(eoi[10]),
    .C(_23516_),
    .Y(_23540_));
 sky130_fd_sc_hd__a21oi_4 _30048_ (.A1(_23539_),
    .A2(_23540_),
    .B1(_23533_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand3_4 _30049_ (.A(_18439_),
    .B(\irq_pending[11] ),
    .C(_23534_),
    .Y(_23541_));
 sky130_fd_sc_hd__buf_1 _30050_ (.A(_23541_),
    .X(_23542_));
 sky130_fd_sc_hd__buf_1 _30051_ (.A(_23542_),
    .X(_23543_));
 sky130_fd_sc_hd__buf_1 _30052_ (.A(_23479_),
    .X(_23544_));
 sky130_fd_sc_hd__nand2_4 _30053_ (.A(_23544_),
    .B(eoi[11]),
    .Y(_23545_));
 sky130_fd_sc_hd__a21o_4 _30054_ (.A1(_23543_),
    .A2(_23545_),
    .B1(_23530_),
    .X(_23546_));
 sky130_fd_sc_hd__buf_1 _30055_ (.A(_23515_),
    .X(_23547_));
 sky130_fd_sc_hd__nand3_4 _30056_ (.A(_23523_),
    .B(eoi[11]),
    .C(_23547_),
    .Y(_23548_));
 sky130_fd_sc_hd__a21oi_4 _30057_ (.A1(_23546_),
    .A2(_23548_),
    .B1(_23533_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand3_4 _30058_ (.A(_18423_),
    .B(\irq_pending[12] ),
    .C(_23534_),
    .Y(_23549_));
 sky130_fd_sc_hd__buf_1 _30059_ (.A(_23549_),
    .X(_23550_));
 sky130_fd_sc_hd__buf_1 _30060_ (.A(_23550_),
    .X(_23551_));
 sky130_fd_sc_hd__nand2_4 _30061_ (.A(_23544_),
    .B(eoi[12]),
    .Y(_23552_));
 sky130_fd_sc_hd__a21o_4 _30062_ (.A1(_23551_),
    .A2(_23552_),
    .B1(_23530_),
    .X(_23553_));
 sky130_fd_sc_hd__buf_1 _30063_ (.A(_23459_),
    .X(_23554_));
 sky130_fd_sc_hd__nand3_4 _30064_ (.A(_23554_),
    .B(eoi[12]),
    .C(_23547_),
    .Y(_23555_));
 sky130_fd_sc_hd__a21oi_4 _30065_ (.A1(_23553_),
    .A2(_23555_),
    .B1(_23533_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand3_4 _30066_ (.A(_18445_),
    .B(\irq_pending[13] ),
    .C(_23534_),
    .Y(_23556_));
 sky130_fd_sc_hd__buf_1 _30067_ (.A(_23556_),
    .X(_23557_));
 sky130_fd_sc_hd__buf_1 _30068_ (.A(_23557_),
    .X(_23558_));
 sky130_fd_sc_hd__nand2_4 _30069_ (.A(_23544_),
    .B(eoi[13]),
    .Y(_23559_));
 sky130_fd_sc_hd__buf_1 _30070_ (.A(_23529_),
    .X(_23560_));
 sky130_fd_sc_hd__a21o_4 _30071_ (.A1(_23558_),
    .A2(_23559_),
    .B1(_23560_),
    .X(_23561_));
 sky130_fd_sc_hd__nand3_4 _30072_ (.A(_23554_),
    .B(eoi[13]),
    .C(_23547_),
    .Y(_23562_));
 sky130_fd_sc_hd__buf_1 _30073_ (.A(_19425_),
    .X(_23563_));
 sky130_fd_sc_hd__buf_1 _30074_ (.A(_23563_),
    .X(_23564_));
 sky130_fd_sc_hd__a21oi_4 _30075_ (.A1(_23561_),
    .A2(_23562_),
    .B1(_23564_),
    .Y(_00218_));
 sky130_fd_sc_hd__buf_1 _30076_ (.A(_23501_),
    .X(_23565_));
 sky130_fd_sc_hd__nand3_4 _30077_ (.A(_18437_),
    .B(\irq_pending[14] ),
    .C(_23565_),
    .Y(_23566_));
 sky130_fd_sc_hd__buf_1 _30078_ (.A(_23566_),
    .X(_23567_));
 sky130_fd_sc_hd__buf_1 _30079_ (.A(_23567_),
    .X(_23568_));
 sky130_fd_sc_hd__nand2_4 _30080_ (.A(_23544_),
    .B(eoi[14]),
    .Y(_23569_));
 sky130_fd_sc_hd__a21o_4 _30081_ (.A1(_23568_),
    .A2(_23569_),
    .B1(_23560_),
    .X(_23570_));
 sky130_fd_sc_hd__nand3_4 _30082_ (.A(_23554_),
    .B(eoi[14]),
    .C(_23547_),
    .Y(_23571_));
 sky130_fd_sc_hd__a21oi_4 _30083_ (.A1(_23570_),
    .A2(_23571_),
    .B1(_23564_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand3_4 _30084_ (.A(_18442_),
    .B(\irq_pending[15] ),
    .C(_23565_),
    .Y(_23572_));
 sky130_fd_sc_hd__buf_1 _30085_ (.A(_23572_),
    .X(_23573_));
 sky130_fd_sc_hd__buf_1 _30086_ (.A(_23573_),
    .X(_23574_));
 sky130_fd_sc_hd__buf_1 _30087_ (.A(_19128_),
    .X(_23575_));
 sky130_fd_sc_hd__buf_1 _30088_ (.A(_23575_),
    .X(_23576_));
 sky130_fd_sc_hd__nand2_4 _30089_ (.A(_23576_),
    .B(eoi[15]),
    .Y(_23577_));
 sky130_fd_sc_hd__a21o_4 _30090_ (.A1(_23574_),
    .A2(_23577_),
    .B1(_23560_),
    .X(_23578_));
 sky130_fd_sc_hd__buf_1 _30091_ (.A(_23515_),
    .X(_23579_));
 sky130_fd_sc_hd__nand3_4 _30092_ (.A(_23554_),
    .B(eoi[15]),
    .C(_23579_),
    .Y(_23580_));
 sky130_fd_sc_hd__a21oi_4 _30093_ (.A1(_23578_),
    .A2(_23580_),
    .B1(_23564_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand3_4 _30094_ (.A(_18433_),
    .B(\irq_pending[16] ),
    .C(_23565_),
    .Y(_23581_));
 sky130_fd_sc_hd__buf_1 _30095_ (.A(_23581_),
    .X(_23582_));
 sky130_fd_sc_hd__buf_1 _30096_ (.A(_23582_),
    .X(_23583_));
 sky130_fd_sc_hd__nand2_4 _30097_ (.A(_23576_),
    .B(eoi[16]),
    .Y(_23584_));
 sky130_fd_sc_hd__a21o_4 _30098_ (.A1(_23583_),
    .A2(_23584_),
    .B1(_23560_),
    .X(_23585_));
 sky130_fd_sc_hd__buf_1 _30099_ (.A(_23458_),
    .X(_23586_));
 sky130_fd_sc_hd__buf_1 _30100_ (.A(_23586_),
    .X(_23587_));
 sky130_fd_sc_hd__nand3_4 _30101_ (.A(_23587_),
    .B(eoi[16]),
    .C(_23579_),
    .Y(_23588_));
 sky130_fd_sc_hd__a21oi_4 _30102_ (.A1(_23585_),
    .A2(_23588_),
    .B1(_23564_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand3_4 _30103_ (.A(_18449_),
    .B(\irq_pending[17] ),
    .C(_23565_),
    .Y(_23589_));
 sky130_fd_sc_hd__buf_1 _30104_ (.A(_23589_),
    .X(_23590_));
 sky130_fd_sc_hd__buf_1 _30105_ (.A(_23590_),
    .X(_23591_));
 sky130_fd_sc_hd__nand2_4 _30106_ (.A(_23576_),
    .B(eoi[17]),
    .Y(_23592_));
 sky130_fd_sc_hd__buf_1 _30107_ (.A(_23529_),
    .X(_23593_));
 sky130_fd_sc_hd__a21o_4 _30108_ (.A1(_23591_),
    .A2(_23592_),
    .B1(_23593_),
    .X(_23594_));
 sky130_fd_sc_hd__nand3_4 _30109_ (.A(_23587_),
    .B(eoi[17]),
    .C(_23579_),
    .Y(_23595_));
 sky130_fd_sc_hd__buf_1 _30110_ (.A(_23563_),
    .X(_23596_));
 sky130_fd_sc_hd__a21oi_4 _30111_ (.A1(_23594_),
    .A2(_23595_),
    .B1(_23596_),
    .Y(_00222_));
 sky130_fd_sc_hd__buf_1 _30112_ (.A(_18903_),
    .X(_23597_));
 sky130_fd_sc_hd__nand3_4 _30113_ (.A(_18450_),
    .B(\irq_pending[18] ),
    .C(_23597_),
    .Y(_23598_));
 sky130_fd_sc_hd__buf_1 _30114_ (.A(_23598_),
    .X(_23599_));
 sky130_fd_sc_hd__nand2_4 _30115_ (.A(_23576_),
    .B(eoi[18]),
    .Y(_23600_));
 sky130_fd_sc_hd__a21o_4 _30116_ (.A1(_23599_),
    .A2(_23600_),
    .B1(_23593_),
    .X(_23601_));
 sky130_fd_sc_hd__nand3_4 _30117_ (.A(_23587_),
    .B(eoi[18]),
    .C(_23579_),
    .Y(_23602_));
 sky130_fd_sc_hd__a21oi_4 _30118_ (.A1(_23601_),
    .A2(_23602_),
    .B1(_23596_),
    .Y(_00223_));
 sky130_fd_sc_hd__buf_1 _30119_ (.A(_23501_),
    .X(_23603_));
 sky130_fd_sc_hd__nand3_4 _30120_ (.A(_18426_),
    .B(\irq_pending[19] ),
    .C(_23603_),
    .Y(_23604_));
 sky130_fd_sc_hd__buf_1 _30121_ (.A(_23604_),
    .X(_23605_));
 sky130_fd_sc_hd__buf_1 _30122_ (.A(_23605_),
    .X(_23606_));
 sky130_fd_sc_hd__buf_1 _30123_ (.A(_23575_),
    .X(_23607_));
 sky130_fd_sc_hd__nand2_4 _30124_ (.A(_23607_),
    .B(eoi[19]),
    .Y(_23608_));
 sky130_fd_sc_hd__a21o_4 _30125_ (.A1(_23606_),
    .A2(_23608_),
    .B1(_23593_),
    .X(_23609_));
 sky130_fd_sc_hd__buf_1 _30126_ (.A(_23515_),
    .X(_23610_));
 sky130_fd_sc_hd__nand3_4 _30127_ (.A(_23587_),
    .B(eoi[19]),
    .C(_23610_),
    .Y(_23611_));
 sky130_fd_sc_hd__a21oi_4 _30128_ (.A1(_23609_),
    .A2(_23611_),
    .B1(_23596_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand3_4 _30129_ (.A(_18440_),
    .B(\irq_pending[20] ),
    .C(_23603_),
    .Y(_23612_));
 sky130_fd_sc_hd__buf_1 _30130_ (.A(_23612_),
    .X(_23613_));
 sky130_fd_sc_hd__buf_1 _30131_ (.A(_23613_),
    .X(_23614_));
 sky130_fd_sc_hd__nand2_4 _30132_ (.A(_23607_),
    .B(eoi[20]),
    .Y(_23615_));
 sky130_fd_sc_hd__a21o_4 _30133_ (.A1(_23614_),
    .A2(_23615_),
    .B1(_23593_),
    .X(_23616_));
 sky130_fd_sc_hd__buf_1 _30134_ (.A(_23586_),
    .X(_23617_));
 sky130_fd_sc_hd__nand3_4 _30135_ (.A(_23617_),
    .B(eoi[20]),
    .C(_23610_),
    .Y(_23618_));
 sky130_fd_sc_hd__a21oi_4 _30136_ (.A1(_23616_),
    .A2(_23618_),
    .B1(_23596_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand3_4 _30137_ (.A(_18443_),
    .B(\irq_pending[21] ),
    .C(_23603_),
    .Y(_23619_));
 sky130_fd_sc_hd__buf_1 _30138_ (.A(_23619_),
    .X(_23620_));
 sky130_fd_sc_hd__buf_1 _30139_ (.A(_23620_),
    .X(_23621_));
 sky130_fd_sc_hd__nand2_4 _30140_ (.A(_23607_),
    .B(eoi[21]),
    .Y(_23622_));
 sky130_fd_sc_hd__buf_1 _30141_ (.A(_23529_),
    .X(_23623_));
 sky130_fd_sc_hd__a21o_4 _30142_ (.A1(_23621_),
    .A2(_23622_),
    .B1(_23623_),
    .X(_23624_));
 sky130_fd_sc_hd__nand3_4 _30143_ (.A(_23617_),
    .B(eoi[21]),
    .C(_23610_),
    .Y(_23625_));
 sky130_fd_sc_hd__buf_1 _30144_ (.A(_23563_),
    .X(_23626_));
 sky130_fd_sc_hd__a21oi_4 _30145_ (.A1(_23624_),
    .A2(_23625_),
    .B1(_23626_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand3_4 _30146_ (.A(_18427_),
    .B(\irq_pending[22] ),
    .C(_23597_),
    .Y(_23627_));
 sky130_fd_sc_hd__buf_1 _30147_ (.A(_23627_),
    .X(_23628_));
 sky130_fd_sc_hd__nand2_4 _30148_ (.A(_23607_),
    .B(eoi[22]),
    .Y(_23629_));
 sky130_fd_sc_hd__a21o_4 _30149_ (.A1(_23628_),
    .A2(_23629_),
    .B1(_23623_),
    .X(_23630_));
 sky130_fd_sc_hd__nand3_4 _30150_ (.A(_23617_),
    .B(eoi[22]),
    .C(_23610_),
    .Y(_23631_));
 sky130_fd_sc_hd__a21oi_4 _30151_ (.A1(_23630_),
    .A2(_23631_),
    .B1(_23626_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand3_4 _30152_ (.A(_18424_),
    .B(\irq_pending[23] ),
    .C(_23603_),
    .Y(_23632_));
 sky130_fd_sc_hd__buf_1 _30153_ (.A(_23632_),
    .X(_23633_));
 sky130_fd_sc_hd__buf_1 _30154_ (.A(_23633_),
    .X(_23634_));
 sky130_fd_sc_hd__buf_1 _30155_ (.A(_23575_),
    .X(_23635_));
 sky130_fd_sc_hd__nand2_4 _30156_ (.A(_23635_),
    .B(eoi[23]),
    .Y(_23636_));
 sky130_fd_sc_hd__a21o_4 _30157_ (.A1(_23634_),
    .A2(_23636_),
    .B1(_23623_),
    .X(_23637_));
 sky130_fd_sc_hd__buf_1 _30158_ (.A(_23461_),
    .X(_23638_));
 sky130_fd_sc_hd__nand3_4 _30159_ (.A(_23617_),
    .B(eoi[23]),
    .C(_23638_),
    .Y(_23639_));
 sky130_fd_sc_hd__a21oi_4 _30160_ (.A1(_23637_),
    .A2(_23639_),
    .B1(_23626_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand3_4 _30161_ (.A(_18458_),
    .B(\irq_pending[24] ),
    .C(_23471_),
    .Y(_23640_));
 sky130_fd_sc_hd__buf_1 _30162_ (.A(_23640_),
    .X(_23641_));
 sky130_fd_sc_hd__buf_1 _30163_ (.A(_23641_),
    .X(_23642_));
 sky130_fd_sc_hd__nand2_4 _30164_ (.A(_23635_),
    .B(eoi[24]),
    .Y(_23643_));
 sky130_fd_sc_hd__a21o_4 _30165_ (.A1(_23642_),
    .A2(_23643_),
    .B1(_23623_),
    .X(_23644_));
 sky130_fd_sc_hd__buf_1 _30166_ (.A(_23586_),
    .X(_23645_));
 sky130_fd_sc_hd__nand3_4 _30167_ (.A(_23645_),
    .B(eoi[24]),
    .C(_23638_),
    .Y(_23646_));
 sky130_fd_sc_hd__a21oi_4 _30168_ (.A1(_23644_),
    .A2(_23646_),
    .B1(_23626_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand3_4 _30169_ (.A(_18452_),
    .B(\irq_pending[25] ),
    .C(_23471_),
    .Y(_23647_));
 sky130_fd_sc_hd__buf_1 _30170_ (.A(_23647_),
    .X(_23648_));
 sky130_fd_sc_hd__buf_1 _30171_ (.A(_23648_),
    .X(_23649_));
 sky130_fd_sc_hd__nand2_4 _30172_ (.A(_23635_),
    .B(eoi[25]),
    .Y(_23650_));
 sky130_fd_sc_hd__buf_1 _30173_ (.A(_19080_),
    .X(_23651_));
 sky130_fd_sc_hd__a21o_4 _30174_ (.A1(_23649_),
    .A2(_23650_),
    .B1(_23651_),
    .X(_23652_));
 sky130_fd_sc_hd__nand3_4 _30175_ (.A(_23645_),
    .B(eoi[25]),
    .C(_23638_),
    .Y(_23653_));
 sky130_fd_sc_hd__buf_1 _30176_ (.A(_23563_),
    .X(_23654_));
 sky130_fd_sc_hd__a21oi_4 _30177_ (.A1(_23652_),
    .A2(_23653_),
    .B1(_23654_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand3_4 _30178_ (.A(_18453_),
    .B(\irq_pending[26] ),
    .C(_23471_),
    .Y(_23655_));
 sky130_fd_sc_hd__buf_1 _30179_ (.A(_23655_),
    .X(_23656_));
 sky130_fd_sc_hd__buf_1 _30180_ (.A(_23656_),
    .X(_23657_));
 sky130_fd_sc_hd__nand2_4 _30181_ (.A(_23635_),
    .B(eoi[26]),
    .Y(_23658_));
 sky130_fd_sc_hd__a21o_4 _30182_ (.A1(_23657_),
    .A2(_23658_),
    .B1(_23651_),
    .X(_23659_));
 sky130_fd_sc_hd__nand3_4 _30183_ (.A(_23645_),
    .B(eoi[26]),
    .C(_23638_),
    .Y(_23660_));
 sky130_fd_sc_hd__a21oi_4 _30184_ (.A1(_23659_),
    .A2(_23660_),
    .B1(_23654_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand3_4 _30185_ (.A(_18455_),
    .B(\irq_pending[27] ),
    .C(_23597_),
    .Y(_23661_));
 sky130_fd_sc_hd__buf_1 _30186_ (.A(_23661_),
    .X(_23662_));
 sky130_fd_sc_hd__buf_1 _30187_ (.A(_23575_),
    .X(_23663_));
 sky130_fd_sc_hd__nand2_4 _30188_ (.A(_23663_),
    .B(eoi[27]),
    .Y(_23664_));
 sky130_fd_sc_hd__a21o_4 _30189_ (.A1(_23662_),
    .A2(_23664_),
    .B1(_23651_),
    .X(_23665_));
 sky130_fd_sc_hd__buf_1 _30190_ (.A(_23461_),
    .X(_23666_));
 sky130_fd_sc_hd__nand3_4 _30191_ (.A(_23645_),
    .B(eoi[27]),
    .C(_23666_),
    .Y(_23667_));
 sky130_fd_sc_hd__a21oi_4 _30192_ (.A1(_23665_),
    .A2(_23667_),
    .B1(_23654_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand3_4 _30193_ (.A(_18446_),
    .B(\irq_pending[28] ),
    .C(_23454_),
    .Y(_23668_));
 sky130_fd_sc_hd__nand2_4 _30194_ (.A(_23663_),
    .B(eoi[28]),
    .Y(_23669_));
 sky130_fd_sc_hd__a21o_4 _30195_ (.A1(_23668_),
    .A2(_23669_),
    .B1(_23651_),
    .X(_23670_));
 sky130_fd_sc_hd__buf_1 _30196_ (.A(_23586_),
    .X(_23671_));
 sky130_fd_sc_hd__nand3_4 _30197_ (.A(_23671_),
    .B(eoi[28]),
    .C(_23666_),
    .Y(_23672_));
 sky130_fd_sc_hd__a21oi_4 _30198_ (.A1(_23670_),
    .A2(_23672_),
    .B1(_23654_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand3_4 _30199_ (.A(_18420_),
    .B(\irq_pending[29] ),
    .C(_23597_),
    .Y(_23673_));
 sky130_fd_sc_hd__buf_1 _30200_ (.A(_23673_),
    .X(_23674_));
 sky130_fd_sc_hd__nand2_4 _30201_ (.A(_23663_),
    .B(eoi[29]),
    .Y(_23675_));
 sky130_fd_sc_hd__a21o_4 _30202_ (.A1(_23674_),
    .A2(_23675_),
    .B1(_19081_),
    .X(_23676_));
 sky130_fd_sc_hd__nand3_4 _30203_ (.A(_23671_),
    .B(eoi[29]),
    .C(_23666_),
    .Y(_23677_));
 sky130_fd_sc_hd__buf_1 _30204_ (.A(_19425_),
    .X(_23678_));
 sky130_fd_sc_hd__buf_1 _30205_ (.A(_23678_),
    .X(_23679_));
 sky130_fd_sc_hd__a21oi_4 _30206_ (.A1(_23676_),
    .A2(_23677_),
    .B1(_23679_),
    .Y(_00235_));
 sky130_fd_sc_hd__nand3_4 _30207_ (.A(_18456_),
    .B(\irq_pending[30] ),
    .C(_23485_),
    .Y(_23680_));
 sky130_fd_sc_hd__buf_1 _30208_ (.A(_23680_),
    .X(_23681_));
 sky130_fd_sc_hd__nand2_4 _30209_ (.A(_23663_),
    .B(eoi[30]),
    .Y(_23682_));
 sky130_fd_sc_hd__a21o_4 _30210_ (.A1(_23681_),
    .A2(_23682_),
    .B1(_19081_),
    .X(_23683_));
 sky130_fd_sc_hd__nand3_4 _30211_ (.A(_23671_),
    .B(eoi[30]),
    .C(_23666_),
    .Y(_23684_));
 sky130_fd_sc_hd__a21oi_4 _30212_ (.A1(_23683_),
    .A2(_23684_),
    .B1(_23679_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand3_4 _30213_ (.A(_18459_),
    .B(\irq_pending[31] ),
    .C(_23485_),
    .Y(_23685_));
 sky130_fd_sc_hd__buf_1 _30214_ (.A(_23685_),
    .X(_23686_));
 sky130_fd_sc_hd__nand2_4 _30215_ (.A(_23479_),
    .B(eoi[31]),
    .Y(_23687_));
 sky130_fd_sc_hd__a21o_4 _30216_ (.A1(_23686_),
    .A2(_23687_),
    .B1(_19081_),
    .X(_23688_));
 sky130_fd_sc_hd__nand3_4 _30217_ (.A(_23671_),
    .B(eoi[31]),
    .C(_23462_),
    .Y(_23689_));
 sky130_fd_sc_hd__a21oi_4 _30218_ (.A1(_23688_),
    .A2(_23689_),
    .B1(_23679_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand3_4 _30219_ (.A(mem_rdata[19]),
    .B(_18872_),
    .C(_18873_),
    .Y(_23690_));
 sky130_fd_sc_hd__a21bo_4 _30220_ (.A1(\mem_rdata_q[19] ),
    .A2(_18199_),
    .B1_N(_23690_),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__buf_1 _30221_ (.A(_19049_),
    .X(_23691_));
 sky130_fd_sc_hd__buf_1 _30222_ (.A(_18360_),
    .X(_23692_));
 sky130_fd_sc_hd__buf_1 _30223_ (.A(_18892_),
    .X(_23693_));
 sky130_fd_sc_hd__buf_1 _30224_ (.A(_23693_),
    .X(_23694_));
 sky130_fd_sc_hd__buf_1 _30225_ (.A(_23694_),
    .X(_23695_));
 sky130_fd_sc_hd__and4_4 _30226_ (.A(_23692_),
    .B(_23096_),
    .C(_23695_),
    .D(\mem_rdata_latched[19] ),
    .X(_23696_));
 sky130_fd_sc_hd__nand2_4 _30227_ (.A(\mem_rdata_latched[3] ),
    .B(_18197_),
    .Y(_23697_));
 sky130_fd_sc_hd__and2_4 _30228_ (.A(\mem_rdata_latched[1] ),
    .B(\mem_rdata_latched[0] ),
    .X(_23698_));
 sky130_vsdinv _30229_ (.A(_23698_),
    .Y(_23699_));
 sky130_fd_sc_hd__nor4_4 _30230_ (.A(\mem_rdata_latched[25] ),
    .B(\mem_rdata_latched[28] ),
    .C(_23697_),
    .D(_23699_),
    .Y(_23700_));
 sky130_fd_sc_hd__and3_4 _30231_ (.A(_18214_),
    .B(_18217_),
    .C(_18221_),
    .X(_23701_));
 sky130_fd_sc_hd__and4_4 _30232_ (.A(_23701_),
    .B(_18881_),
    .C(_18883_),
    .D(_18885_),
    .X(_23702_));
 sky130_fd_sc_hd__buf_1 _30233_ (.A(_23702_),
    .X(_23703_));
 sky130_fd_sc_hd__nand4_4 _30234_ (.A(_18209_),
    .B(_23700_),
    .C(_23703_),
    .D(_19050_),
    .Y(_23704_));
 sky130_vsdinv _30235_ (.A(_23704_),
    .Y(_23705_));
 sky130_fd_sc_hd__a211o_4 _30236_ (.A1(\decoded_rs1[4] ),
    .A2(_23691_),
    .B1(_23696_),
    .C1(_23705_),
    .X(_00205_));
 sky130_fd_sc_hd__buf_1 _30237_ (.A(_19050_),
    .X(_23706_));
 sky130_fd_sc_hd__buf_1 _30238_ (.A(_23706_),
    .X(_23707_));
 sky130_fd_sc_hd__buf_1 _30239_ (.A(_18360_),
    .X(_23708_));
 sky130_fd_sc_hd__buf_1 _30240_ (.A(_23708_),
    .X(_23709_));
 sky130_fd_sc_hd__buf_1 _30241_ (.A(_23693_),
    .X(_23710_));
 sky130_fd_sc_hd__buf_1 _30242_ (.A(_23710_),
    .X(_23711_));
 sky130_fd_sc_hd__buf_1 _30243_ (.A(_23711_),
    .X(_23712_));
 sky130_fd_sc_hd__buf_1 _30244_ (.A(_23712_),
    .X(_23713_));
 sky130_fd_sc_hd__nand4_4 _30245_ (.A(_22981_),
    .B(_23709_),
    .C(_23713_),
    .D(\mem_rdata_latched[30] ),
    .Y(_23714_));
 sky130_fd_sc_hd__o21ai_4 _30246_ (.A1(_22335_),
    .A2(_23707_),
    .B1(_23714_),
    .Y(_00165_));
 sky130_fd_sc_hd__buf_1 _30247_ (.A(_19049_),
    .X(_23715_));
 sky130_fd_sc_hd__buf_1 _30248_ (.A(_23715_),
    .X(_23716_));
 sky130_fd_sc_hd__buf_1 _30249_ (.A(_18359_),
    .X(_23717_));
 sky130_fd_sc_hd__and4_4 _30250_ (.A(_23717_),
    .B(_18835_),
    .C(_23695_),
    .D(\mem_rdata_latched[27] ),
    .X(_23718_));
 sky130_fd_sc_hd__a21o_4 _30251_ (.A1(\decoded_imm_uj[7] ),
    .A2(_23716_),
    .B1(_23718_),
    .X(_00193_));
 sky130_fd_sc_hd__buf_1 _30252_ (.A(_19124_),
    .X(_23719_));
 sky130_fd_sc_hd__buf_1 _30253_ (.A(_23719_),
    .X(_23720_));
 sky130_fd_sc_hd__nand4_4 _30254_ (.A(_23720_),
    .B(_23709_),
    .C(_23713_),
    .D(\mem_rdata_latched[26] ),
    .Y(_23721_));
 sky130_fd_sc_hd__o21ai_4 _30255_ (.A1(_22198_),
    .A2(_23707_),
    .B1(_23721_),
    .Y(_00192_));
 sky130_vsdinv _30256_ (.A(\mem_rdata_q[21] ),
    .Y(_23722_));
 sky130_fd_sc_hd__buf_1 _30257_ (.A(_18871_),
    .X(_23723_));
 sky130_fd_sc_hd__buf_1 _30258_ (.A(_18200_),
    .X(_23724_));
 sky130_fd_sc_hd__buf_1 _30259_ (.A(_18201_),
    .X(_23725_));
 sky130_fd_sc_hd__nand3_4 _30260_ (.A(mem_rdata[21]),
    .B(_23724_),
    .C(_23725_),
    .Y(_23726_));
 sky130_fd_sc_hd__o21ai_4 _30261_ (.A1(_23722_),
    .A2(_23723_),
    .B1(_23726_),
    .Y(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__buf_1 _30262_ (.A(_23691_),
    .X(_23727_));
 sky130_fd_sc_hd__buf_1 _30263_ (.A(_23717_),
    .X(_23728_));
 sky130_fd_sc_hd__buf_1 _30264_ (.A(_23694_),
    .X(_23729_));
 sky130_fd_sc_hd__buf_1 _30265_ (.A(_23729_),
    .X(_23730_));
 sky130_fd_sc_hd__nand4_4 _30266_ (.A(_18843_),
    .B(_23728_),
    .C(_23730_),
    .D(\mem_rdata_latched[21] ),
    .Y(_23731_));
 sky130_fd_sc_hd__a21bo_4 _30267_ (.A1(\decoded_imm_uj[1] ),
    .A2(_23727_),
    .B1_N(_23731_),
    .X(_00175_));
 sky130_fd_sc_hd__buf_1 _30268_ (.A(\mem_rdata_q[22] ),
    .X(_23732_));
 sky130_fd_sc_hd__buf_1 _30269_ (.A(_18199_),
    .X(_23733_));
 sky130_fd_sc_hd__buf_1 _30270_ (.A(_18206_),
    .X(_23734_));
 sky130_fd_sc_hd__buf_1 _30271_ (.A(_23734_),
    .X(_23735_));
 sky130_fd_sc_hd__buf_1 _30272_ (.A(_18207_),
    .X(_23736_));
 sky130_fd_sc_hd__buf_1 _30273_ (.A(_23736_),
    .X(_23737_));
 sky130_fd_sc_hd__nand3_4 _30274_ (.A(mem_rdata[22]),
    .B(_23735_),
    .C(_23737_),
    .Y(_23738_));
 sky130_fd_sc_hd__a21bo_4 _30275_ (.A1(_23732_),
    .A2(_23733_),
    .B1_N(_23738_),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__buf_1 _30276_ (.A(_23096_),
    .X(_23739_));
 sky130_fd_sc_hd__buf_1 _30277_ (.A(_23695_),
    .X(_23740_));
 sky130_fd_sc_hd__nand4_4 _30278_ (.A(_23739_),
    .B(_23728_),
    .C(_23740_),
    .D(\mem_rdata_latched[22] ),
    .Y(_23741_));
 sky130_fd_sc_hd__o21ai_4 _30279_ (.A1(_21976_),
    .A2(_23707_),
    .B1(_23741_),
    .Y(_00186_));
 sky130_fd_sc_hd__buf_1 _30280_ (.A(\mem_rdata_q[23] ),
    .X(_23742_));
 sky130_fd_sc_hd__nand3_4 _30281_ (.A(mem_rdata[23]),
    .B(_23735_),
    .C(_23737_),
    .Y(_23743_));
 sky130_fd_sc_hd__a21bo_4 _30282_ (.A1(_23742_),
    .A2(_23733_),
    .B1_N(_23743_),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__nand4_4 _30283_ (.A(_23739_),
    .B(_23728_),
    .C(_23730_),
    .D(\mem_rdata_latched[23] ),
    .Y(_23744_));
 sky130_fd_sc_hd__o21ai_4 _30284_ (.A1(_22051_),
    .A2(_23707_),
    .B1(_23744_),
    .Y(_00189_));
 sky130_fd_sc_hd__buf_1 _30285_ (.A(_19050_),
    .X(_23745_));
 sky130_fd_sc_hd__buf_1 _30286_ (.A(_23745_),
    .X(_23746_));
 sky130_fd_sc_hd__nand4_4 _30287_ (.A(_23720_),
    .B(_23709_),
    .C(_23713_),
    .D(\mem_rdata_latched[25] ),
    .Y(_23747_));
 sky130_fd_sc_hd__o21ai_4 _30288_ (.A1(_22138_),
    .A2(_23746_),
    .B1(_23747_),
    .Y(_00191_));
 sky130_fd_sc_hd__buf_1 _30289_ (.A(_23692_),
    .X(_23748_));
 sky130_fd_sc_hd__nand4_4 _30290_ (.A(_23720_),
    .B(_23748_),
    .C(_23713_),
    .D(\mem_rdata_latched[28] ),
    .Y(_23749_));
 sky130_fd_sc_hd__o21ai_4 _30291_ (.A1(_22230_),
    .A2(_23746_),
    .B1(_23749_),
    .Y(_00194_));
 sky130_fd_sc_hd__buf_1 _30292_ (.A(_23712_),
    .X(_23750_));
 sky130_fd_sc_hd__nand4_4 _30293_ (.A(_23720_),
    .B(_23748_),
    .C(_23750_),
    .D(\mem_rdata_latched[29] ),
    .Y(_23751_));
 sky130_fd_sc_hd__o21ai_4 _30294_ (.A1(_22298_),
    .A2(_23746_),
    .B1(_23751_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand4_4 _30295_ (.A(_18835_),
    .B(_23717_),
    .C(_23729_),
    .D(\mem_rdata_latched[31] ),
    .Y(_23752_));
 sky130_fd_sc_hd__buf_1 _30296_ (.A(_23752_),
    .X(_23753_));
 sky130_fd_sc_hd__o21ai_4 _30297_ (.A1(_22588_),
    .A2(_23746_),
    .B1(_23753_),
    .Y(_00176_));
 sky130_fd_sc_hd__buf_1 _30298_ (.A(_23745_),
    .X(_23754_));
 sky130_fd_sc_hd__o21ai_4 _30299_ (.A1(_22657_),
    .A2(_23754_),
    .B1(_23753_),
    .Y(_00177_));
 sky130_fd_sc_hd__o21ai_4 _30300_ (.A1(_22649_),
    .A2(_23754_),
    .B1(_23753_),
    .Y(_00178_));
 sky130_fd_sc_hd__o21ai_4 _30301_ (.A1(_22712_),
    .A2(_23754_),
    .B1(_23753_),
    .Y(_00179_));
 sky130_fd_sc_hd__buf_1 _30302_ (.A(_23752_),
    .X(_23755_));
 sky130_fd_sc_hd__o21ai_4 _30303_ (.A1(_22709_),
    .A2(_23754_),
    .B1(_23755_),
    .Y(_00180_));
 sky130_fd_sc_hd__buf_1 _30304_ (.A(_23745_),
    .X(_23756_));
 sky130_fd_sc_hd__o21ai_4 _30305_ (.A1(_22739_),
    .A2(_23756_),
    .B1(_23755_),
    .Y(_00181_));
 sky130_fd_sc_hd__o21ai_4 _30306_ (.A1(_22793_),
    .A2(_23756_),
    .B1(_23755_),
    .Y(_00182_));
 sky130_fd_sc_hd__o21ai_4 _30307_ (.A1(_22830_),
    .A2(_23756_),
    .B1(_23755_),
    .Y(_00183_));
 sky130_fd_sc_hd__buf_1 _30308_ (.A(_23752_),
    .X(_23757_));
 sky130_fd_sc_hd__o21ai_4 _30309_ (.A1(_22823_),
    .A2(_23756_),
    .B1(_23757_),
    .Y(_00184_));
 sky130_fd_sc_hd__buf_1 _30310_ (.A(_23745_),
    .X(_23758_));
 sky130_fd_sc_hd__o21ai_4 _30311_ (.A1(_22860_),
    .A2(_23758_),
    .B1(_23757_),
    .Y(_00185_));
 sky130_fd_sc_hd__o21ai_4 _30312_ (.A1(_22885_),
    .A2(_23758_),
    .B1(_23757_),
    .Y(_00187_));
 sky130_fd_sc_hd__a21bo_4 _30313_ (.A1(\decoded_imm_uj[31] ),
    .A2(_23727_),
    .B1_N(_23757_),
    .X(_00188_));
 sky130_vsdinv _30314_ (.A(\mem_rdata_q[24] ),
    .Y(_23759_));
 sky130_fd_sc_hd__nand3_4 _30315_ (.A(mem_rdata[24]),
    .B(_23724_),
    .C(_23725_),
    .Y(_23760_));
 sky130_fd_sc_hd__o21ai_4 _30316_ (.A1(_23759_),
    .A2(_23723_),
    .B1(_23760_),
    .Y(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__nand4_4 _30317_ (.A(_22929_),
    .B(_23708_),
    .C(_23730_),
    .D(\mem_rdata_latched[24] ),
    .Y(_23761_));
 sky130_fd_sc_hd__o21ai_4 _30318_ (.A1(_22114_),
    .A2(_23758_),
    .B1(_23761_),
    .Y(_00190_));
 sky130_vsdinv _30319_ (.A(\mem_rdata_q[20] ),
    .Y(_23762_));
 sky130_fd_sc_hd__nand3_4 _30320_ (.A(mem_rdata[20]),
    .B(_23735_),
    .C(_23737_),
    .Y(_23763_));
 sky130_fd_sc_hd__o21ai_4 _30321_ (.A1(_23762_),
    .A2(_23723_),
    .B1(_23763_),
    .Y(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__nand4_4 _30322_ (.A(_23739_),
    .B(_23728_),
    .C(_23730_),
    .D(\mem_rdata_latched[20] ),
    .Y(_23764_));
 sky130_fd_sc_hd__o21ai_4 _30323_ (.A1(_22358_),
    .A2(_23758_),
    .B1(_23764_),
    .Y(_00166_));
 sky130_fd_sc_hd__and2_4 _30324_ (.A(_23691_),
    .B(_21924_),
    .X(_00164_));
 sky130_fd_sc_hd__nand3_4 _30325_ (.A(mem_rdata[15]),
    .B(_18200_),
    .C(_18201_),
    .Y(_23765_));
 sky130_fd_sc_hd__a21bo_4 _30326_ (.A1(\mem_rdata_q[15] ),
    .A2(_18199_),
    .B1_N(_23765_),
    .X(\mem_rdata_latched[15] ));
 sky130_vsdinv _30327_ (.A(\mem_rdata_q[16] ),
    .Y(_23766_));
 sky130_fd_sc_hd__nand3_4 _30328_ (.A(mem_rdata[16]),
    .B(_23734_),
    .C(_23736_),
    .Y(_23767_));
 sky130_fd_sc_hd__o21ai_4 _30329_ (.A1(_23766_),
    .A2(_18871_),
    .B1(_23767_),
    .Y(\mem_rdata_latched[16] ));
 sky130_vsdinv _30330_ (.A(\mem_rdata_q[17] ),
    .Y(_23768_));
 sky130_fd_sc_hd__nand3_4 _30331_ (.A(mem_rdata[17]),
    .B(_23734_),
    .C(_23736_),
    .Y(_23769_));
 sky130_fd_sc_hd__o21ai_4 _30332_ (.A1(_23768_),
    .A2(_18871_),
    .B1(_23769_),
    .Y(\mem_rdata_latched[17] ));
 sky130_vsdinv _30333_ (.A(\mem_rdata_q[18] ),
    .Y(_23770_));
 sky130_fd_sc_hd__nand3_4 _30334_ (.A(mem_rdata[18]),
    .B(_23734_),
    .C(_23736_),
    .Y(_23771_));
 sky130_fd_sc_hd__o21ai_4 _30335_ (.A1(_23770_),
    .A2(_18831_),
    .B1(_23771_),
    .Y(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__nand4_4 _30336_ (.A(\mem_rdata_latched[26] ),
    .B(_23700_),
    .C(_23703_),
    .D(_18209_),
    .Y(_23772_));
 sky130_fd_sc_hd__buf_1 _30337_ (.A(_18232_),
    .X(_23773_));
 sky130_fd_sc_hd__and4_4 _30338_ (.A(_18401_),
    .B(_23773_),
    .C(_23711_),
    .D(\mem_rdata_latched[15] ),
    .X(_23774_));
 sky130_fd_sc_hd__and2_4 _30339_ (.A(_23772_),
    .B(_23774_),
    .X(_23775_));
 sky130_fd_sc_hd__a21o_4 _30340_ (.A1(\decoded_rs1[0] ),
    .A2(_23716_),
    .B1(_23775_),
    .X(_00201_));
 sky130_fd_sc_hd__and4_4 _30341_ (.A(_18401_),
    .B(_23773_),
    .C(_23711_),
    .D(\mem_rdata_latched[16] ),
    .X(_23776_));
 sky130_fd_sc_hd__and2_4 _30342_ (.A(_23772_),
    .B(_23776_),
    .X(_23777_));
 sky130_fd_sc_hd__a21o_4 _30343_ (.A1(\decoded_rs1[1] ),
    .A2(_23716_),
    .B1(_23777_),
    .X(_00202_));
 sky130_fd_sc_hd__and4_4 _30344_ (.A(_18401_),
    .B(_23773_),
    .C(_23711_),
    .D(\mem_rdata_latched[17] ),
    .X(_23778_));
 sky130_fd_sc_hd__and2_4 _30345_ (.A(_23772_),
    .B(_23778_),
    .X(_23779_));
 sky130_fd_sc_hd__a21o_4 _30346_ (.A1(\decoded_rs1[2] ),
    .A2(_23716_),
    .B1(_23779_),
    .X(_00203_));
 sky130_fd_sc_hd__buf_1 _30347_ (.A(_23715_),
    .X(_23780_));
 sky130_fd_sc_hd__buf_1 _30348_ (.A(_19048_),
    .X(_23781_));
 sky130_fd_sc_hd__and4_4 _30349_ (.A(_18360_),
    .B(_23773_),
    .C(_23781_),
    .D(\mem_rdata_latched[18] ),
    .X(_23782_));
 sky130_fd_sc_hd__and2_4 _30350_ (.A(_23772_),
    .B(_23782_),
    .X(_23783_));
 sky130_fd_sc_hd__a21o_4 _30351_ (.A1(\decoded_rs1[3] ),
    .A2(_23780_),
    .B1(_23783_),
    .X(_00204_));
 sky130_fd_sc_hd__buf_1 _30352_ (.A(is_alu_reg_reg),
    .X(_23784_));
 sky130_fd_sc_hd__buf_1 _30353_ (.A(_23784_),
    .X(_23785_));
 sky130_fd_sc_hd__nand2_4 _30354_ (.A(_18215_),
    .B(_18222_),
    .Y(_23786_));
 sky130_fd_sc_hd__nand4_4 _30355_ (.A(_18835_),
    .B(_23717_),
    .C(_23729_),
    .D(\mem_rdata_latched[4] ),
    .Y(_23787_));
 sky130_fd_sc_hd__and4_4 _30356_ (.A(\mem_rdata_latched[1] ),
    .B(\mem_rdata_latched[0] ),
    .C(_18197_),
    .D(_18205_),
    .X(_23788_));
 sky130_fd_sc_hd__buf_1 _30357_ (.A(_23788_),
    .X(_23789_));
 sky130_vsdinv _30358_ (.A(_23789_),
    .Y(_23790_));
 sky130_fd_sc_hd__nor3_4 _30359_ (.A(_23786_),
    .B(_23787_),
    .C(_23790_),
    .Y(_23791_));
 sky130_fd_sc_hd__a21o_4 _30360_ (.A1(_23785_),
    .A2(_23780_),
    .B1(_23791_),
    .X(_00363_));
 sky130_fd_sc_hd__buf_1 _30361_ (.A(is_alu_reg_imm),
    .X(_23792_));
 sky130_fd_sc_hd__buf_1 _30362_ (.A(_23792_),
    .X(_23793_));
 sky130_fd_sc_hd__nor4_4 _30363_ (.A(\mem_rdata_latched[5] ),
    .B(\mem_rdata_latched[6] ),
    .C(_23787_),
    .D(_23790_),
    .Y(_23794_));
 sky130_fd_sc_hd__a21o_4 _30364_ (.A1(_23793_),
    .A2(_23780_),
    .B1(_23794_),
    .X(_00362_));
 sky130_fd_sc_hd__buf_1 _30365_ (.A(_19051_),
    .X(_23795_));
 sky130_fd_sc_hd__nor2_4 _30366_ (.A(_23715_),
    .B(_23790_),
    .Y(_23796_));
 sky130_fd_sc_hd__nand4_4 _30367_ (.A(\mem_rdata_latched[5] ),
    .B(_23796_),
    .C(_18217_),
    .D(_18222_),
    .Y(_23797_));
 sky130_fd_sc_hd__o21ai_4 _30368_ (.A1(_18808_),
    .A2(_23795_),
    .B1(_23797_),
    .Y(_00369_));
 sky130_fd_sc_hd__nor2_4 _30369_ (.A(decoder_pseudo_trigger),
    .B(_19134_),
    .Y(_23798_));
 sky130_vsdinv _30370_ (.A(_23798_),
    .Y(_23799_));
 sky130_fd_sc_hd__buf_1 _30371_ (.A(_23799_),
    .X(_23800_));
 sky130_fd_sc_hd__buf_1 _30372_ (.A(_23800_),
    .X(_23801_));
 sky130_fd_sc_hd__buf_1 _30373_ (.A(_23801_),
    .X(_23802_));
 sky130_fd_sc_hd__buf_1 _30374_ (.A(_23799_),
    .X(_23803_));
 sky130_fd_sc_hd__buf_1 _30375_ (.A(_23803_),
    .X(_23804_));
 sky130_vsdinv _30376_ (.A(is_alu_reg_imm),
    .Y(_23805_));
 sky130_fd_sc_hd__buf_1 _30377_ (.A(\mem_rdata_q[13] ),
    .X(_23806_));
 sky130_fd_sc_hd__buf_1 _30378_ (.A(_23806_),
    .X(_23807_));
 sky130_fd_sc_hd__buf_1 _30379_ (.A(_18870_),
    .X(_23808_));
 sky130_fd_sc_hd__nor2_4 _30380_ (.A(_23807_),
    .B(_23808_),
    .Y(_23809_));
 sky130_vsdinv _30381_ (.A(instr_jalr),
    .Y(_23810_));
 sky130_fd_sc_hd__o21a_4 _30382_ (.A1(_23805_),
    .A2(_23809_),
    .B1(_23810_),
    .X(_23811_));
 sky130_fd_sc_hd__nor2_4 _30383_ (.A(_23804_),
    .B(_23811_),
    .Y(_23812_));
 sky130_fd_sc_hd__a21o_4 _30384_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(_23802_),
    .B1(_23812_),
    .X(_00366_));
 sky130_fd_sc_hd__buf_1 _30385_ (.A(_23798_),
    .X(_23813_));
 sky130_fd_sc_hd__buf_1 _30386_ (.A(_23813_),
    .X(_23814_));
 sky130_fd_sc_hd__buf_1 _30387_ (.A(_23814_),
    .X(_23815_));
 sky130_fd_sc_hd__buf_1 _30388_ (.A(_23815_),
    .X(_23816_));
 sky130_fd_sc_hd__buf_1 _30389_ (.A(\mem_rdata_q[27] ),
    .X(_23817_));
 sky130_fd_sc_hd__nor2_4 _30390_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[31] ),
    .Y(_23818_));
 sky130_fd_sc_hd__buf_1 _30391_ (.A(\mem_rdata_q[29] ),
    .X(_23819_));
 sky130_vsdinv _30392_ (.A(_23819_),
    .Y(_23820_));
 sky130_fd_sc_hd__nand3_4 _30393_ (.A(_23818_),
    .B(_23820_),
    .C(\mem_rdata_q[30] ),
    .Y(_23821_));
 sky130_fd_sc_hd__nor4_4 _30394_ (.A(_18198_),
    .B(_23817_),
    .C(\mem_rdata_q[25] ),
    .D(_23821_),
    .Y(_23822_));
 sky130_fd_sc_hd__buf_1 _30395_ (.A(\mem_rdata_q[14] ),
    .X(_23823_));
 sky130_fd_sc_hd__buf_1 _30396_ (.A(_23823_),
    .X(_23824_));
 sky130_fd_sc_hd__nand2_4 _30397_ (.A(_23822_),
    .B(_23824_),
    .Y(_23825_));
 sky130_fd_sc_hd__nor2_4 _30398_ (.A(\mem_rdata_q[26] ),
    .B(\mem_rdata_q[27] ),
    .Y(_23826_));
 sky130_fd_sc_hd__nor2_4 _30399_ (.A(_23819_),
    .B(\mem_rdata_q[30] ),
    .Y(_23827_));
 sky130_fd_sc_hd__buf_1 _30400_ (.A(_18827_),
    .X(_23828_));
 sky130_fd_sc_hd__and4_4 _30401_ (.A(_23826_),
    .B(_23818_),
    .C(_23827_),
    .D(_23828_),
    .X(_23829_));
 sky130_vsdinv _30402_ (.A(_23829_),
    .Y(_23830_));
 sky130_fd_sc_hd__buf_1 _30403_ (.A(_23806_),
    .X(_23831_));
 sky130_fd_sc_hd__nand2_4 _30404_ (.A(_23814_),
    .B(_23792_),
    .Y(_23832_));
 sky130_fd_sc_hd__a2111o_4 _30405_ (.A1(_23825_),
    .A2(_23830_),
    .B1(_23808_),
    .C1(_23831_),
    .D1(_23832_),
    .X(_23833_));
 sky130_fd_sc_hd__o21ai_4 _30406_ (.A1(_21183_),
    .A2(_23816_),
    .B1(_23833_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand3_4 _30407_ (.A(_23706_),
    .B(_23701_),
    .C(_23789_),
    .Y(_23834_));
 sky130_fd_sc_hd__o21ai_4 _30408_ (.A1(_18287_),
    .A2(_23795_),
    .B1(_23834_),
    .Y(_00367_));
 sky130_fd_sc_hd__nor3_4 _30409_ (.A(_19142_),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(is_alu_reg_imm),
    .Y(_23835_));
 sky130_fd_sc_hd__buf_1 _30410_ (.A(_23835_),
    .X(_23836_));
 sky130_fd_sc_hd__buf_1 _30411_ (.A(is_sb_sh_sw),
    .X(_23837_));
 sky130_fd_sc_hd__a22oi_4 _30412_ (.A1(_22176_),
    .A2(_21924_),
    .B1(_23837_),
    .B2(\mem_rdata_q[7] ),
    .Y(_23838_));
 sky130_fd_sc_hd__o21a_4 _30413_ (.A1(_23762_),
    .A2(_23836_),
    .B1(_23838_),
    .X(_23839_));
 sky130_fd_sc_hd__nor2_4 _30414_ (.A(_23804_),
    .B(_23839_),
    .Y(_23840_));
 sky130_fd_sc_hd__a21o_4 _30415_ (.A1(_21345_),
    .A2(_23802_),
    .B1(_23840_),
    .X(_00132_));
 sky130_vsdinv _30416_ (.A(\mem_rdata_q[8] ),
    .Y(_23841_));
 sky130_fd_sc_hd__nor2_4 _30417_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(_23837_),
    .Y(_23842_));
 sky130_fd_sc_hd__a2bb2oi_4 _30418_ (.A1_N(_23841_),
    .A2_N(_23842_),
    .B1(_22544_),
    .B2(\decoded_imm_uj[1] ),
    .Y(_23843_));
 sky130_fd_sc_hd__o21ai_4 _30419_ (.A1(_23722_),
    .A2(_23836_),
    .B1(_23843_),
    .Y(_23844_));
 sky130_fd_sc_hd__buf_1 _30420_ (.A(_23798_),
    .X(_23845_));
 sky130_fd_sc_hd__buf_1 _30421_ (.A(_23845_),
    .X(_23846_));
 sky130_fd_sc_hd__buf_1 _30422_ (.A(_23846_),
    .X(_23847_));
 sky130_fd_sc_hd__nand2_4 _30423_ (.A(_23844_),
    .B(_23847_),
    .Y(_23848_));
 sky130_fd_sc_hd__o21ai_4 _30424_ (.A1(_21373_),
    .A2(_23816_),
    .B1(_23848_),
    .Y(_00143_));
 sky130_vsdinv _30425_ (.A(_23835_),
    .Y(_23849_));
 sky130_vsdinv _30426_ (.A(\mem_rdata_q[9] ),
    .Y(_23850_));
 sky130_fd_sc_hd__a2bb2o_4 _30427_ (.A1_N(_23850_),
    .A2_N(_23842_),
    .B1(_18775_),
    .B2(\decoded_imm_uj[2] ),
    .X(_23851_));
 sky130_fd_sc_hd__a21o_4 _30428_ (.A1(_23732_),
    .A2(_23849_),
    .B1(_23851_),
    .X(_23852_));
 sky130_fd_sc_hd__buf_1 _30429_ (.A(_23845_),
    .X(_23853_));
 sky130_fd_sc_hd__and2_4 _30430_ (.A(_23852_),
    .B(_23853_),
    .X(_23854_));
 sky130_fd_sc_hd__a21o_4 _30431_ (.A1(_21147_),
    .A2(_23802_),
    .B1(_23854_),
    .X(_00154_));
 sky130_vsdinv _30432_ (.A(\mem_rdata_q[10] ),
    .Y(_23855_));
 sky130_fd_sc_hd__a2bb2o_4 _30433_ (.A1_N(_23855_),
    .A2_N(_23842_),
    .B1(_22176_),
    .B2(\decoded_imm_uj[3] ),
    .X(_23856_));
 sky130_fd_sc_hd__a21o_4 _30434_ (.A1(_23742_),
    .A2(_23849_),
    .B1(_23856_),
    .X(_23857_));
 sky130_fd_sc_hd__buf_1 _30435_ (.A(_23846_),
    .X(_23858_));
 sky130_fd_sc_hd__nand2_4 _30436_ (.A(_23857_),
    .B(_23858_),
    .Y(_23859_));
 sky130_fd_sc_hd__o21ai_4 _30437_ (.A1(_21160_),
    .A2(_23816_),
    .B1(_23859_),
    .Y(_00157_));
 sky130_vsdinv _30438_ (.A(\mem_rdata_q[11] ),
    .Y(_23860_));
 sky130_fd_sc_hd__o22a_4 _30439_ (.A1(_21923_),
    .A2(_22114_),
    .B1(_23860_),
    .B2(_23842_),
    .X(_23861_));
 sky130_fd_sc_hd__o21ai_4 _30440_ (.A1(_23759_),
    .A2(_23836_),
    .B1(_23861_),
    .Y(_23862_));
 sky130_fd_sc_hd__nand2_4 _30441_ (.A(_23862_),
    .B(_23858_),
    .Y(_23863_));
 sky130_fd_sc_hd__o21ai_4 _30442_ (.A1(_21173_),
    .A2(_23816_),
    .B1(_23863_),
    .Y(_00158_));
 sky130_fd_sc_hd__buf_1 _30443_ (.A(_21922_),
    .X(_23864_));
 sky130_fd_sc_hd__buf_1 _30444_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_23865_));
 sky130_fd_sc_hd__nand4_4 _30445_ (.A(_23810_),
    .B(_18287_),
    .C(_18807_),
    .D(_23805_),
    .Y(_23866_));
 sky130_fd_sc_hd__nor2_4 _30446_ (.A(_23865_),
    .B(_23866_),
    .Y(_23867_));
 sky130_fd_sc_hd__buf_1 _30447_ (.A(_23867_),
    .X(_23868_));
 sky130_fd_sc_hd__o22a_4 _30448_ (.A1(_23864_),
    .A2(_22138_),
    .B1(_23828_),
    .B2(_23868_),
    .X(_23869_));
 sky130_fd_sc_hd__nor2_4 _30449_ (.A(_23804_),
    .B(_23869_),
    .Y(_23870_));
 sky130_fd_sc_hd__a21o_4 _30450_ (.A1(_21186_),
    .A2(_23802_),
    .B1(_23870_),
    .X(_00159_));
 sky130_fd_sc_hd__buf_1 _30451_ (.A(_23801_),
    .X(_23871_));
 sky130_fd_sc_hd__buf_1 _30452_ (.A(_23803_),
    .X(_23872_));
 sky130_vsdinv _30453_ (.A(_18198_),
    .Y(_23873_));
 sky130_fd_sc_hd__o22a_4 _30454_ (.A1(_23864_),
    .A2(_22198_),
    .B1(_23873_),
    .B2(_23868_),
    .X(_23874_));
 sky130_fd_sc_hd__nor2_4 _30455_ (.A(_23872_),
    .B(_23874_),
    .Y(_23875_));
 sky130_fd_sc_hd__a21o_4 _30456_ (.A1(_21193_),
    .A2(_23871_),
    .B1(_23875_),
    .X(_00160_));
 sky130_vsdinv _30457_ (.A(_23817_),
    .Y(_23876_));
 sky130_fd_sc_hd__a2bb2oi_4 _30458_ (.A1_N(_23876_),
    .A2_N(_23868_),
    .B1(_21950_),
    .B2(\decoded_imm_uj[7] ),
    .Y(_23877_));
 sky130_fd_sc_hd__nor2_4 _30459_ (.A(_23872_),
    .B(_23877_),
    .Y(_23878_));
 sky130_fd_sc_hd__a21o_4 _30460_ (.A1(_21201_),
    .A2(_23871_),
    .B1(_23878_),
    .X(_00161_));
 sky130_fd_sc_hd__o22a_4 _30461_ (.A1(_23864_),
    .A2(_22230_),
    .B1(_18830_),
    .B2(_23868_),
    .X(_23879_));
 sky130_fd_sc_hd__nor2_4 _30462_ (.A(_23872_),
    .B(_23879_),
    .Y(_23880_));
 sky130_fd_sc_hd__a21o_4 _30463_ (.A1(_21207_),
    .A2(_23871_),
    .B1(_23880_),
    .X(_00162_));
 sky130_fd_sc_hd__o22a_4 _30464_ (.A1(_23864_),
    .A2(_22298_),
    .B1(_23820_),
    .B2(_23867_),
    .X(_23881_));
 sky130_fd_sc_hd__nor2_4 _30465_ (.A(_23872_),
    .B(_23881_),
    .Y(_23882_));
 sky130_fd_sc_hd__a21o_4 _30466_ (.A1(_21531_),
    .A2(_23871_),
    .B1(_23882_),
    .X(_00163_));
 sky130_fd_sc_hd__buf_1 _30467_ (.A(_23800_),
    .X(_23883_));
 sky130_fd_sc_hd__buf_1 _30468_ (.A(_23883_),
    .X(_23884_));
 sky130_fd_sc_hd__buf_1 _30469_ (.A(_23800_),
    .X(_23885_));
 sky130_fd_sc_hd__nand3_4 _30470_ (.A(_23836_),
    .B(_18864_),
    .C(_18808_),
    .Y(_23886_));
 sky130_fd_sc_hd__buf_1 _30471_ (.A(\mem_rdata_q[30] ),
    .X(_23887_));
 sky130_fd_sc_hd__a22oi_4 _30472_ (.A1(_22544_),
    .A2(\decoded_imm_uj[10] ),
    .B1(_23886_),
    .B2(_23887_),
    .Y(_23888_));
 sky130_fd_sc_hd__nor2_4 _30473_ (.A(_23885_),
    .B(_23888_),
    .Y(_23889_));
 sky130_fd_sc_hd__a21o_4 _30474_ (.A1(_21222_),
    .A2(_23884_),
    .B1(_23889_),
    .X(_00133_));
 sky130_fd_sc_hd__buf_1 _30475_ (.A(\mem_rdata_q[31] ),
    .X(_23890_));
 sky130_fd_sc_hd__a22oi_4 _30476_ (.A1(_22176_),
    .A2(\decoded_imm_uj[11] ),
    .B1(_23865_),
    .B2(\mem_rdata_q[7] ),
    .Y(_23891_));
 sky130_fd_sc_hd__a21boi_4 _30477_ (.A1(_23866_),
    .A2(_23890_),
    .B1_N(_23891_),
    .Y(_23892_));
 sky130_fd_sc_hd__nor2_4 _30478_ (.A(_23885_),
    .B(_23892_),
    .Y(_23893_));
 sky130_fd_sc_hd__a21o_4 _30479_ (.A1(_21232_),
    .A2(_23884_),
    .B1(_23893_),
    .X(_00134_));
 sky130_fd_sc_hd__o21ai_4 _30480_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(_23866_),
    .B1(\mem_rdata_q[31] ),
    .Y(_23894_));
 sky130_fd_sc_hd__buf_1 _30481_ (.A(_23894_),
    .X(_23895_));
 sky130_fd_sc_hd__buf_1 _30482_ (.A(_23895_),
    .X(_23896_));
 sky130_fd_sc_hd__nand2_4 _30483_ (.A(_22507_),
    .B(\decoded_imm_uj[12] ),
    .Y(_23897_));
 sky130_fd_sc_hd__buf_1 _30484_ (.A(instr_auipc),
    .X(_23898_));
 sky130_fd_sc_hd__buf_1 _30485_ (.A(instr_lui),
    .X(_23899_));
 sky130_fd_sc_hd__buf_1 _30486_ (.A(\mem_rdata_q[12] ),
    .X(_23900_));
 sky130_fd_sc_hd__o21ai_4 _30487_ (.A1(_23898_),
    .A2(_23899_),
    .B1(_23900_),
    .Y(_23901_));
 sky130_fd_sc_hd__nand3_4 _30488_ (.A(_23896_),
    .B(_23897_),
    .C(_23901_),
    .Y(_23902_));
 sky130_fd_sc_hd__and2_4 _30489_ (.A(_23902_),
    .B(_23853_),
    .X(_23903_));
 sky130_fd_sc_hd__a21o_4 _30490_ (.A1(_21239_),
    .A2(_23884_),
    .B1(_23903_),
    .X(_00135_));
 sky130_fd_sc_hd__nand2_4 _30491_ (.A(_22507_),
    .B(\decoded_imm_uj[13] ),
    .Y(_23904_));
 sky130_fd_sc_hd__buf_1 _30492_ (.A(instr_auipc),
    .X(_23905_));
 sky130_fd_sc_hd__o21ai_4 _30493_ (.A1(_23905_),
    .A2(_23899_),
    .B1(_23807_),
    .Y(_23906_));
 sky130_fd_sc_hd__nand3_4 _30494_ (.A(_23896_),
    .B(_23904_),
    .C(_23906_),
    .Y(_23907_));
 sky130_fd_sc_hd__buf_1 _30495_ (.A(_23813_),
    .X(_23908_));
 sky130_fd_sc_hd__buf_1 _30496_ (.A(_23908_),
    .X(_23909_));
 sky130_fd_sc_hd__and2_4 _30497_ (.A(_23907_),
    .B(_23909_),
    .X(_23910_));
 sky130_fd_sc_hd__a21o_4 _30498_ (.A1(_21603_),
    .A2(_23884_),
    .B1(_23910_),
    .X(_00136_));
 sky130_fd_sc_hd__buf_1 _30499_ (.A(_23883_),
    .X(_23911_));
 sky130_fd_sc_hd__buf_1 _30500_ (.A(_23905_),
    .X(_23912_));
 sky130_fd_sc_hd__buf_1 _30501_ (.A(instr_lui),
    .X(_23913_));
 sky130_fd_sc_hd__buf_1 _30502_ (.A(_23913_),
    .X(_23914_));
 sky130_fd_sc_hd__o21ai_4 _30503_ (.A1(_23912_),
    .A2(_23914_),
    .B1(_23823_),
    .Y(_23915_));
 sky130_fd_sc_hd__nand2_4 _30504_ (.A(_22619_),
    .B(\decoded_imm_uj[14] ),
    .Y(_23916_));
 sky130_fd_sc_hd__nand3_4 _30505_ (.A(_23896_),
    .B(_23915_),
    .C(_23916_),
    .Y(_23917_));
 sky130_fd_sc_hd__and2_4 _30506_ (.A(_23917_),
    .B(_23909_),
    .X(_23918_));
 sky130_fd_sc_hd__a21o_4 _30507_ (.A1(_21253_),
    .A2(_23911_),
    .B1(_23918_),
    .X(_00137_));
 sky130_fd_sc_hd__o21ai_4 _30508_ (.A1(_23912_),
    .A2(_23914_),
    .B1(\mem_rdata_q[15] ),
    .Y(_23919_));
 sky130_fd_sc_hd__nand2_4 _30509_ (.A(_22619_),
    .B(_22446_),
    .Y(_23920_));
 sky130_fd_sc_hd__nand3_4 _30510_ (.A(_23896_),
    .B(_23919_),
    .C(_23920_),
    .Y(_23921_));
 sky130_fd_sc_hd__and2_4 _30511_ (.A(_23921_),
    .B(_23909_),
    .X(_23922_));
 sky130_fd_sc_hd__a21o_4 _30512_ (.A1(_21258_),
    .A2(_23911_),
    .B1(_23922_),
    .X(_00138_));
 sky130_fd_sc_hd__buf_1 _30513_ (.A(_23894_),
    .X(_23923_));
 sky130_fd_sc_hd__buf_1 _30514_ (.A(_23905_),
    .X(_23924_));
 sky130_fd_sc_hd__o21ai_4 _30515_ (.A1(_23924_),
    .A2(_23914_),
    .B1(\mem_rdata_q[16] ),
    .Y(_23925_));
 sky130_fd_sc_hd__nand2_4 _30516_ (.A(_22619_),
    .B(\decoded_imm_uj[16] ),
    .Y(_23926_));
 sky130_fd_sc_hd__nand3_4 _30517_ (.A(_23923_),
    .B(_23925_),
    .C(_23926_),
    .Y(_23927_));
 sky130_fd_sc_hd__and2_4 _30518_ (.A(_23927_),
    .B(_23909_),
    .X(_23928_));
 sky130_fd_sc_hd__a21o_4 _30519_ (.A1(_21264_),
    .A2(_23911_),
    .B1(_23928_),
    .X(_00139_));
 sky130_fd_sc_hd__buf_1 _30520_ (.A(_23913_),
    .X(_23929_));
 sky130_fd_sc_hd__o21ai_4 _30521_ (.A1(_23924_),
    .A2(_23929_),
    .B1(\mem_rdata_q[17] ),
    .Y(_23930_));
 sky130_fd_sc_hd__buf_1 _30522_ (.A(_22618_),
    .X(_23931_));
 sky130_fd_sc_hd__nand2_4 _30523_ (.A(_23931_),
    .B(\decoded_imm_uj[17] ),
    .Y(_23932_));
 sky130_fd_sc_hd__nand3_4 _30524_ (.A(_23923_),
    .B(_23930_),
    .C(_23932_),
    .Y(_23933_));
 sky130_fd_sc_hd__buf_1 _30525_ (.A(_23908_),
    .X(_23934_));
 sky130_fd_sc_hd__and2_4 _30526_ (.A(_23933_),
    .B(_23934_),
    .X(_23935_));
 sky130_fd_sc_hd__a21o_4 _30527_ (.A1(_21270_),
    .A2(_23911_),
    .B1(_23935_),
    .X(_00140_));
 sky130_fd_sc_hd__buf_1 _30528_ (.A(_23883_),
    .X(_23936_));
 sky130_fd_sc_hd__o21ai_4 _30529_ (.A1(_23924_),
    .A2(_23929_),
    .B1(\mem_rdata_q[18] ),
    .Y(_23937_));
 sky130_fd_sc_hd__nand2_4 _30530_ (.A(_23931_),
    .B(\decoded_imm_uj[18] ),
    .Y(_23938_));
 sky130_fd_sc_hd__nand3_4 _30531_ (.A(_23923_),
    .B(_23937_),
    .C(_23938_),
    .Y(_23939_));
 sky130_fd_sc_hd__and2_4 _30532_ (.A(_23939_),
    .B(_23934_),
    .X(_23940_));
 sky130_fd_sc_hd__a21o_4 _30533_ (.A1(_21274_),
    .A2(_23936_),
    .B1(_23940_),
    .X(_00141_));
 sky130_fd_sc_hd__o21ai_4 _30534_ (.A1(_23924_),
    .A2(_23929_),
    .B1(\mem_rdata_q[19] ),
    .Y(_23941_));
 sky130_fd_sc_hd__nand2_4 _30535_ (.A(_23931_),
    .B(\decoded_imm_uj[19] ),
    .Y(_23942_));
 sky130_fd_sc_hd__nand3_4 _30536_ (.A(_23923_),
    .B(_23941_),
    .C(_23942_),
    .Y(_23943_));
 sky130_fd_sc_hd__and2_4 _30537_ (.A(_23943_),
    .B(_23934_),
    .X(_23944_));
 sky130_fd_sc_hd__a21o_4 _30538_ (.A1(_21281_),
    .A2(_23936_),
    .B1(_23944_),
    .X(_00142_));
 sky130_fd_sc_hd__buf_1 _30539_ (.A(_23894_),
    .X(_23945_));
 sky130_fd_sc_hd__buf_1 _30540_ (.A(_23905_),
    .X(_23946_));
 sky130_fd_sc_hd__o21ai_4 _30541_ (.A1(_23946_),
    .A2(_23929_),
    .B1(\mem_rdata_q[20] ),
    .Y(_23947_));
 sky130_fd_sc_hd__nand2_4 _30542_ (.A(_23931_),
    .B(\decoded_imm_uj[20] ),
    .Y(_23948_));
 sky130_fd_sc_hd__nand3_4 _30543_ (.A(_23945_),
    .B(_23947_),
    .C(_23948_),
    .Y(_23949_));
 sky130_fd_sc_hd__and2_4 _30544_ (.A(_23949_),
    .B(_23934_),
    .X(_23950_));
 sky130_fd_sc_hd__a21o_4 _30545_ (.A1(_21286_),
    .A2(_23936_),
    .B1(_23950_),
    .X(_00144_));
 sky130_fd_sc_hd__buf_1 _30546_ (.A(_23913_),
    .X(_23951_));
 sky130_fd_sc_hd__o21ai_4 _30547_ (.A1(_23946_),
    .A2(_23951_),
    .B1(\mem_rdata_q[21] ),
    .Y(_23952_));
 sky130_fd_sc_hd__buf_1 _30548_ (.A(_22618_),
    .X(_23953_));
 sky130_fd_sc_hd__nand2_4 _30549_ (.A(_23953_),
    .B(\decoded_imm_uj[21] ),
    .Y(_23954_));
 sky130_fd_sc_hd__nand3_4 _30550_ (.A(_23945_),
    .B(_23952_),
    .C(_23954_),
    .Y(_23955_));
 sky130_fd_sc_hd__buf_1 _30551_ (.A(_23908_),
    .X(_23956_));
 sky130_fd_sc_hd__and2_4 _30552_ (.A(_23955_),
    .B(_23956_),
    .X(_23957_));
 sky130_fd_sc_hd__a21o_4 _30553_ (.A1(_21292_),
    .A2(_23936_),
    .B1(_23957_),
    .X(_00145_));
 sky130_fd_sc_hd__buf_1 _30554_ (.A(_23883_),
    .X(_23958_));
 sky130_fd_sc_hd__o21ai_4 _30555_ (.A1(_23946_),
    .A2(_23951_),
    .B1(_23732_),
    .Y(_23959_));
 sky130_fd_sc_hd__nand2_4 _30556_ (.A(_23953_),
    .B(\decoded_imm_uj[22] ),
    .Y(_23960_));
 sky130_fd_sc_hd__nand3_4 _30557_ (.A(_23945_),
    .B(_23959_),
    .C(_23960_),
    .Y(_23961_));
 sky130_fd_sc_hd__and2_4 _30558_ (.A(_23961_),
    .B(_23956_),
    .X(_23962_));
 sky130_fd_sc_hd__a21o_4 _30559_ (.A1(_21296_),
    .A2(_23958_),
    .B1(_23962_),
    .X(_00146_));
 sky130_fd_sc_hd__o21ai_4 _30560_ (.A1(_23946_),
    .A2(_23951_),
    .B1(_23742_),
    .Y(_23963_));
 sky130_fd_sc_hd__nand2_4 _30561_ (.A(_23953_),
    .B(\decoded_imm_uj[23] ),
    .Y(_23964_));
 sky130_fd_sc_hd__nand3_4 _30562_ (.A(_23945_),
    .B(_23963_),
    .C(_23964_),
    .Y(_23965_));
 sky130_fd_sc_hd__and2_4 _30563_ (.A(_23965_),
    .B(_23956_),
    .X(_23966_));
 sky130_fd_sc_hd__a21o_4 _30564_ (.A1(\decoded_imm[23] ),
    .A2(_23958_),
    .B1(_23966_),
    .X(_00147_));
 sky130_fd_sc_hd__buf_1 _30565_ (.A(_23894_),
    .X(_23967_));
 sky130_fd_sc_hd__buf_1 _30566_ (.A(instr_auipc),
    .X(_23968_));
 sky130_fd_sc_hd__o21ai_4 _30567_ (.A1(_23968_),
    .A2(_23951_),
    .B1(\mem_rdata_q[24] ),
    .Y(_23969_));
 sky130_fd_sc_hd__nand2_4 _30568_ (.A(_23953_),
    .B(\decoded_imm_uj[24] ),
    .Y(_23970_));
 sky130_fd_sc_hd__nand3_4 _30569_ (.A(_23967_),
    .B(_23969_),
    .C(_23970_),
    .Y(_23971_));
 sky130_fd_sc_hd__and2_4 _30570_ (.A(_23971_),
    .B(_23956_),
    .X(_23972_));
 sky130_fd_sc_hd__a21o_4 _30571_ (.A1(_21305_),
    .A2(_23958_),
    .B1(_23972_),
    .X(_00148_));
 sky130_fd_sc_hd__buf_1 _30572_ (.A(_23913_),
    .X(_23973_));
 sky130_fd_sc_hd__buf_1 _30573_ (.A(\mem_rdata_q[25] ),
    .X(_23974_));
 sky130_fd_sc_hd__o21ai_4 _30574_ (.A1(_23968_),
    .A2(_23973_),
    .B1(_23974_),
    .Y(_23975_));
 sky130_fd_sc_hd__buf_1 _30575_ (.A(_22618_),
    .X(_23976_));
 sky130_fd_sc_hd__nand2_4 _30576_ (.A(_23976_),
    .B(\decoded_imm_uj[25] ),
    .Y(_23977_));
 sky130_fd_sc_hd__nand3_4 _30577_ (.A(_23967_),
    .B(_23975_),
    .C(_23977_),
    .Y(_23978_));
 sky130_fd_sc_hd__buf_1 _30578_ (.A(_23908_),
    .X(_23979_));
 sky130_fd_sc_hd__and2_4 _30579_ (.A(_23978_),
    .B(_23979_),
    .X(_23980_));
 sky130_fd_sc_hd__a21o_4 _30580_ (.A1(_21311_),
    .A2(_23958_),
    .B1(_23980_),
    .X(_00149_));
 sky130_fd_sc_hd__buf_1 _30581_ (.A(_23803_),
    .X(_23981_));
 sky130_fd_sc_hd__buf_1 _30582_ (.A(_18198_),
    .X(_23982_));
 sky130_fd_sc_hd__o21ai_4 _30583_ (.A1(_23968_),
    .A2(_23973_),
    .B1(_23982_),
    .Y(_23983_));
 sky130_fd_sc_hd__nand2_4 _30584_ (.A(_23976_),
    .B(\decoded_imm_uj[26] ),
    .Y(_23984_));
 sky130_fd_sc_hd__nand3_4 _30585_ (.A(_23967_),
    .B(_23983_),
    .C(_23984_),
    .Y(_23985_));
 sky130_fd_sc_hd__and2_4 _30586_ (.A(_23985_),
    .B(_23979_),
    .X(_23986_));
 sky130_fd_sc_hd__a21o_4 _30587_ (.A1(_21318_),
    .A2(_23981_),
    .B1(_23986_),
    .X(_00150_));
 sky130_fd_sc_hd__o21ai_4 _30588_ (.A1(_23968_),
    .A2(_23973_),
    .B1(_23817_),
    .Y(_23987_));
 sky130_fd_sc_hd__nand2_4 _30589_ (.A(_23976_),
    .B(\decoded_imm_uj[27] ),
    .Y(_23988_));
 sky130_fd_sc_hd__nand3_4 _30590_ (.A(_23967_),
    .B(_23987_),
    .C(_23988_),
    .Y(_23989_));
 sky130_fd_sc_hd__and2_4 _30591_ (.A(_23989_),
    .B(_23979_),
    .X(_23990_));
 sky130_fd_sc_hd__a21o_4 _30592_ (.A1(_21321_),
    .A2(_23981_),
    .B1(_23990_),
    .X(_00151_));
 sky130_fd_sc_hd__o21ai_4 _30593_ (.A1(_23898_),
    .A2(_23973_),
    .B1(\mem_rdata_q[28] ),
    .Y(_23991_));
 sky130_fd_sc_hd__nand2_4 _30594_ (.A(_23976_),
    .B(\decoded_imm_uj[28] ),
    .Y(_23992_));
 sky130_fd_sc_hd__nand3_4 _30595_ (.A(_23895_),
    .B(_23991_),
    .C(_23992_),
    .Y(_23993_));
 sky130_fd_sc_hd__and2_4 _30596_ (.A(_23993_),
    .B(_23979_),
    .X(_23994_));
 sky130_fd_sc_hd__a21o_4 _30597_ (.A1(_21326_),
    .A2(_23981_),
    .B1(_23994_),
    .X(_00152_));
 sky130_fd_sc_hd__o21ai_4 _30598_ (.A1(_23898_),
    .A2(_23899_),
    .B1(_23819_),
    .Y(_23995_));
 sky130_fd_sc_hd__nand2_4 _30599_ (.A(_21949_),
    .B(\decoded_imm_uj[29] ),
    .Y(_23996_));
 sky130_fd_sc_hd__nand3_4 _30600_ (.A(_23895_),
    .B(_23995_),
    .C(_23996_),
    .Y(_23997_));
 sky130_fd_sc_hd__buf_1 _30601_ (.A(_23814_),
    .X(_23998_));
 sky130_fd_sc_hd__and2_4 _30602_ (.A(_23997_),
    .B(_23998_),
    .X(_23999_));
 sky130_fd_sc_hd__a21o_4 _30603_ (.A1(_21331_),
    .A2(_23981_),
    .B1(_23999_),
    .X(_00153_));
 sky130_fd_sc_hd__buf_1 _30604_ (.A(_23803_),
    .X(_24000_));
 sky130_fd_sc_hd__o21ai_4 _30605_ (.A1(_23898_),
    .A2(_23899_),
    .B1(_23887_),
    .Y(_24001_));
 sky130_fd_sc_hd__nand2_4 _30606_ (.A(_21949_),
    .B(\decoded_imm_uj[30] ),
    .Y(_24002_));
 sky130_fd_sc_hd__nand3_4 _30607_ (.A(_23895_),
    .B(_24001_),
    .C(_24002_),
    .Y(_24003_));
 sky130_fd_sc_hd__and2_4 _30608_ (.A(_24003_),
    .B(_23998_),
    .X(_24004_));
 sky130_fd_sc_hd__a21o_4 _30609_ (.A1(_21336_),
    .A2(_24000_),
    .B1(_24004_),
    .X(_00155_));
 sky130_fd_sc_hd__buf_1 _30610_ (.A(_23813_),
    .X(_24005_));
 sky130_fd_sc_hd__buf_1 _30611_ (.A(_24005_),
    .X(_24006_));
 sky130_fd_sc_hd__buf_1 _30612_ (.A(_24006_),
    .X(_24007_));
 sky130_fd_sc_hd__buf_1 _30613_ (.A(_23865_),
    .X(_24008_));
 sky130_fd_sc_hd__o41ai_4 _30614_ (.A1(_23912_),
    .A2(_23914_),
    .A3(_24008_),
    .A4(_23866_),
    .B1(_23890_),
    .Y(_24009_));
 sky130_fd_sc_hd__nand2_4 _30615_ (.A(_21950_),
    .B(\decoded_imm_uj[31] ),
    .Y(_24010_));
 sky130_fd_sc_hd__a21o_4 _30616_ (.A1(_24009_),
    .A2(_24010_),
    .B1(_23885_),
    .X(_24011_));
 sky130_fd_sc_hd__o21ai_4 _30617_ (.A1(_21341_),
    .A2(_24007_),
    .B1(_24011_),
    .Y(_00156_));
 sky130_fd_sc_hd__o21ai_4 _30618_ (.A1(_19167_),
    .A2(_23795_),
    .B1(_23764_),
    .Y(_00206_));
 sky130_fd_sc_hd__o21ai_4 _30619_ (.A1(_19178_),
    .A2(_23795_),
    .B1(_23731_),
    .Y(_00207_));
 sky130_fd_sc_hd__buf_1 _30620_ (.A(_19051_),
    .X(_24012_));
 sky130_fd_sc_hd__o21ai_4 _30621_ (.A1(_19173_),
    .A2(_24012_),
    .B1(_23741_),
    .Y(_00208_));
 sky130_fd_sc_hd__o21ai_4 _30622_ (.A1(_19184_),
    .A2(_24012_),
    .B1(_23744_),
    .Y(_00209_));
 sky130_fd_sc_hd__a21bo_4 _30623_ (.A1(\decoded_rs2[4] ),
    .A2(_23727_),
    .B1_N(_23761_),
    .X(_00210_));
 sky130_fd_sc_hd__buf_1 _30624_ (.A(_23719_),
    .X(_24013_));
 sky130_fd_sc_hd__nand4_4 _30625_ (.A(_24013_),
    .B(_23748_),
    .C(_23750_),
    .D(\mem_rdata_latched[12] ),
    .Y(_24014_));
 sky130_fd_sc_hd__o21ai_4 _30626_ (.A1(_22361_),
    .A2(_24012_),
    .B1(_24014_),
    .Y(_00167_));
 sky130_fd_sc_hd__and4_4 _30627_ (.A(_23708_),
    .B(_18507_),
    .C(_23712_),
    .D(\mem_rdata_latched[13] ),
    .X(_24015_));
 sky130_fd_sc_hd__a21o_4 _30628_ (.A1(\decoded_imm_uj[13] ),
    .A2(_23780_),
    .B1(_24015_),
    .X(_00168_));
 sky130_fd_sc_hd__nand4_4 _30629_ (.A(_24013_),
    .B(_23748_),
    .C(_23750_),
    .D(\mem_rdata_latched[14] ),
    .Y(_24016_));
 sky130_fd_sc_hd__o21ai_4 _30630_ (.A1(_22417_),
    .A2(_24012_),
    .B1(_24016_),
    .Y(_00169_));
 sky130_fd_sc_hd__buf_1 _30631_ (.A(_23715_),
    .X(_24017_));
 sky130_fd_sc_hd__a21o_4 _30632_ (.A1(_22446_),
    .A2(_24017_),
    .B1(_23774_),
    .X(_00170_));
 sky130_fd_sc_hd__a21o_4 _30633_ (.A1(\decoded_imm_uj[16] ),
    .A2(_24017_),
    .B1(_23776_),
    .X(_00171_));
 sky130_fd_sc_hd__a21o_4 _30634_ (.A1(\decoded_imm_uj[17] ),
    .A2(_24017_),
    .B1(_23778_),
    .X(_00172_));
 sky130_fd_sc_hd__a21o_4 _30635_ (.A1(\decoded_imm_uj[18] ),
    .A2(_24017_),
    .B1(_23782_),
    .X(_00173_));
 sky130_fd_sc_hd__buf_1 _30636_ (.A(_19049_),
    .X(_24018_));
 sky130_fd_sc_hd__a21o_4 _30637_ (.A1(\decoded_imm_uj[19] ),
    .A2(_24018_),
    .B1(_23696_),
    .X(_00174_));
 sky130_vsdinv _30638_ (.A(\mem_rdata_q[7] ),
    .Y(_24019_));
 sky130_fd_sc_hd__nand3_4 _30639_ (.A(mem_rdata[7]),
    .B(_23724_),
    .C(_23725_),
    .Y(_24020_));
 sky130_fd_sc_hd__o21ai_4 _30640_ (.A1(_24019_),
    .A2(_18876_),
    .B1(_24020_),
    .Y(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__and4_4 _30641_ (.A(_23708_),
    .B(_18507_),
    .C(_23712_),
    .D(\mem_rdata_latched[7] ),
    .X(_24021_));
 sky130_fd_sc_hd__a21o_4 _30642_ (.A1(\decoded_rd[0] ),
    .A2(_24018_),
    .B1(_24021_),
    .X(_00196_));
 sky130_fd_sc_hd__buf_1 _30643_ (.A(_18876_),
    .X(_24022_));
 sky130_fd_sc_hd__buf_1 _30644_ (.A(_23724_),
    .X(_24023_));
 sky130_fd_sc_hd__buf_1 _30645_ (.A(_23725_),
    .X(_24024_));
 sky130_fd_sc_hd__nand3_4 _30646_ (.A(mem_rdata[8]),
    .B(_24023_),
    .C(_24024_),
    .Y(_24025_));
 sky130_fd_sc_hd__o21ai_4 _30647_ (.A1(_23841_),
    .A2(_24022_),
    .B1(_24025_),
    .Y(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__buf_1 _30648_ (.A(_19051_),
    .X(_24026_));
 sky130_fd_sc_hd__buf_1 _30649_ (.A(_23692_),
    .X(_24027_));
 sky130_fd_sc_hd__nand4_4 _30650_ (.A(_24013_),
    .B(_24027_),
    .C(_23750_),
    .D(\mem_rdata_latched[8] ),
    .Y(_24028_));
 sky130_fd_sc_hd__o21ai_4 _30651_ (.A1(_19083_),
    .A2(_24026_),
    .B1(_24028_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand3_4 _30652_ (.A(mem_rdata[9]),
    .B(_24023_),
    .C(_24024_),
    .Y(_24029_));
 sky130_fd_sc_hd__o21ai_4 _30653_ (.A1(_23850_),
    .A2(_24022_),
    .B1(_24029_),
    .Y(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__nand4_4 _30654_ (.A(_24013_),
    .B(_24027_),
    .C(_23740_),
    .D(\mem_rdata_latched[9] ),
    .Y(_24030_));
 sky130_fd_sc_hd__o21ai_4 _30655_ (.A1(_19088_),
    .A2(_24026_),
    .B1(_24030_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand3_4 _30656_ (.A(mem_rdata[10]),
    .B(_24023_),
    .C(_24024_),
    .Y(_24031_));
 sky130_fd_sc_hd__o21ai_4 _30657_ (.A1(_23855_),
    .A2(_24022_),
    .B1(_24031_),
    .Y(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__nand4_4 _30658_ (.A(_23097_),
    .B(_24027_),
    .C(_23740_),
    .D(\mem_rdata_latched[10] ),
    .Y(_24032_));
 sky130_fd_sc_hd__o21ai_4 _30659_ (.A1(_19093_),
    .A2(_24026_),
    .B1(_24032_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand3_4 _30660_ (.A(mem_rdata[11]),
    .B(_23735_),
    .C(_24024_),
    .Y(_24033_));
 sky130_fd_sc_hd__o21ai_4 _30661_ (.A1(_23860_),
    .A2(_24022_),
    .B1(_24033_),
    .Y(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__nand4_4 _30662_ (.A(_23097_),
    .B(_24027_),
    .C(_23740_),
    .D(\mem_rdata_latched[11] ),
    .Y(_24034_));
 sky130_fd_sc_hd__o21ai_4 _30663_ (.A1(_19105_),
    .A2(_24026_),
    .B1(_24034_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand4_4 _30664_ (.A(_23873_),
    .B(_23818_),
    .C(_23827_),
    .D(_23974_),
    .Y(_24035_));
 sky130_fd_sc_hd__buf_1 _30665_ (.A(_23817_),
    .X(_24036_));
 sky130_vsdinv _30666_ (.A(\mem_rdata_q[3] ),
    .Y(_24037_));
 sky130_fd_sc_hd__nor4_4 _30667_ (.A(_24037_),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[4] ),
    .D(\mem_rdata_q[6] ),
    .Y(_24038_));
 sky130_vsdinv _30668_ (.A(\mem_rdata_q[2] ),
    .Y(_24039_));
 sky130_fd_sc_hd__nand3_4 _30669_ (.A(_24039_),
    .B(\mem_rdata_q[1] ),
    .C(\mem_rdata_q[0] ),
    .Y(_24040_));
 sky130_vsdinv _30670_ (.A(_24040_),
    .Y(_24041_));
 sky130_fd_sc_hd__nand4_4 _30671_ (.A(_24036_),
    .B(_24038_),
    .C(_23815_),
    .D(_24041_),
    .Y(_24042_));
 sky130_fd_sc_hd__buf_1 _30672_ (.A(_19163_),
    .X(_24043_));
 sky130_fd_sc_hd__buf_1 _30673_ (.A(_24043_),
    .X(_24044_));
 sky130_fd_sc_hd__buf_1 _30674_ (.A(_23885_),
    .X(_24045_));
 sky130_fd_sc_hd__a2bb2o_4 _30675_ (.A1_N(_24035_),
    .A2_N(_24042_),
    .B1(_24044_),
    .B2(_24045_),
    .X(_00290_));
 sky130_fd_sc_hd__nand4_4 _30676_ (.A(_18203_),
    .B(_23700_),
    .C(_23703_),
    .D(_23718_),
    .Y(_24046_));
 sky130_fd_sc_hd__o21ai_4 _30677_ (.A1(_22103_),
    .A2(_19052_),
    .B1(_24046_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand3_4 _30678_ (.A(_23818_),
    .B(_23827_),
    .C(_23974_),
    .Y(_24047_));
 sky130_fd_sc_hd__nand2_4 _30679_ (.A(_24005_),
    .B(_23982_),
    .Y(_24048_));
 sky130_fd_sc_hd__nor3_4 _30680_ (.A(_24036_),
    .B(_24047_),
    .C(_24048_),
    .Y(_24049_));
 sky130_fd_sc_hd__a32o_4 _30681_ (.A1(_24049_),
    .A2(_24041_),
    .A3(_24038_),
    .B1(_21060_),
    .B2(_24000_),
    .X(_00267_));
 sky130_vsdinv _30682_ (.A(_19141_),
    .Y(_24050_));
 sky130_fd_sc_hd__and3_4 _30683_ (.A(_23700_),
    .B(_23703_),
    .C(_18209_),
    .X(_24051_));
 sky130_fd_sc_hd__nand3_4 _30684_ (.A(_24051_),
    .B(\mem_rdata_latched[26] ),
    .C(_23706_),
    .Y(_24052_));
 sky130_fd_sc_hd__o21ai_4 _30685_ (.A1(_24050_),
    .A2(_19052_),
    .B1(_24052_),
    .Y(_00274_));
 sky130_fd_sc_hd__buf_1 _30686_ (.A(decoder_pseudo_trigger),
    .X(_24053_));
 sky130_fd_sc_hd__buf_1 _30687_ (.A(_21958_),
    .X(_24054_));
 sky130_fd_sc_hd__nor3_4 _30688_ (.A(_24036_),
    .B(_24053_),
    .C(_24054_),
    .Y(_24055_));
 sky130_fd_sc_hd__nand3_4 _30689_ (.A(_24038_),
    .B(_24041_),
    .C(_24055_),
    .Y(_24056_));
 sky130_fd_sc_hd__a2bb2o_4 _30690_ (.A1_N(_24035_),
    .A2_N(_24056_),
    .B1(_19096_),
    .B2(_24045_),
    .X(_00276_));
 sky130_vsdinv _30691_ (.A(instr_getq),
    .Y(_24057_));
 sky130_fd_sc_hd__buf_1 _30692_ (.A(_23829_),
    .X(_24058_));
 sky130_fd_sc_hd__buf_1 _30693_ (.A(_24058_),
    .X(_24059_));
 sky130_fd_sc_hd__nand4_4 _30694_ (.A(_23858_),
    .B(_24038_),
    .C(_24059_),
    .D(_24041_),
    .Y(_24060_));
 sky130_fd_sc_hd__o21ai_4 _30695_ (.A1(_24057_),
    .A2(_24007_),
    .B1(_24060_),
    .Y(_00258_));
 sky130_fd_sc_hd__nor4_4 _30696_ (.A(\mem_rdata_q[8] ),
    .B(\mem_rdata_q[9] ),
    .C(\mem_rdata_q[10] ),
    .D(\mem_rdata_q[11] ),
    .Y(_24061_));
 sky130_fd_sc_hd__nor3_4 _30697_ (.A(_23900_),
    .B(_23806_),
    .C(_23823_),
    .Y(_24062_));
 sky130_fd_sc_hd__nand4_4 _30698_ (.A(_23759_),
    .B(_24061_),
    .C(_24019_),
    .D(_24062_),
    .Y(_24063_));
 sky130_fd_sc_hd__nand3_4 _30699_ (.A(_23766_),
    .B(_23768_),
    .C(_23770_),
    .Y(_24064_));
 sky130_fd_sc_hd__nor3_4 _30700_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[15] ),
    .C(_24064_),
    .Y(_24065_));
 sky130_fd_sc_hd__nor2_4 _30701_ (.A(\mem_rdata_q[22] ),
    .B(\mem_rdata_q[23] ),
    .Y(_24066_));
 sky130_fd_sc_hd__and3_4 _30702_ (.A(_23813_),
    .B(_23722_),
    .C(_24066_),
    .X(_24067_));
 sky130_fd_sc_hd__buf_1 _30703_ (.A(_24067_),
    .X(_24068_));
 sky130_fd_sc_hd__nand4_4 _30704_ (.A(_24037_),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[4] ),
    .D(\mem_rdata_q[6] ),
    .Y(_24069_));
 sky130_fd_sc_hd__nor2_4 _30705_ (.A(_24040_),
    .B(_24069_),
    .Y(_24070_));
 sky130_fd_sc_hd__nand4_4 _30706_ (.A(_24059_),
    .B(_24065_),
    .C(_24068_),
    .D(_24070_),
    .Y(_24071_));
 sky130_fd_sc_hd__a2bb2o_4 _30707_ (.A1_N(_24063_),
    .A2_N(_24071_),
    .B1(instr_ecall_ebreak),
    .B2(_24045_),
    .X(_00257_));
 sky130_fd_sc_hd__buf_1 _30708_ (.A(_18319_),
    .X(_24072_));
 sky130_fd_sc_hd__buf_1 _30709_ (.A(_24072_),
    .X(_24073_));
 sky130_fd_sc_hd__buf_1 _30710_ (.A(_24073_),
    .X(_24074_));
 sky130_fd_sc_hd__nand2_4 _30711_ (.A(_23828_),
    .B(_23759_),
    .Y(_24075_));
 sky130_fd_sc_hd__nand4_4 _30712_ (.A(_18830_),
    .B(_23820_),
    .C(_23887_),
    .D(_23890_),
    .Y(_24076_));
 sky130_fd_sc_hd__nor4_4 _30713_ (.A(_23982_),
    .B(_23876_),
    .C(_24075_),
    .D(_24076_),
    .Y(_24077_));
 sky130_fd_sc_hd__buf_1 _30714_ (.A(decoder_pseudo_trigger),
    .X(_24078_));
 sky130_fd_sc_hd__nor3_4 _30715_ (.A(\mem_rdata_q[20] ),
    .B(_24078_),
    .C(_22708_),
    .Y(_24079_));
 sky130_fd_sc_hd__and4_4 _30716_ (.A(_24077_),
    .B(\mem_rdata_q[21] ),
    .C(_24066_),
    .D(_24079_),
    .X(_24080_));
 sky130_fd_sc_hd__nor3_4 _30717_ (.A(\mem_rdata_q[12] ),
    .B(\mem_rdata_q[14] ),
    .C(_18875_),
    .Y(_24081_));
 sky130_fd_sc_hd__and3_4 _30718_ (.A(_24065_),
    .B(_24070_),
    .C(_24081_),
    .X(_24082_));
 sky130_fd_sc_hd__buf_1 _30719_ (.A(_24082_),
    .X(_24083_));
 sky130_fd_sc_hd__nand2_4 _30720_ (.A(_24080_),
    .B(_24083_),
    .Y(_24084_));
 sky130_fd_sc_hd__o21ai_4 _30721_ (.A1(_24074_),
    .A2(_24007_),
    .B1(_24084_),
    .Y(_00273_));
 sky130_fd_sc_hd__buf_1 _30722_ (.A(_18318_),
    .X(_24085_));
 sky130_fd_sc_hd__buf_1 _30723_ (.A(_24085_),
    .X(_24086_));
 sky130_fd_sc_hd__buf_1 _30724_ (.A(_24086_),
    .X(_24087_));
 sky130_fd_sc_hd__nand4_4 _30725_ (.A(_23873_),
    .B(_23876_),
    .C(_23828_),
    .D(_23762_),
    .Y(_24088_));
 sky130_fd_sc_hd__nor2_4 _30726_ (.A(_24076_),
    .B(_24088_),
    .Y(_24089_));
 sky130_fd_sc_hd__nor3_4 _30727_ (.A(\mem_rdata_q[24] ),
    .B(_24078_),
    .C(_23011_),
    .Y(_24090_));
 sky130_fd_sc_hd__and4_4 _30728_ (.A(_24089_),
    .B(\mem_rdata_q[21] ),
    .C(_24066_),
    .D(_24090_),
    .X(_24091_));
 sky130_fd_sc_hd__nand2_4 _30729_ (.A(_24091_),
    .B(_24083_),
    .Y(_24092_));
 sky130_fd_sc_hd__o21ai_4 _30730_ (.A1(_24087_),
    .A2(_24007_),
    .B1(_24092_),
    .Y(_00272_));
 sky130_fd_sc_hd__buf_1 _30731_ (.A(_18320_),
    .X(_24093_));
 sky130_fd_sc_hd__buf_1 _30732_ (.A(_24093_),
    .X(_24094_));
 sky130_fd_sc_hd__buf_1 _30733_ (.A(_24094_),
    .X(_24095_));
 sky130_fd_sc_hd__buf_1 _30734_ (.A(_24006_),
    .X(_24096_));
 sky130_fd_sc_hd__nand3_4 _30735_ (.A(_24083_),
    .B(_24068_),
    .C(_24077_),
    .Y(_24097_));
 sky130_fd_sc_hd__o21ai_4 _30736_ (.A1(_24095_),
    .A2(_24096_),
    .B1(_24097_),
    .Y(_00271_));
 sky130_fd_sc_hd__nor4_4 _30737_ (.A(_23982_),
    .B(_24036_),
    .C(_24075_),
    .D(_24076_),
    .Y(_24098_));
 sky130_fd_sc_hd__nand3_4 _30738_ (.A(_24083_),
    .B(_24068_),
    .C(_24098_),
    .Y(_24099_));
 sky130_fd_sc_hd__o21ai_4 _30739_ (.A1(_18321_),
    .A2(_24096_),
    .B1(_24099_),
    .Y(_00270_));
 sky130_fd_sc_hd__buf_1 _30740_ (.A(_23799_),
    .X(_24100_));
 sky130_fd_sc_hd__buf_1 _30741_ (.A(_24100_),
    .X(_24101_));
 sky130_fd_sc_hd__buf_1 _30742_ (.A(_23845_),
    .X(_24102_));
 sky130_fd_sc_hd__buf_1 _30743_ (.A(_24102_),
    .X(_24103_));
 sky130_fd_sc_hd__buf_1 _30744_ (.A(\mem_rdata_q[14] ),
    .X(_24104_));
 sky130_fd_sc_hd__and4_4 _30745_ (.A(_18875_),
    .B(_23900_),
    .C(_24104_),
    .D(_23792_),
    .X(_24105_));
 sky130_fd_sc_hd__nand3_4 _30746_ (.A(_23822_),
    .B(_24103_),
    .C(_24105_),
    .Y(_24106_));
 sky130_fd_sc_hd__a21bo_4 _30747_ (.A1(instr_srai),
    .A2(_24101_),
    .B1_N(_24106_),
    .X(_00285_));
 sky130_fd_sc_hd__buf_1 _30748_ (.A(_24005_),
    .X(_24107_));
 sky130_fd_sc_hd__nand3_4 _30749_ (.A(_24059_),
    .B(_24107_),
    .C(_24105_),
    .Y(_24108_));
 sky130_fd_sc_hd__a21bo_4 _30750_ (.A1(instr_srli),
    .A2(_24101_),
    .B1_N(_24108_),
    .X(_00287_));
 sky130_fd_sc_hd__buf_1 _30751_ (.A(instr_slli),
    .X(_24109_));
 sky130_fd_sc_hd__buf_1 _30752_ (.A(_24109_),
    .X(_24110_));
 sky130_fd_sc_hd__nor3_4 _30753_ (.A(_23806_),
    .B(_23823_),
    .C(_23808_),
    .Y(_24111_));
 sky130_fd_sc_hd__and4_4 _30754_ (.A(_24058_),
    .B(_23792_),
    .C(_23846_),
    .D(_24111_),
    .X(_24112_));
 sky130_fd_sc_hd__a21o_4 _30755_ (.A1(_24110_),
    .A2(_24000_),
    .B1(_24112_),
    .X(_00279_));
 sky130_fd_sc_hd__nand2_4 _30756_ (.A(_23846_),
    .B(_23837_),
    .Y(_24113_));
 sky130_vsdinv _30757_ (.A(_24081_),
    .Y(_24114_));
 sky130_fd_sc_hd__buf_1 _30758_ (.A(_23800_),
    .X(_24115_));
 sky130_fd_sc_hd__buf_1 _30759_ (.A(_24115_),
    .X(_24116_));
 sky130_fd_sc_hd__a2bb2o_4 _30760_ (.A1_N(_24113_),
    .A2_N(_24114_),
    .B1(instr_sw),
    .B2(_24116_),
    .X(_00289_));
 sky130_fd_sc_hd__buf_1 _30761_ (.A(_23853_),
    .X(_24117_));
 sky130_fd_sc_hd__buf_1 _30762_ (.A(_24111_),
    .X(_24118_));
 sky130_vsdinv _30763_ (.A(_24113_),
    .Y(_24119_));
 sky130_fd_sc_hd__a2bb2o_4 _30764_ (.A1_N(_18833_),
    .A2_N(_24117_),
    .B1(_24118_),
    .B2(_24119_),
    .X(_00277_));
 sky130_fd_sc_hd__buf_1 _30765_ (.A(_24062_),
    .X(_24120_));
 sky130_fd_sc_hd__a2bb2o_4 _30766_ (.A1_N(_18845_),
    .A2_N(_24117_),
    .B1(_24120_),
    .B2(_24119_),
    .X(_00275_));
 sky130_fd_sc_hd__nand2_4 _30767_ (.A(_23814_),
    .B(is_lb_lh_lw_lbu_lhu),
    .Y(_24121_));
 sky130_vsdinv _30768_ (.A(_24121_),
    .Y(_24122_));
 sky130_fd_sc_hd__a32o_4 _30769_ (.A1(_24122_),
    .A2(_23824_),
    .A3(_23809_),
    .B1(instr_lhu),
    .B2(_23804_),
    .X(_00264_));
 sky130_fd_sc_hd__buf_1 _30770_ (.A(\mem_rdata_q[12] ),
    .X(_24123_));
 sky130_fd_sc_hd__nor3_4 _30771_ (.A(_24123_),
    .B(_23831_),
    .C(_18878_),
    .Y(_24124_));
 sky130_vsdinv _30772_ (.A(_24124_),
    .Y(_24125_));
 sky130_fd_sc_hd__a2bb2o_4 _30773_ (.A1_N(_24121_),
    .A2_N(_24125_),
    .B1(instr_lbu),
    .B2(_24116_),
    .X(_00262_));
 sky130_fd_sc_hd__a2bb2o_4 _30774_ (.A1_N(_24121_),
    .A2_N(_24114_),
    .B1(instr_lw),
    .B2(_24116_),
    .X(_00266_));
 sky130_vsdinv _30775_ (.A(instr_lh),
    .Y(_24126_));
 sky130_fd_sc_hd__a2bb2o_4 _30776_ (.A1_N(_24126_),
    .A2_N(_24117_),
    .B1(_24118_),
    .B2(_24122_),
    .X(_00263_));
 sky130_vsdinv _30777_ (.A(_24120_),
    .Y(_24127_));
 sky130_fd_sc_hd__a2bb2o_4 _30778_ (.A1_N(_24121_),
    .A2_N(_24127_),
    .B1(instr_lb),
    .B2(_24116_),
    .X(_00261_));
 sky130_fd_sc_hd__nor3_4 _30779_ (.A(_18214_),
    .B(_18222_),
    .C(\mem_rdata_latched[4] ),
    .Y(_24128_));
 sky130_fd_sc_hd__nand4_4 _30780_ (.A(_23007_),
    .B(_24128_),
    .C(_23695_),
    .D(_23692_),
    .Y(_24129_));
 sky130_fd_sc_hd__nand4_4 _30781_ (.A(\mem_rdata_latched[2] ),
    .B(\mem_rdata_latched[1] ),
    .C(\mem_rdata_latched[0] ),
    .D(_18205_),
    .Y(_24130_));
 sky130_fd_sc_hd__or4_4 _30782_ (.A(\mem_rdata_latched[12] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[14] ),
    .D(_24130_),
    .X(_24131_));
 sky130_fd_sc_hd__a2bb2o_4 _30783_ (.A1_N(_24129_),
    .A2_N(_24131_),
    .B1(_19142_),
    .B2(_23727_),
    .X(_00260_));
 sky130_fd_sc_hd__nor4_4 _30784_ (.A(_18197_),
    .B(_18205_),
    .C(_23699_),
    .D(_24129_),
    .Y(_24132_));
 sky130_fd_sc_hd__a21o_4 _30785_ (.A1(_18777_),
    .A2(_24018_),
    .B1(_24132_),
    .X(_00259_));
 sky130_fd_sc_hd__nor4_4 _30786_ (.A(\mem_rdata_latched[5] ),
    .B(\mem_rdata_latched[6] ),
    .C(_24130_),
    .D(_23787_),
    .Y(_24133_));
 sky130_fd_sc_hd__a21o_4 _30787_ (.A1(_23912_),
    .A2(_24018_),
    .B1(_24133_),
    .X(_00250_));
 sky130_fd_sc_hd__o32ai_4 _30788_ (.A1(_23786_),
    .A2(_24130_),
    .A3(_23787_),
    .B1(_21360_),
    .B2(_19052_),
    .Y(_00265_));
 sky130_fd_sc_hd__buf_1 _30789_ (.A(_23845_),
    .X(_24134_));
 sky130_fd_sc_hd__buf_1 _30790_ (.A(_24134_),
    .X(_24135_));
 sky130_fd_sc_hd__nand2_4 _30791_ (.A(_24135_),
    .B(\mem_rdata_q[0] ),
    .Y(_24136_));
 sky130_fd_sc_hd__a21bo_4 _30792_ (.A1(pcpi_insn[0]),
    .A2(_24101_),
    .B1_N(_24136_),
    .X(_00460_));
 sky130_fd_sc_hd__nand2_4 _30793_ (.A(_24135_),
    .B(\mem_rdata_q[1] ),
    .Y(_24137_));
 sky130_fd_sc_hd__a21bo_4 _30794_ (.A1(pcpi_insn[1]),
    .A2(_24101_),
    .B1_N(_24137_),
    .X(_00471_));
 sky130_fd_sc_hd__buf_1 _30795_ (.A(_23998_),
    .X(_24138_));
 sky130_fd_sc_hd__nand2_4 _30796_ (.A(_24138_),
    .B(\mem_rdata_q[2] ),
    .Y(_24139_));
 sky130_fd_sc_hd__o21ai_4 _30797_ (.A1(_18812_),
    .A2(_24096_),
    .B1(_24139_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_4 _30798_ (.A(_24138_),
    .B(\mem_rdata_q[3] ),
    .Y(_24140_));
 sky130_fd_sc_hd__o21ai_4 _30799_ (.A1(_18811_),
    .A2(_24096_),
    .B1(_24140_),
    .Y(_00485_));
 sky130_fd_sc_hd__buf_1 _30800_ (.A(_24100_),
    .X(_24141_));
 sky130_fd_sc_hd__nand2_4 _30801_ (.A(_24135_),
    .B(\mem_rdata_q[4] ),
    .Y(_24142_));
 sky130_fd_sc_hd__a21bo_4 _30802_ (.A1(pcpi_insn[4]),
    .A2(_24141_),
    .B1_N(_24142_),
    .X(_00486_));
 sky130_fd_sc_hd__nand2_4 _30803_ (.A(_24135_),
    .B(\mem_rdata_q[5] ),
    .Y(_24143_));
 sky130_fd_sc_hd__a21bo_4 _30804_ (.A1(pcpi_insn[5]),
    .A2(_24141_),
    .B1_N(_24143_),
    .X(_00487_));
 sky130_fd_sc_hd__buf_1 _30805_ (.A(_24006_),
    .X(_24144_));
 sky130_fd_sc_hd__buf_1 _30806_ (.A(_23998_),
    .X(_24145_));
 sky130_fd_sc_hd__nand2_4 _30807_ (.A(_24145_),
    .B(\mem_rdata_q[6] ),
    .Y(_24146_));
 sky130_fd_sc_hd__o21ai_4 _30808_ (.A1(_18815_),
    .A2(_24144_),
    .B1(_24146_),
    .Y(_00488_));
 sky130_fd_sc_hd__buf_1 _30809_ (.A(_24134_),
    .X(_24147_));
 sky130_fd_sc_hd__nand2_4 _30810_ (.A(_24147_),
    .B(\mem_rdata_q[7] ),
    .Y(_24148_));
 sky130_fd_sc_hd__a21bo_4 _30811_ (.A1(pcpi_insn[7]),
    .A2(_24141_),
    .B1_N(_24148_),
    .X(_00489_));
 sky130_fd_sc_hd__nand2_4 _30812_ (.A(_24147_),
    .B(\mem_rdata_q[8] ),
    .Y(_24149_));
 sky130_fd_sc_hd__a21bo_4 _30813_ (.A1(pcpi_insn[8]),
    .A2(_24141_),
    .B1_N(_24149_),
    .X(_00490_));
 sky130_fd_sc_hd__buf_1 _30814_ (.A(_24100_),
    .X(_24150_));
 sky130_fd_sc_hd__nand2_4 _30815_ (.A(_24147_),
    .B(\mem_rdata_q[9] ),
    .Y(_24151_));
 sky130_fd_sc_hd__a21bo_4 _30816_ (.A1(pcpi_insn[9]),
    .A2(_24150_),
    .B1_N(_24151_),
    .X(_00491_));
 sky130_fd_sc_hd__nand2_4 _30817_ (.A(_24147_),
    .B(\mem_rdata_q[10] ),
    .Y(_24152_));
 sky130_fd_sc_hd__a21bo_4 _30818_ (.A1(pcpi_insn[10]),
    .A2(_24150_),
    .B1_N(_24152_),
    .X(_00461_));
 sky130_fd_sc_hd__buf_1 _30819_ (.A(_24134_),
    .X(_24153_));
 sky130_fd_sc_hd__nand2_4 _30820_ (.A(_24153_),
    .B(\mem_rdata_q[11] ),
    .Y(_24154_));
 sky130_fd_sc_hd__a21bo_4 _30821_ (.A1(pcpi_insn[11]),
    .A2(_24150_),
    .B1_N(_24154_),
    .X(_00462_));
 sky130_vsdinv _30822_ (.A(pcpi_insn[12]),
    .Y(_24155_));
 sky130_fd_sc_hd__nand2_4 _30823_ (.A(_24145_),
    .B(_24123_),
    .Y(_24156_));
 sky130_fd_sc_hd__o21ai_4 _30824_ (.A1(_24155_),
    .A2(_24144_),
    .B1(_24156_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_4 _30825_ (.A(_24153_),
    .B(_23831_),
    .Y(_24157_));
 sky130_fd_sc_hd__a21bo_4 _30826_ (.A1(pcpi_insn[13]),
    .A2(_24150_),
    .B1_N(_24157_),
    .X(_00464_));
 sky130_fd_sc_hd__nand2_4 _30827_ (.A(_24145_),
    .B(_23824_),
    .Y(_24158_));
 sky130_fd_sc_hd__o21ai_4 _30828_ (.A1(_18824_),
    .A2(_24144_),
    .B1(_24158_),
    .Y(_00465_));
 sky130_fd_sc_hd__buf_1 _30829_ (.A(_23801_),
    .X(_24159_));
 sky130_fd_sc_hd__nand2_4 _30830_ (.A(_24153_),
    .B(\mem_rdata_q[15] ),
    .Y(_24160_));
 sky130_fd_sc_hd__a21bo_4 _30831_ (.A1(pcpi_insn[15]),
    .A2(_24159_),
    .B1_N(_24160_),
    .X(_00466_));
 sky130_fd_sc_hd__nand2_4 _30832_ (.A(_24153_),
    .B(\mem_rdata_q[16] ),
    .Y(_24161_));
 sky130_fd_sc_hd__a21bo_4 _30833_ (.A1(pcpi_insn[16]),
    .A2(_24159_),
    .B1_N(_24161_),
    .X(_00467_));
 sky130_fd_sc_hd__buf_1 _30834_ (.A(_24134_),
    .X(_24162_));
 sky130_fd_sc_hd__nand2_4 _30835_ (.A(_24162_),
    .B(\mem_rdata_q[17] ),
    .Y(_24163_));
 sky130_fd_sc_hd__a21bo_4 _30836_ (.A1(pcpi_insn[17]),
    .A2(_24159_),
    .B1_N(_24163_),
    .X(_00468_));
 sky130_fd_sc_hd__nand2_4 _30837_ (.A(_24162_),
    .B(\mem_rdata_q[18] ),
    .Y(_24164_));
 sky130_fd_sc_hd__a21bo_4 _30838_ (.A1(pcpi_insn[18]),
    .A2(_24159_),
    .B1_N(_24164_),
    .X(_00469_));
 sky130_fd_sc_hd__buf_1 _30839_ (.A(_23801_),
    .X(_24165_));
 sky130_fd_sc_hd__nand2_4 _30840_ (.A(_24162_),
    .B(\mem_rdata_q[19] ),
    .Y(_24166_));
 sky130_fd_sc_hd__a21bo_4 _30841_ (.A1(pcpi_insn[19]),
    .A2(_24165_),
    .B1_N(_24166_),
    .X(_00470_));
 sky130_vsdinv _30842_ (.A(_24079_),
    .Y(_24167_));
 sky130_fd_sc_hd__o21a_4 _30843_ (.A1(pcpi_insn[20]),
    .A2(_24117_),
    .B1(_24167_),
    .X(_00472_));
 sky130_fd_sc_hd__nand2_4 _30844_ (.A(_23858_),
    .B(_23722_),
    .Y(_24168_));
 sky130_fd_sc_hd__o21a_4 _30845_ (.A1(pcpi_insn[21]),
    .A2(_24138_),
    .B1(_24168_),
    .X(_00473_));
 sky130_fd_sc_hd__nand2_4 _30846_ (.A(_24162_),
    .B(_23732_),
    .Y(_24169_));
 sky130_fd_sc_hd__a21bo_4 _30847_ (.A1(pcpi_insn[22]),
    .A2(_24165_),
    .B1_N(_24169_),
    .X(_00474_));
 sky130_fd_sc_hd__buf_1 _30848_ (.A(_24102_),
    .X(_24170_));
 sky130_fd_sc_hd__nand2_4 _30849_ (.A(_24170_),
    .B(_23742_),
    .Y(_24171_));
 sky130_fd_sc_hd__a21bo_4 _30850_ (.A1(pcpi_insn[23]),
    .A2(_24165_),
    .B1_N(_24171_),
    .X(_00475_));
 sky130_vsdinv _30851_ (.A(_24090_),
    .Y(_24172_));
 sky130_fd_sc_hd__o21a_4 _30852_ (.A1(pcpi_insn[24]),
    .A2(_24138_),
    .B1(_24172_),
    .X(_00476_));
 sky130_fd_sc_hd__nand2_4 _30853_ (.A(_24170_),
    .B(_23974_),
    .Y(_24173_));
 sky130_fd_sc_hd__a21bo_4 _30854_ (.A1(pcpi_insn[25]),
    .A2(_24165_),
    .B1_N(_24173_),
    .X(_00477_));
 sky130_fd_sc_hd__o21ai_4 _30855_ (.A1(_18816_),
    .A2(_24144_),
    .B1(_24048_),
    .Y(_00478_));
 sky130_fd_sc_hd__a21oi_4 _30856_ (.A1(_24045_),
    .A2(_18819_),
    .B1(_24055_),
    .Y(_00479_));
 sky130_fd_sc_hd__buf_1 _30857_ (.A(_24006_),
    .X(_24174_));
 sky130_fd_sc_hd__nand2_4 _30858_ (.A(_24145_),
    .B(\mem_rdata_q[28] ),
    .Y(_24175_));
 sky130_fd_sc_hd__o21ai_4 _30859_ (.A1(_18818_),
    .A2(_24174_),
    .B1(_24175_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_4 _30860_ (.A(_23847_),
    .B(_23819_),
    .Y(_24176_));
 sky130_fd_sc_hd__o21ai_4 _30861_ (.A1(_18814_),
    .A2(_24174_),
    .B1(_24176_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_4 _30862_ (.A(_23847_),
    .B(_23887_),
    .Y(_24177_));
 sky130_fd_sc_hd__o21ai_4 _30863_ (.A1(_18820_),
    .A2(_24174_),
    .B1(_24177_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_4 _30864_ (.A(_23847_),
    .B(_23890_),
    .Y(_24178_));
 sky130_fd_sc_hd__o21ai_4 _30865_ (.A1(_18823_),
    .A2(_24174_),
    .B1(_24178_),
    .Y(_00484_));
 sky130_fd_sc_hd__buf_1 _30866_ (.A(trap),
    .X(_24179_));
 sky130_fd_sc_hd__buf_1 _30867_ (.A(_24179_),
    .X(_24180_));
 sky130_fd_sc_hd__nand2_4 _30868_ (.A(_18843_),
    .B(_24180_),
    .Y(_24181_));
 sky130_fd_sc_hd__nor2_4 _30869_ (.A(_24179_),
    .B(_18227_),
    .Y(_24182_));
 sky130_fd_sc_hd__buf_1 _30870_ (.A(_24182_),
    .X(_24183_));
 sky130_fd_sc_hd__nor2_4 _30871_ (.A(_23729_),
    .B(_18254_),
    .Y(_24184_));
 sky130_fd_sc_hd__nor3_4 _30872_ (.A(_18891_),
    .B(_18892_),
    .C(_18235_),
    .Y(_24185_));
 sky130_fd_sc_hd__buf_1 _30873_ (.A(_24185_),
    .X(_24186_));
 sky130_fd_sc_hd__nor3_4 _30874_ (.A(_18280_),
    .B(_18897_),
    .C(_24186_),
    .Y(_24187_));
 sky130_fd_sc_hd__buf_1 _30875_ (.A(\mem_state[1] ),
    .X(_24188_));
 sky130_fd_sc_hd__nor2_4 _30876_ (.A(_23710_),
    .B(_21391_),
    .Y(_24189_));
 sky130_fd_sc_hd__nor2_4 _30877_ (.A(_23733_),
    .B(_24189_),
    .Y(_24190_));
 sky130_fd_sc_hd__nor3_4 _30878_ (.A(_18887_),
    .B(_24188_),
    .C(_24190_),
    .Y(_24191_));
 sky130_fd_sc_hd__or3_4 _30879_ (.A(_24184_),
    .B(_24187_),
    .C(_24191_),
    .X(_24192_));
 sky130_fd_sc_hd__a2bb2o_4 _30880_ (.A1_N(_18887_),
    .A2_N(_24181_),
    .B1(_24183_),
    .B2(_24192_),
    .X(_00421_));
 sky130_fd_sc_hd__nor3_4 _30881_ (.A(_18886_),
    .B(_24188_),
    .C(_18834_),
    .Y(_24193_));
 sky130_fd_sc_hd__nand3_4 _30882_ (.A(_23733_),
    .B(_18887_),
    .C(_24188_),
    .Y(_24194_));
 sky130_vsdinv _30883_ (.A(_24194_),
    .Y(_24195_));
 sky130_fd_sc_hd__nand4_4 _30884_ (.A(_18886_),
    .B(_23723_),
    .C(_18888_),
    .D(_24189_),
    .Y(_24196_));
 sky130_vsdinv _30885_ (.A(_24196_),
    .Y(_24197_));
 sky130_fd_sc_hd__o41ai_4 _30886_ (.A1(_24193_),
    .A2(_24184_),
    .A3(_24195_),
    .A4(_24197_),
    .B1(_24183_),
    .Y(_24198_));
 sky130_fd_sc_hd__o21ai_4 _30887_ (.A1(_18888_),
    .A2(_24181_),
    .B1(_24198_),
    .Y(_00422_));
 sky130_fd_sc_hd__a21o_4 _30888_ (.A1(_24185_),
    .A2(_18245_),
    .B1(_18896_),
    .X(_24199_));
 sky130_fd_sc_hd__nor3_4 _30889_ (.A(_18225_),
    .B(trap),
    .C(_24199_),
    .Y(_24200_));
 sky130_fd_sc_hd__buf_1 _30890_ (.A(_24200_),
    .X(_24201_));
 sky130_fd_sc_hd__buf_1 _30891_ (.A(_24201_),
    .X(_24202_));
 sky130_fd_sc_hd__buf_1 _30892_ (.A(_24202_),
    .X(_24203_));
 sky130_fd_sc_hd__buf_1 _30893_ (.A(_24183_),
    .X(_24204_));
 sky130_vsdinv _30894_ (.A(\mem_wordsize[2] ),
    .Y(_24205_));
 sky130_fd_sc_hd__nand2_4 _30895_ (.A(_24205_),
    .B(_18297_),
    .Y(_24206_));
 sky130_fd_sc_hd__nor2_4 _30896_ (.A(_18295_),
    .B(\mem_wordsize[1] ),
    .Y(_24207_));
 sky130_fd_sc_hd__a21oi_4 _30897_ (.A1(_24206_),
    .A2(_21367_),
    .B1(_24207_),
    .Y(_24208_));
 sky130_vsdinv _30898_ (.A(_24208_),
    .Y(_24209_));
 sky130_fd_sc_hd__buf_1 _30899_ (.A(_24209_),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__a211o_4 _30900_ (.A1(_24186_),
    .A2(_18246_),
    .B1(_18263_),
    .C1(_18896_),
    .X(_24210_));
 sky130_fd_sc_hd__buf_1 _30901_ (.A(_24210_),
    .X(_24211_));
 sky130_fd_sc_hd__o32ai_4 _30902_ (.A1(_18886_),
    .A2(_24188_),
    .A3(_24186_),
    .B1(mem_la_wstrb[0]),
    .B2(_24211_),
    .Y(_24212_));
 sky130_fd_sc_hd__a2bb2oi_4 _30903_ (.A1_N(mem_wstrb[0]),
    .A2_N(_24203_),
    .B1(_24204_),
    .B2(_24212_),
    .Y(_00456_));
 sky130_vsdinv _30904_ (.A(mem_wstrb[1]),
    .Y(_24213_));
 sky130_fd_sc_hd__o21ai_4 _30905_ (.A1(_18897_),
    .A2(_24186_),
    .B1(_24182_),
    .Y(_24214_));
 sky130_fd_sc_hd__buf_1 _30906_ (.A(_18227_),
    .X(_24215_));
 sky130_fd_sc_hd__buf_1 _30907_ (.A(_18841_),
    .X(_24216_));
 sky130_fd_sc_hd__buf_1 _30908_ (.A(_18620_),
    .X(_24217_));
 sky130_fd_sc_hd__buf_1 _30909_ (.A(_24217_),
    .X(_24218_));
 sky130_fd_sc_hd__buf_1 _30910_ (.A(_18841_),
    .X(_24219_));
 sky130_fd_sc_hd__nor2_4 _30911_ (.A(_24219_),
    .B(_21351_),
    .Y(_24220_));
 sky130_fd_sc_hd__o22a_4 _30912_ (.A1(_24216_),
    .A2(_18847_),
    .B1(_24218_),
    .B2(_24220_),
    .X(_24221_));
 sky130_vsdinv _30913_ (.A(_24221_),
    .Y(mem_la_wstrb[1]));
 sky130_fd_sc_hd__buf_1 _30914_ (.A(_24199_),
    .X(_24222_));
 sky130_fd_sc_hd__nor3_4 _30915_ (.A(_24215_),
    .B(mem_la_wstrb[1]),
    .C(_24222_),
    .Y(_24223_));
 sky130_fd_sc_hd__a211o_4 _30916_ (.A1(_24213_),
    .A2(_24211_),
    .B1(_24214_),
    .C1(_24223_),
    .X(_24224_));
 sky130_fd_sc_hd__o21ai_4 _30917_ (.A1(_24213_),
    .A2(_24204_),
    .B1(_24224_),
    .Y(_00457_));
 sky130_vsdinv _30918_ (.A(mem_wstrb[2]),
    .Y(_24225_));
 sky130_fd_sc_hd__buf_1 _30919_ (.A(_24206_),
    .X(_24226_));
 sky130_fd_sc_hd__buf_1 _30920_ (.A(_24207_),
    .X(_24227_));
 sky130_fd_sc_hd__buf_1 _30921_ (.A(_24227_),
    .X(_24228_));
 sky130_fd_sc_hd__buf_1 _30922_ (.A(_24228_),
    .X(_24229_));
 sky130_fd_sc_hd__a21o_4 _30923_ (.A1(_24226_),
    .A2(_21380_),
    .B1(_24229_),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__nor3_4 _30924_ (.A(_24215_),
    .B(mem_la_wstrb[2]),
    .C(_24222_),
    .Y(_24230_));
 sky130_fd_sc_hd__a211o_4 _30925_ (.A1(_24225_),
    .A2(_24210_),
    .B1(_24214_),
    .C1(_24230_),
    .X(_24231_));
 sky130_fd_sc_hd__o21ai_4 _30926_ (.A1(_24225_),
    .A2(_24204_),
    .B1(_24231_),
    .Y(_00458_));
 sky130_vsdinv _30927_ (.A(mem_wstrb[3]),
    .Y(_24232_));
 sky130_fd_sc_hd__o22a_4 _30928_ (.A1(_24216_),
    .A2(_18847_),
    .B1(_21369_),
    .B2(_24220_),
    .X(_24233_));
 sky130_vsdinv _30929_ (.A(_24233_),
    .Y(mem_la_wstrb[3]));
 sky130_fd_sc_hd__nor3_4 _30930_ (.A(_24215_),
    .B(mem_la_wstrb[3]),
    .C(_24222_),
    .Y(_24234_));
 sky130_fd_sc_hd__a211o_4 _30931_ (.A1(_24232_),
    .A2(_24210_),
    .B1(_24214_),
    .C1(_24234_),
    .X(_24235_));
 sky130_fd_sc_hd__o21ai_4 _30932_ (.A1(_24232_),
    .A2(_24204_),
    .B1(_24235_),
    .Y(_00459_));
 sky130_fd_sc_hd__buf_1 _30933_ (.A(_18661_),
    .X(_24236_));
 sky130_fd_sc_hd__buf_1 _30934_ (.A(_24228_),
    .X(_24237_));
 sky130_fd_sc_hd__buf_1 _30935_ (.A(_24237_),
    .X(_24238_));
 sky130_vsdinv _30936_ (.A(_18847_),
    .Y(_24239_));
 sky130_fd_sc_hd__buf_1 _30937_ (.A(_24239_),
    .X(_24240_));
 sky130_fd_sc_hd__buf_1 _30938_ (.A(_24240_),
    .X(_24241_));
 sky130_fd_sc_hd__a2bb2o_4 _30939_ (.A1_N(_21110_),
    .A2_N(_24241_),
    .B1(_18842_),
    .B2(_24236_),
    .X(_24242_));
 sky130_fd_sc_hd__a21o_4 _30940_ (.A1(_24236_),
    .A2(_24238_),
    .B1(_24242_),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__buf_1 _30941_ (.A(pcpi_rs2[9]),
    .X(_24243_));
 sky130_fd_sc_hd__a2bb2o_4 _30942_ (.A1_N(_21126_),
    .A2_N(_24241_),
    .B1(_18842_),
    .B2(_24243_),
    .X(_24244_));
 sky130_fd_sc_hd__a21o_4 _30943_ (.A1(_24243_),
    .A2(_24238_),
    .B1(_24244_),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__buf_1 _30944_ (.A(_21140_),
    .X(_24245_));
 sky130_fd_sc_hd__buf_1 _30945_ (.A(_24245_),
    .X(_24246_));
 sky130_fd_sc_hd__a2bb2o_4 _30946_ (.A1_N(_24246_),
    .A2_N(_24241_),
    .B1(_18842_),
    .B2(_21227_),
    .X(_24247_));
 sky130_fd_sc_hd__a21o_4 _30947_ (.A1(_21228_),
    .A2(_24238_),
    .B1(_24247_),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__buf_1 _30948_ (.A(_18658_),
    .X(_24248_));
 sky130_fd_sc_hd__buf_1 _30949_ (.A(_21153_),
    .X(_24249_));
 sky130_fd_sc_hd__buf_1 _30950_ (.A(_18841_),
    .X(_24250_));
 sky130_fd_sc_hd__a2bb2o_4 _30951_ (.A1_N(_24249_),
    .A2_N(_24241_),
    .B1(_24250_),
    .B2(_24248_),
    .X(_24251_));
 sky130_fd_sc_hd__a21o_4 _30952_ (.A1(_24248_),
    .A2(_24238_),
    .B1(_24251_),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__buf_1 _30953_ (.A(_18647_),
    .X(_24252_));
 sky130_fd_sc_hd__buf_1 _30954_ (.A(_24237_),
    .X(_01473_));
 sky130_fd_sc_hd__buf_1 _30955_ (.A(_24240_),
    .X(_01474_));
 sky130_fd_sc_hd__a2bb2o_4 _30956_ (.A1_N(_21166_),
    .A2_N(_01474_),
    .B1(_24250_),
    .B2(_24252_),
    .X(_01475_));
 sky130_fd_sc_hd__a21o_4 _30957_ (.A1(_24252_),
    .A2(_01473_),
    .B1(_01475_),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__buf_1 _30958_ (.A(pcpi_rs2[13]),
    .X(_01476_));
 sky130_fd_sc_hd__a2bb2o_4 _30959_ (.A1_N(_21179_),
    .A2_N(_01474_),
    .B1(_24250_),
    .B2(_01476_),
    .X(_01477_));
 sky130_fd_sc_hd__a21o_4 _30960_ (.A1(_01476_),
    .A2(_01473_),
    .B1(_01477_),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__buf_1 _30961_ (.A(pcpi_rs2[14]),
    .X(_01478_));
 sky130_fd_sc_hd__a2bb2o_4 _30962_ (.A1_N(_21190_),
    .A2_N(_01474_),
    .B1(_24250_),
    .B2(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__a21o_4 _30963_ (.A1(_01478_),
    .A2(_01473_),
    .B1(_01479_),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__buf_1 _30964_ (.A(_18643_),
    .X(_01480_));
 sky130_fd_sc_hd__buf_1 _30965_ (.A(_24219_),
    .X(_01481_));
 sky130_fd_sc_hd__a2bb2o_4 _30966_ (.A1_N(_21198_),
    .A2_N(_01474_),
    .B1(_01481_),
    .B2(_01480_),
    .X(_01482_));
 sky130_fd_sc_hd__a21o_4 _30967_ (.A1(_01480_),
    .A2(_01473_),
    .B1(_01482_),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__buf_1 _30968_ (.A(_24237_),
    .X(_01483_));
 sky130_fd_sc_hd__buf_1 _30969_ (.A(_24205_),
    .X(_01484_));
 sky130_fd_sc_hd__buf_1 _30970_ (.A(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__buf_1 _30971_ (.A(_01485_),
    .X(_01486_));
 sky130_fd_sc_hd__buf_1 _30972_ (.A(_24239_),
    .X(_01487_));
 sky130_fd_sc_hd__buf_1 _30973_ (.A(_01487_),
    .X(_01488_));
 sky130_fd_sc_hd__nand3_4 _30974_ (.A(_01486_),
    .B(_01488_),
    .C(_18712_),
    .Y(_01489_));
 sky130_fd_sc_hd__o21ai_4 _30975_ (.A1(_21110_),
    .A2(_01483_),
    .B1(_01489_),
    .Y(mem_la_wdata[16]));
 sky130_fd_sc_hd__nand3_4 _30976_ (.A(_01486_),
    .B(_01488_),
    .C(_18717_),
    .Y(_01490_));
 sky130_fd_sc_hd__o21ai_4 _30977_ (.A1(_21127_),
    .A2(_01483_),
    .B1(_01490_),
    .Y(mem_la_wdata[17]));
 sky130_fd_sc_hd__buf_1 _30978_ (.A(_24245_),
    .X(_01491_));
 sky130_fd_sc_hd__buf_1 _30979_ (.A(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__nand3_4 _30980_ (.A(_01486_),
    .B(_01488_),
    .C(_18706_),
    .Y(_01493_));
 sky130_fd_sc_hd__o21ai_4 _30981_ (.A1(_01492_),
    .A2(_01483_),
    .B1(_01493_),
    .Y(mem_la_wdata[18]));
 sky130_fd_sc_hd__buf_1 _30982_ (.A(_24249_),
    .X(_01494_));
 sky130_fd_sc_hd__nand3_4 _30983_ (.A(_01486_),
    .B(_01488_),
    .C(_18696_),
    .Y(_01495_));
 sky130_fd_sc_hd__o21ai_4 _30984_ (.A1(_01494_),
    .A2(_01483_),
    .B1(_01495_),
    .Y(mem_la_wdata[19]));
 sky130_fd_sc_hd__buf_1 _30985_ (.A(_24237_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_1 _30986_ (.A(_01485_),
    .X(_01497_));
 sky130_fd_sc_hd__buf_1 _30987_ (.A(_01487_),
    .X(_01498_));
 sky130_fd_sc_hd__nand3_4 _30988_ (.A(_01497_),
    .B(_01498_),
    .C(_18668_),
    .Y(_01499_));
 sky130_fd_sc_hd__o21ai_4 _30989_ (.A1(_21167_),
    .A2(_01496_),
    .B1(_01499_),
    .Y(mem_la_wdata[20]));
 sky130_fd_sc_hd__nand3_4 _30990_ (.A(_01497_),
    .B(_01498_),
    .C(_18682_),
    .Y(_01500_));
 sky130_fd_sc_hd__o21ai_4 _30991_ (.A1(_21179_),
    .A2(_01496_),
    .B1(_01500_),
    .Y(mem_la_wdata[21]));
 sky130_fd_sc_hd__nand3_4 _30992_ (.A(_01497_),
    .B(_01498_),
    .C(_18677_),
    .Y(_01501_));
 sky130_fd_sc_hd__o21ai_4 _30993_ (.A1(_21190_),
    .A2(_01496_),
    .B1(_01501_),
    .Y(mem_la_wdata[22]));
 sky130_fd_sc_hd__nand3_4 _30994_ (.A(_01497_),
    .B(_01498_),
    .C(_18689_),
    .Y(_01502_));
 sky130_fd_sc_hd__o21ai_4 _30995_ (.A1(_21198_),
    .A2(_01496_),
    .B1(_01502_),
    .Y(mem_la_wdata[23]));
 sky130_fd_sc_hd__buf_1 _30996_ (.A(_24227_),
    .X(_01503_));
 sky130_fd_sc_hd__buf_1 _30997_ (.A(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__a21o_4 _30998_ (.A1(_18734_),
    .A2(_01504_),
    .B1(_24242_),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__a21o_4 _30999_ (.A1(_18767_),
    .A2(_01504_),
    .B1(_24244_),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__a21o_4 _31000_ (.A1(_18722_),
    .A2(_01504_),
    .B1(_24247_),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__a21o_4 _31001_ (.A1(_18762_),
    .A2(_01504_),
    .B1(_24251_),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__buf_1 _31002_ (.A(_01503_),
    .X(_01505_));
 sky130_fd_sc_hd__a21o_4 _31003_ (.A1(_18747_),
    .A2(_01505_),
    .B1(_01475_),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__buf_1 _31004_ (.A(_18752_),
    .X(_01506_));
 sky130_fd_sc_hd__a21o_4 _31005_ (.A1(_01506_),
    .A2(_01505_),
    .B1(_01477_),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__a21o_4 _31006_ (.A1(_18737_),
    .A2(_01505_),
    .B1(_01479_),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__a21o_4 _31007_ (.A1(_21339_),
    .A2(_01505_),
    .B1(_01482_),
    .X(mem_la_wdata[31]));
 sky130_vsdinv _31008_ (.A(trap),
    .Y(_01507_));
 sky130_fd_sc_hd__and4_4 _31009_ (.A(_18895_),
    .B(_18374_),
    .C(_18280_),
    .D(_01507_),
    .X(_01508_));
 sky130_vsdinv _31010_ (.A(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__buf_1 _31011_ (.A(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__buf_1 _31012_ (.A(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__buf_1 _31013_ (.A(_24179_),
    .X(_01512_));
 sky130_fd_sc_hd__buf_1 _31014_ (.A(_18889_),
    .X(_01513_));
 sky130_fd_sc_hd__nor3_4 _31015_ (.A(_21110_),
    .B(_01512_),
    .C(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__a21o_4 _31016_ (.A1(_01511_),
    .A2(mem_wdata[0]),
    .B1(_01514_),
    .X(_00424_));
 sky130_fd_sc_hd__nor3_4 _31017_ (.A(_21127_),
    .B(_01512_),
    .C(_01513_),
    .Y(_01515_));
 sky130_fd_sc_hd__a21o_4 _31018_ (.A1(_01511_),
    .A2(mem_wdata[1]),
    .B1(_01515_),
    .X(_00435_));
 sky130_fd_sc_hd__buf_1 _31019_ (.A(_24179_),
    .X(_01516_));
 sky130_fd_sc_hd__nor3_4 _31020_ (.A(_21144_),
    .B(_01516_),
    .C(_01513_),
    .Y(_01517_));
 sky130_fd_sc_hd__a21o_4 _31021_ (.A1(_01511_),
    .A2(mem_wdata[2]),
    .B1(_01517_),
    .X(_00446_));
 sky130_fd_sc_hd__buf_1 _31022_ (.A(_01494_),
    .X(_01518_));
 sky130_fd_sc_hd__nor3_4 _31023_ (.A(_01518_),
    .B(_01516_),
    .C(_01513_),
    .Y(_01519_));
 sky130_fd_sc_hd__a21o_4 _31024_ (.A1(_01511_),
    .A2(mem_wdata[3]),
    .B1(_01519_),
    .X(_00449_));
 sky130_fd_sc_hd__buf_1 _31025_ (.A(_01510_),
    .X(_01520_));
 sky130_fd_sc_hd__buf_1 _31026_ (.A(_21167_),
    .X(_01521_));
 sky130_fd_sc_hd__buf_1 _31027_ (.A(_18889_),
    .X(_01522_));
 sky130_fd_sc_hd__nor3_4 _31028_ (.A(_01521_),
    .B(_01516_),
    .C(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__a21o_4 _31029_ (.A1(_01520_),
    .A2(mem_wdata[4]),
    .B1(_01523_),
    .X(_00450_));
 sky130_fd_sc_hd__nor3_4 _31030_ (.A(_21179_),
    .B(_01516_),
    .C(_01522_),
    .Y(_01524_));
 sky130_fd_sc_hd__a21o_4 _31031_ (.A1(_01520_),
    .A2(mem_wdata[5]),
    .B1(_01524_),
    .X(_00451_));
 sky130_fd_sc_hd__nor3_4 _31032_ (.A(_21190_),
    .B(_24180_),
    .C(_01522_),
    .Y(_01525_));
 sky130_fd_sc_hd__a21o_4 _31033_ (.A1(_01520_),
    .A2(mem_wdata[6]),
    .B1(_01525_),
    .X(_00452_));
 sky130_fd_sc_hd__nor3_4 _31034_ (.A(_21198_),
    .B(_24180_),
    .C(_01522_),
    .Y(_01526_));
 sky130_fd_sc_hd__a21o_4 _31035_ (.A1(_01520_),
    .A2(mem_wdata[7]),
    .B1(_01526_),
    .X(_00453_));
 sky130_fd_sc_hd__buf_1 _31036_ (.A(_01509_),
    .X(_01527_));
 sky130_fd_sc_hd__buf_1 _31037_ (.A(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__buf_1 _31038_ (.A(_01508_),
    .X(_01529_));
 sky130_fd_sc_hd__buf_1 _31039_ (.A(_01529_),
    .X(_01530_));
 sky130_fd_sc_hd__and2_4 _31040_ (.A(mem_la_wdata[8]),
    .B(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__a21o_4 _31041_ (.A1(mem_wdata[8]),
    .A2(_01528_),
    .B1(_01531_),
    .X(_00454_));
 sky130_fd_sc_hd__and2_4 _31042_ (.A(mem_la_wdata[9]),
    .B(_01530_),
    .X(_01532_));
 sky130_fd_sc_hd__a21o_4 _31043_ (.A1(mem_wdata[9]),
    .A2(_01528_),
    .B1(_01532_),
    .X(_00455_));
 sky130_fd_sc_hd__and2_4 _31044_ (.A(mem_la_wdata[10]),
    .B(_01530_),
    .X(_01533_));
 sky130_fd_sc_hd__a21o_4 _31045_ (.A1(mem_wdata[10]),
    .A2(_01528_),
    .B1(_01533_),
    .X(_00425_));
 sky130_fd_sc_hd__and2_4 _31046_ (.A(mem_la_wdata[11]),
    .B(_01530_),
    .X(_01534_));
 sky130_fd_sc_hd__a21o_4 _31047_ (.A1(mem_wdata[11]),
    .A2(_01528_),
    .B1(_01534_),
    .X(_00426_));
 sky130_fd_sc_hd__buf_1 _31048_ (.A(_01527_),
    .X(_01535_));
 sky130_fd_sc_hd__buf_1 _31049_ (.A(_01529_),
    .X(_01536_));
 sky130_fd_sc_hd__and2_4 _31050_ (.A(mem_la_wdata[12]),
    .B(_01536_),
    .X(_01537_));
 sky130_fd_sc_hd__a21o_4 _31051_ (.A1(mem_wdata[12]),
    .A2(_01535_),
    .B1(_01537_),
    .X(_00427_));
 sky130_fd_sc_hd__and2_4 _31052_ (.A(mem_la_wdata[13]),
    .B(_01536_),
    .X(_01538_));
 sky130_fd_sc_hd__a21o_4 _31053_ (.A1(mem_wdata[13]),
    .A2(_01535_),
    .B1(_01538_),
    .X(_00428_));
 sky130_fd_sc_hd__and2_4 _31054_ (.A(mem_la_wdata[14]),
    .B(_01536_),
    .X(_01539_));
 sky130_fd_sc_hd__a21o_4 _31055_ (.A1(mem_wdata[14]),
    .A2(_01535_),
    .B1(_01539_),
    .X(_00429_));
 sky130_fd_sc_hd__and2_4 _31056_ (.A(mem_la_wdata[15]),
    .B(_01536_),
    .X(_01540_));
 sky130_fd_sc_hd__a21o_4 _31057_ (.A1(mem_wdata[15]),
    .A2(_01535_),
    .B1(_01540_),
    .X(_00430_));
 sky130_fd_sc_hd__buf_1 _31058_ (.A(_01510_),
    .X(_01541_));
 sky130_fd_sc_hd__buf_1 _31059_ (.A(_01507_),
    .X(_01542_));
 sky130_fd_sc_hd__nand3_4 _31060_ (.A(mem_la_write),
    .B(mem_la_wdata[16]),
    .C(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21bo_4 _31061_ (.A1(mem_wdata[16]),
    .A2(_01541_),
    .B1_N(_01543_),
    .X(_00431_));
 sky130_fd_sc_hd__nand3_4 _31062_ (.A(mem_la_write),
    .B(mem_la_wdata[17]),
    .C(_01542_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21bo_4 _31063_ (.A1(mem_wdata[17]),
    .A2(_01541_),
    .B1_N(_01544_),
    .X(_00432_));
 sky130_fd_sc_hd__nand3_4 _31064_ (.A(mem_la_write),
    .B(mem_la_wdata[18]),
    .C(_01542_),
    .Y(_01545_));
 sky130_fd_sc_hd__a21bo_4 _31065_ (.A1(mem_wdata[18]),
    .A2(_01541_),
    .B1_N(_01545_),
    .X(_00433_));
 sky130_fd_sc_hd__buf_1 _31066_ (.A(_18890_),
    .X(_01546_));
 sky130_fd_sc_hd__nand3_4 _31067_ (.A(_01546_),
    .B(mem_la_wdata[19]),
    .C(_01542_),
    .Y(_01547_));
 sky130_fd_sc_hd__a21bo_4 _31068_ (.A1(mem_wdata[19]),
    .A2(_01541_),
    .B1_N(_01547_),
    .X(_00434_));
 sky130_fd_sc_hd__buf_1 _31069_ (.A(_01510_),
    .X(_01548_));
 sky130_fd_sc_hd__buf_1 _31070_ (.A(_01507_),
    .X(_01549_));
 sky130_fd_sc_hd__nand3_4 _31071_ (.A(_01546_),
    .B(mem_la_wdata[20]),
    .C(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__a21bo_4 _31072_ (.A1(mem_wdata[20]),
    .A2(_01548_),
    .B1_N(_01550_),
    .X(_00436_));
 sky130_fd_sc_hd__nand3_4 _31073_ (.A(_01546_),
    .B(mem_la_wdata[21]),
    .C(_01549_),
    .Y(_01551_));
 sky130_fd_sc_hd__a21bo_4 _31074_ (.A1(mem_wdata[21]),
    .A2(_01548_),
    .B1_N(_01551_),
    .X(_00437_));
 sky130_fd_sc_hd__nand3_4 _31075_ (.A(_01546_),
    .B(mem_la_wdata[22]),
    .C(_01549_),
    .Y(_01552_));
 sky130_fd_sc_hd__a21bo_4 _31076_ (.A1(mem_wdata[22]),
    .A2(_01548_),
    .B1_N(_01552_),
    .X(_00438_));
 sky130_fd_sc_hd__nand3_4 _31077_ (.A(_18890_),
    .B(mem_la_wdata[23]),
    .C(_01549_),
    .Y(_01553_));
 sky130_fd_sc_hd__a21bo_4 _31078_ (.A1(mem_wdata[23]),
    .A2(_01548_),
    .B1_N(_01553_),
    .X(_00439_));
 sky130_fd_sc_hd__buf_1 _31079_ (.A(_01527_),
    .X(_01554_));
 sky130_fd_sc_hd__buf_1 _31080_ (.A(_01529_),
    .X(_01555_));
 sky130_fd_sc_hd__and2_4 _31081_ (.A(mem_la_wdata[24]),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__a21o_4 _31082_ (.A1(mem_wdata[24]),
    .A2(_01554_),
    .B1(_01556_),
    .X(_00440_));
 sky130_fd_sc_hd__and2_4 _31083_ (.A(mem_la_wdata[25]),
    .B(_01555_),
    .X(_01557_));
 sky130_fd_sc_hd__a21o_4 _31084_ (.A1(mem_wdata[25]),
    .A2(_01554_),
    .B1(_01557_),
    .X(_00441_));
 sky130_fd_sc_hd__and2_4 _31085_ (.A(mem_la_wdata[26]),
    .B(_01555_),
    .X(_01558_));
 sky130_fd_sc_hd__a21o_4 _31086_ (.A1(mem_wdata[26]),
    .A2(_01554_),
    .B1(_01558_),
    .X(_00442_));
 sky130_fd_sc_hd__and2_4 _31087_ (.A(mem_la_wdata[27]),
    .B(_01555_),
    .X(_01559_));
 sky130_fd_sc_hd__a21o_4 _31088_ (.A1(mem_wdata[27]),
    .A2(_01554_),
    .B1(_01559_),
    .X(_00443_));
 sky130_fd_sc_hd__buf_1 _31089_ (.A(_01527_),
    .X(_01560_));
 sky130_fd_sc_hd__buf_1 _31090_ (.A(_01529_),
    .X(_01561_));
 sky130_fd_sc_hd__and2_4 _31091_ (.A(mem_la_wdata[28]),
    .B(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__a21o_4 _31092_ (.A1(mem_wdata[28]),
    .A2(_01560_),
    .B1(_01562_),
    .X(_00444_));
 sky130_fd_sc_hd__and2_4 _31093_ (.A(mem_la_wdata[29]),
    .B(_01561_),
    .X(_01563_));
 sky130_fd_sc_hd__a21o_4 _31094_ (.A1(mem_wdata[29]),
    .A2(_01560_),
    .B1(_01563_),
    .X(_00445_));
 sky130_fd_sc_hd__and2_4 _31095_ (.A(mem_la_wdata[30]),
    .B(_01561_),
    .X(_01564_));
 sky130_fd_sc_hd__a21o_4 _31096_ (.A1(mem_wdata[30]),
    .A2(_01560_),
    .B1(_01564_),
    .X(_00447_));
 sky130_fd_sc_hd__and2_4 _31097_ (.A(mem_la_wdata[31]),
    .B(_01561_),
    .X(_01565_));
 sky130_fd_sc_hd__a21o_4 _31098_ (.A1(mem_wdata[31]),
    .A2(_01560_),
    .B1(_01565_),
    .X(_00448_));
 sky130_fd_sc_hd__buf_1 _31099_ (.A(_22733_),
    .X(_01566_));
 sky130_fd_sc_hd__buf_1 _31100_ (.A(_01566_),
    .X(_01567_));
 sky130_fd_sc_hd__buf_1 _31101_ (.A(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__or2_4 _31102_ (.A(\reg_out[2] ),
    .B(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__o21ai_4 _31103_ (.A1(\reg_next_pc[2] ),
    .A2(_21919_),
    .B1(_01569_),
    .Y(_01570_));
 sky130_vsdinv _31104_ (.A(_18893_),
    .Y(_01571_));
 sky130_fd_sc_hd__buf_1 _31105_ (.A(_01571_),
    .X(_01572_));
 sky130_fd_sc_hd__buf_1 _31106_ (.A(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__buf_1 _31107_ (.A(_18891_),
    .X(_01574_));
 sky130_fd_sc_hd__buf_1 _31108_ (.A(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__nor3_4 _31109_ (.A(_01575_),
    .B(_23781_),
    .C(_21397_),
    .Y(_01576_));
 sky130_fd_sc_hd__a21oi_4 _31110_ (.A1(_01570_),
    .A2(_01573_),
    .B1(_01576_),
    .Y(mem_la_addr[2]));
 sky130_fd_sc_hd__buf_1 _31111_ (.A(_01566_),
    .X(_01577_));
 sky130_fd_sc_hd__buf_1 _31112_ (.A(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__or2_4 _31113_ (.A(\reg_out[3] ),
    .B(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__o21ai_4 _31114_ (.A1(\reg_next_pc[3] ),
    .A2(_21919_),
    .B1(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__nor3_4 _31115_ (.A(_01575_),
    .B(_23781_),
    .C(_21421_),
    .Y(_01581_));
 sky130_fd_sc_hd__a21oi_4 _31116_ (.A1(_01580_),
    .A2(_01573_),
    .B1(_01581_),
    .Y(mem_la_addr[3]));
 sky130_fd_sc_hd__or2_4 _31117_ (.A(\reg_out[4] ),
    .B(_01568_),
    .X(_01582_));
 sky130_fd_sc_hd__a21oi_4 _31118_ (.A1(_01582_),
    .A2(_22090_),
    .B1(_18893_),
    .Y(_01583_));
 sky130_fd_sc_hd__a21oi_4 _31119_ (.A1(_21435_),
    .A2(_18893_),
    .B1(_01583_),
    .Y(mem_la_addr[4]));
 sky130_fd_sc_hd__or2_4 _31120_ (.A(\reg_out[5] ),
    .B(_01578_),
    .X(_01584_));
 sky130_fd_sc_hd__o21ai_4 _31121_ (.A1(\reg_next_pc[5] ),
    .A2(_21919_),
    .B1(_01584_),
    .Y(_01585_));
 sky130_fd_sc_hd__nor3_4 _31122_ (.A(_01575_),
    .B(_23781_),
    .C(_21462_),
    .Y(_01586_));
 sky130_fd_sc_hd__a21oi_4 _31123_ (.A1(_01585_),
    .A2(_01573_),
    .B1(_01586_),
    .Y(mem_la_addr[5]));
 sky130_fd_sc_hd__buf_1 _31124_ (.A(_21918_),
    .X(_01587_));
 sky130_fd_sc_hd__or2_4 _31125_ (.A(\reg_out[6] ),
    .B(_01578_),
    .X(_01588_));
 sky130_fd_sc_hd__o21ai_4 _31126_ (.A1(\reg_next_pc[6] ),
    .A2(_01587_),
    .B1(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__buf_1 _31127_ (.A(_01572_),
    .X(_01590_));
 sky130_fd_sc_hd__buf_1 _31128_ (.A(_19048_),
    .X(_01591_));
 sky130_fd_sc_hd__nor3_4 _31129_ (.A(_01575_),
    .B(_01591_),
    .C(_21479_),
    .Y(_01592_));
 sky130_fd_sc_hd__a21oi_4 _31130_ (.A1(_01589_),
    .A2(_01590_),
    .B1(_01592_),
    .Y(mem_la_addr[6]));
 sky130_fd_sc_hd__or2_4 _31131_ (.A(\reg_out[7] ),
    .B(_01578_),
    .X(_01593_));
 sky130_fd_sc_hd__o21ai_4 _31132_ (.A1(\reg_next_pc[7] ),
    .A2(_01587_),
    .B1(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__buf_1 _31133_ (.A(_01574_),
    .X(_01595_));
 sky130_fd_sc_hd__nor3_4 _31134_ (.A(_01595_),
    .B(_01591_),
    .C(_21493_),
    .Y(_01596_));
 sky130_fd_sc_hd__a21oi_4 _31135_ (.A1(_01594_),
    .A2(_01590_),
    .B1(_01596_),
    .Y(mem_la_addr[7]));
 sky130_fd_sc_hd__buf_1 _31136_ (.A(_01577_),
    .X(_01597_));
 sky130_fd_sc_hd__or2_4 _31137_ (.A(\reg_out[8] ),
    .B(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__o21ai_4 _31138_ (.A1(\reg_next_pc[8] ),
    .A2(_01587_),
    .B1(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__nor3_4 _31139_ (.A(_01595_),
    .B(_01591_),
    .C(_21507_),
    .Y(_01600_));
 sky130_fd_sc_hd__a21oi_4 _31140_ (.A1(_01599_),
    .A2(_01590_),
    .B1(_01600_),
    .Y(mem_la_addr[8]));
 sky130_fd_sc_hd__or2_4 _31141_ (.A(\reg_out[9] ),
    .B(_01597_),
    .X(_01601_));
 sky130_fd_sc_hd__o21ai_4 _31142_ (.A1(\reg_next_pc[9] ),
    .A2(_01587_),
    .B1(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__nor3_4 _31143_ (.A(_01595_),
    .B(_01591_),
    .C(_21530_),
    .Y(_01603_));
 sky130_fd_sc_hd__a21oi_4 _31144_ (.A1(_01602_),
    .A2(_01590_),
    .B1(_01603_),
    .Y(mem_la_addr[9]));
 sky130_fd_sc_hd__buf_1 _31145_ (.A(_21918_),
    .X(_01604_));
 sky130_fd_sc_hd__or2_4 _31146_ (.A(\reg_out[10] ),
    .B(_01597_),
    .X(_01605_));
 sky130_fd_sc_hd__o21ai_4 _31147_ (.A1(\reg_next_pc[10] ),
    .A2(_01604_),
    .B1(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__buf_1 _31148_ (.A(_01571_),
    .X(_01607_));
 sky130_fd_sc_hd__buf_1 _31149_ (.A(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__buf_1 _31150_ (.A(_23693_),
    .X(_01609_));
 sky130_fd_sc_hd__buf_1 _31151_ (.A(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__buf_1 _31152_ (.A(_21545_),
    .X(_01611_));
 sky130_fd_sc_hd__nor3_4 _31153_ (.A(_01595_),
    .B(_01610_),
    .C(_01611_),
    .Y(_01612_));
 sky130_fd_sc_hd__a21oi_4 _31154_ (.A1(_01606_),
    .A2(_01608_),
    .B1(_01612_),
    .Y(mem_la_addr[10]));
 sky130_fd_sc_hd__or2_4 _31155_ (.A(\reg_out[11] ),
    .B(_01597_),
    .X(_01613_));
 sky130_fd_sc_hd__o21ai_4 _31156_ (.A1(\reg_next_pc[11] ),
    .A2(_01604_),
    .B1(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__buf_1 _31157_ (.A(_01574_),
    .X(_01615_));
 sky130_fd_sc_hd__nor3_4 _31158_ (.A(_01615_),
    .B(_01610_),
    .C(_21565_),
    .Y(_01616_));
 sky130_fd_sc_hd__a21oi_4 _31159_ (.A1(_01614_),
    .A2(_01608_),
    .B1(_01616_),
    .Y(mem_la_addr[11]));
 sky130_fd_sc_hd__buf_1 _31160_ (.A(_01577_),
    .X(_01617_));
 sky130_fd_sc_hd__or2_4 _31161_ (.A(\reg_out[12] ),
    .B(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__o21ai_4 _31162_ (.A1(\reg_next_pc[12] ),
    .A2(_01604_),
    .B1(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__nor3_4 _31163_ (.A(_01615_),
    .B(_01610_),
    .C(_21590_),
    .Y(_01620_));
 sky130_fd_sc_hd__a21oi_4 _31164_ (.A1(_01619_),
    .A2(_01608_),
    .B1(_01620_),
    .Y(mem_la_addr[12]));
 sky130_fd_sc_hd__or2_4 _31165_ (.A(\reg_out[13] ),
    .B(_01617_),
    .X(_01621_));
 sky130_fd_sc_hd__o21ai_4 _31166_ (.A1(\reg_next_pc[13] ),
    .A2(_01604_),
    .B1(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__nor3_4 _31167_ (.A(_01615_),
    .B(_01610_),
    .C(_21605_),
    .Y(_01623_));
 sky130_fd_sc_hd__a21oi_4 _31168_ (.A1(_01622_),
    .A2(_01608_),
    .B1(_01623_),
    .Y(mem_la_addr[13]));
 sky130_fd_sc_hd__buf_1 _31169_ (.A(_21917_),
    .X(_01624_));
 sky130_fd_sc_hd__buf_1 _31170_ (.A(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__or2_4 _31171_ (.A(\reg_out[14] ),
    .B(_01617_),
    .X(_01626_));
 sky130_fd_sc_hd__o21ai_4 _31172_ (.A1(\reg_next_pc[14] ),
    .A2(_01625_),
    .B1(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__buf_1 _31173_ (.A(_01607_),
    .X(_01628_));
 sky130_fd_sc_hd__buf_1 _31174_ (.A(_01609_),
    .X(_01629_));
 sky130_fd_sc_hd__buf_1 _31175_ (.A(_18638_),
    .X(_01630_));
 sky130_fd_sc_hd__nor3_4 _31176_ (.A(_01615_),
    .B(_01629_),
    .C(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__a21oi_4 _31177_ (.A1(_01627_),
    .A2(_01628_),
    .B1(_01631_),
    .Y(mem_la_addr[14]));
 sky130_fd_sc_hd__or2_4 _31178_ (.A(\reg_out[15] ),
    .B(_01617_),
    .X(_01632_));
 sky130_fd_sc_hd__o21ai_4 _31179_ (.A1(\reg_next_pc[15] ),
    .A2(_01625_),
    .B1(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__buf_1 _31180_ (.A(_18891_),
    .X(_01634_));
 sky130_fd_sc_hd__buf_1 _31181_ (.A(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__buf_1 _31182_ (.A(_18642_),
    .X(_01636_));
 sky130_fd_sc_hd__nor3_4 _31183_ (.A(_01635_),
    .B(_01629_),
    .C(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21oi_4 _31184_ (.A1(_01633_),
    .A2(_01628_),
    .B1(_01637_),
    .Y(mem_la_addr[15]));
 sky130_fd_sc_hd__buf_1 _31185_ (.A(_01577_),
    .X(_01638_));
 sky130_fd_sc_hd__or2_4 _31186_ (.A(\reg_out[16] ),
    .B(_01638_),
    .X(_01639_));
 sky130_fd_sc_hd__o21ai_4 _31187_ (.A1(\reg_next_pc[16] ),
    .A2(_01625_),
    .B1(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__nor3_4 _31188_ (.A(_01635_),
    .B(_01629_),
    .C(_21678_),
    .Y(_01641_));
 sky130_fd_sc_hd__a21oi_4 _31189_ (.A1(_01640_),
    .A2(_01628_),
    .B1(_01641_),
    .Y(mem_la_addr[16]));
 sky130_fd_sc_hd__or2_4 _31190_ (.A(\reg_out[17] ),
    .B(_01638_),
    .X(_01642_));
 sky130_fd_sc_hd__o21ai_4 _31191_ (.A1(\reg_next_pc[17] ),
    .A2(_01625_),
    .B1(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__nor3_4 _31192_ (.A(_01635_),
    .B(_01629_),
    .C(_18715_),
    .Y(_01644_));
 sky130_fd_sc_hd__a21oi_4 _31193_ (.A1(_01643_),
    .A2(_01628_),
    .B1(_01644_),
    .Y(mem_la_addr[17]));
 sky130_fd_sc_hd__buf_1 _31194_ (.A(_01624_),
    .X(_01645_));
 sky130_fd_sc_hd__or2_4 _31195_ (.A(\reg_out[18] ),
    .B(_01638_),
    .X(_01646_));
 sky130_fd_sc_hd__o21ai_4 _31196_ (.A1(\reg_next_pc[18] ),
    .A2(_01645_),
    .B1(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__buf_1 _31197_ (.A(_01607_),
    .X(_01648_));
 sky130_fd_sc_hd__buf_1 _31198_ (.A(_01609_),
    .X(_01649_));
 sky130_fd_sc_hd__nor3_4 _31199_ (.A(_01635_),
    .B(_01649_),
    .C(_18705_),
    .Y(_01650_));
 sky130_fd_sc_hd__a21oi_4 _31200_ (.A1(_01647_),
    .A2(_01648_),
    .B1(_01650_),
    .Y(mem_la_addr[18]));
 sky130_fd_sc_hd__or2_4 _31201_ (.A(\reg_out[19] ),
    .B(_01638_),
    .X(_01651_));
 sky130_fd_sc_hd__o21ai_4 _31202_ (.A1(\reg_next_pc[19] ),
    .A2(_01645_),
    .B1(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__buf_1 _31203_ (.A(_01634_),
    .X(_01653_));
 sky130_fd_sc_hd__nor3_4 _31204_ (.A(_01653_),
    .B(_01649_),
    .C(_18694_),
    .Y(_01654_));
 sky130_fd_sc_hd__a21oi_4 _31205_ (.A1(_01652_),
    .A2(_01648_),
    .B1(_01654_),
    .Y(mem_la_addr[19]));
 sky130_fd_sc_hd__buf_1 _31206_ (.A(_01566_),
    .X(_01655_));
 sky130_fd_sc_hd__or2_4 _31207_ (.A(\reg_out[20] ),
    .B(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__o21ai_4 _31208_ (.A1(\reg_next_pc[20] ),
    .A2(_01645_),
    .B1(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__nor3_4 _31209_ (.A(_01653_),
    .B(_01649_),
    .C(_21721_),
    .Y(_01658_));
 sky130_fd_sc_hd__a21oi_4 _31210_ (.A1(_01657_),
    .A2(_01648_),
    .B1(_01658_),
    .Y(mem_la_addr[20]));
 sky130_fd_sc_hd__or2_4 _31211_ (.A(\reg_out[21] ),
    .B(_01655_),
    .X(_01659_));
 sky130_fd_sc_hd__o21ai_4 _31212_ (.A1(\reg_next_pc[21] ),
    .A2(_01645_),
    .B1(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nor3_4 _31213_ (.A(_01653_),
    .B(_01649_),
    .C(_21739_),
    .Y(_01661_));
 sky130_fd_sc_hd__a21oi_4 _31214_ (.A1(_01660_),
    .A2(_01648_),
    .B1(_01661_),
    .Y(mem_la_addr[21]));
 sky130_fd_sc_hd__buf_1 _31215_ (.A(_01624_),
    .X(_01662_));
 sky130_fd_sc_hd__or2_4 _31216_ (.A(\reg_out[22] ),
    .B(_01655_),
    .X(_01663_));
 sky130_fd_sc_hd__o21ai_4 _31217_ (.A1(\reg_next_pc[22] ),
    .A2(_01662_),
    .B1(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__buf_1 _31218_ (.A(_01607_),
    .X(_01665_));
 sky130_fd_sc_hd__buf_1 _31219_ (.A(_01609_),
    .X(_01666_));
 sky130_fd_sc_hd__nor3_4 _31220_ (.A(_01653_),
    .B(_01666_),
    .C(_18676_),
    .Y(_01667_));
 sky130_fd_sc_hd__a21oi_4 _31221_ (.A1(_01664_),
    .A2(_01665_),
    .B1(_01667_),
    .Y(mem_la_addr[22]));
 sky130_fd_sc_hd__or2_4 _31222_ (.A(\reg_out[23] ),
    .B(_01655_),
    .X(_01668_));
 sky130_fd_sc_hd__o21ai_4 _31223_ (.A1(\reg_next_pc[23] ),
    .A2(_01662_),
    .B1(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__buf_1 _31224_ (.A(_01634_),
    .X(_01670_));
 sky130_fd_sc_hd__buf_1 _31225_ (.A(_18688_),
    .X(_01671_));
 sky130_fd_sc_hd__nor3_4 _31226_ (.A(_01670_),
    .B(_01666_),
    .C(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__a21oi_4 _31227_ (.A1(_01669_),
    .A2(_01665_),
    .B1(_01672_),
    .Y(mem_la_addr[23]));
 sky130_fd_sc_hd__buf_1 _31228_ (.A(_01566_),
    .X(_01673_));
 sky130_fd_sc_hd__or2_4 _31229_ (.A(\reg_out[24] ),
    .B(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__o21ai_4 _31230_ (.A1(\reg_next_pc[24] ),
    .A2(_01662_),
    .B1(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__nor3_4 _31231_ (.A(_01670_),
    .B(_01666_),
    .C(_18732_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21oi_4 _31232_ (.A1(_01675_),
    .A2(_01665_),
    .B1(_01676_),
    .Y(mem_la_addr[24]));
 sky130_fd_sc_hd__or2_4 _31233_ (.A(\reg_out[25] ),
    .B(_01673_),
    .X(_01677_));
 sky130_fd_sc_hd__o21ai_4 _31234_ (.A1(\reg_next_pc[25] ),
    .A2(_01662_),
    .B1(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__nor3_4 _31235_ (.A(_01670_),
    .B(_01666_),
    .C(_18766_),
    .Y(_01679_));
 sky130_fd_sc_hd__a21oi_4 _31236_ (.A1(_01678_),
    .A2(_01665_),
    .B1(_01679_),
    .Y(mem_la_addr[25]));
 sky130_fd_sc_hd__buf_1 _31237_ (.A(_01624_),
    .X(_01680_));
 sky130_fd_sc_hd__or2_4 _31238_ (.A(\reg_out[26] ),
    .B(_01673_),
    .X(_01681_));
 sky130_fd_sc_hd__o21ai_4 _31239_ (.A1(\reg_next_pc[26] ),
    .A2(_01680_),
    .B1(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__buf_1 _31240_ (.A(_01571_),
    .X(_01683_));
 sky130_fd_sc_hd__buf_1 _31241_ (.A(_23693_),
    .X(_01684_));
 sky130_fd_sc_hd__nor3_4 _31242_ (.A(_01670_),
    .B(_01684_),
    .C(_18721_),
    .Y(_01685_));
 sky130_fd_sc_hd__a21oi_4 _31243_ (.A1(_01682_),
    .A2(_01683_),
    .B1(_01685_),
    .Y(mem_la_addr[26]));
 sky130_fd_sc_hd__or2_4 _31244_ (.A(\reg_out[27] ),
    .B(_01673_),
    .X(_01686_));
 sky130_fd_sc_hd__o21ai_4 _31245_ (.A1(\reg_next_pc[27] ),
    .A2(_01680_),
    .B1(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__buf_1 _31246_ (.A(_01634_),
    .X(_01688_));
 sky130_fd_sc_hd__buf_1 _31247_ (.A(_18757_),
    .X(_01689_));
 sky130_fd_sc_hd__nor3_4 _31248_ (.A(_01688_),
    .B(_01684_),
    .C(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__a21oi_4 _31249_ (.A1(_01687_),
    .A2(_01683_),
    .B1(_01690_),
    .Y(mem_la_addr[27]));
 sky130_vsdinv _31250_ (.A(\reg_next_pc[28] ),
    .Y(_01691_));
 sky130_fd_sc_hd__nor2_4 _31251_ (.A(\reg_out[28] ),
    .B(_01568_),
    .Y(_01692_));
 sky130_fd_sc_hd__a21o_4 _31252_ (.A1(_01691_),
    .A2(_01568_),
    .B1(_01692_),
    .X(_01693_));
 sky130_fd_sc_hd__buf_1 _31253_ (.A(_21833_),
    .X(_01694_));
 sky130_fd_sc_hd__nor3_4 _31254_ (.A(_01688_),
    .B(_01684_),
    .C(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__a21oi_4 _31255_ (.A1(_01693_),
    .A2(_01683_),
    .B1(_01695_),
    .Y(mem_la_addr[28]));
 sky130_fd_sc_hd__or2_4 _31256_ (.A(\reg_out[29] ),
    .B(_01567_),
    .X(_01696_));
 sky130_fd_sc_hd__o21ai_4 _31257_ (.A1(\reg_next_pc[29] ),
    .A2(_01680_),
    .B1(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor3_4 _31258_ (.A(_01688_),
    .B(_01684_),
    .C(_21879_),
    .Y(_01698_));
 sky130_fd_sc_hd__a21oi_4 _31259_ (.A1(_01697_),
    .A2(_01683_),
    .B1(_01698_),
    .Y(mem_la_addr[29]));
 sky130_fd_sc_hd__or2_4 _31260_ (.A(\reg_out[30] ),
    .B(_01567_),
    .X(_01699_));
 sky130_fd_sc_hd__o21ai_4 _31261_ (.A1(\reg_next_pc[30] ),
    .A2(_01680_),
    .B1(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__nor3_4 _31262_ (.A(_01688_),
    .B(_23694_),
    .C(_21871_),
    .Y(_01701_));
 sky130_fd_sc_hd__a21oi_4 _31263_ (.A1(_01700_),
    .A2(_01572_),
    .B1(_01701_),
    .Y(mem_la_addr[30]));
 sky130_fd_sc_hd__or2_4 _31264_ (.A(\reg_out[31] ),
    .B(_01567_),
    .X(_01702_));
 sky130_fd_sc_hd__o21ai_4 _31265_ (.A1(\reg_next_pc[31] ),
    .A2(_21918_),
    .B1(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__nor3_4 _31266_ (.A(_01574_),
    .B(_23694_),
    .C(_21905_),
    .Y(_01704_));
 sky130_fd_sc_hd__a21oi_4 _31267_ (.A1(_01703_),
    .A2(_01572_),
    .B1(_01704_),
    .Y(mem_la_addr[31]));
 sky130_fd_sc_hd__o21a_4 _31268_ (.A1(_01512_),
    .A2(_24211_),
    .B1(mem_addr[0]),
    .X(_00384_));
 sky130_fd_sc_hd__o21a_4 _31269_ (.A1(_01512_),
    .A2(_24211_),
    .B1(mem_addr[1]),
    .X(_00395_));
 sky130_vsdinv _31270_ (.A(_24201_),
    .Y(_01705_));
 sky130_fd_sc_hd__buf_1 _31271_ (.A(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__buf_1 _31272_ (.A(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__and2_4 _31273_ (.A(_24203_),
    .B(mem_la_addr[2]),
    .X(_01708_));
 sky130_fd_sc_hd__a21o_4 _31274_ (.A1(mem_addr[2]),
    .A2(_01707_),
    .B1(_01708_),
    .X(_00406_));
 sky130_fd_sc_hd__and2_4 _31275_ (.A(_24203_),
    .B(mem_la_addr[3]),
    .X(_01709_));
 sky130_fd_sc_hd__a21o_4 _31276_ (.A1(mem_addr[3]),
    .A2(_01707_),
    .B1(_01709_),
    .X(_00409_));
 sky130_fd_sc_hd__and2_4 _31277_ (.A(mem_la_addr[4]),
    .B(_24202_),
    .X(_01710_));
 sky130_fd_sc_hd__a21o_4 _31278_ (.A1(mem_addr[4]),
    .A2(_01707_),
    .B1(_01710_),
    .X(_00410_));
 sky130_fd_sc_hd__and2_4 _31279_ (.A(_24203_),
    .B(mem_la_addr[5]),
    .X(_01711_));
 sky130_fd_sc_hd__a21o_4 _31280_ (.A1(mem_addr[5]),
    .A2(_01707_),
    .B1(_01711_),
    .X(_00411_));
 sky130_fd_sc_hd__buf_1 _31281_ (.A(_01706_),
    .X(_01712_));
 sky130_fd_sc_hd__buf_1 _31282_ (.A(_24200_),
    .X(_01713_));
 sky130_fd_sc_hd__buf_1 _31283_ (.A(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__and2_4 _31284_ (.A(_01714_),
    .B(mem_la_addr[6]),
    .X(_01715_));
 sky130_fd_sc_hd__a21o_4 _31285_ (.A1(mem_addr[6]),
    .A2(_01712_),
    .B1(_01715_),
    .X(_00412_));
 sky130_fd_sc_hd__and2_4 _31286_ (.A(_01714_),
    .B(mem_la_addr[7]),
    .X(_01716_));
 sky130_fd_sc_hd__a21o_4 _31287_ (.A1(mem_addr[7]),
    .A2(_01712_),
    .B1(_01716_),
    .X(_00413_));
 sky130_fd_sc_hd__and2_4 _31288_ (.A(_01714_),
    .B(mem_la_addr[8]),
    .X(_01717_));
 sky130_fd_sc_hd__a21o_4 _31289_ (.A1(mem_addr[8]),
    .A2(_01712_),
    .B1(_01717_),
    .X(_00414_));
 sky130_fd_sc_hd__and2_4 _31290_ (.A(_01714_),
    .B(mem_la_addr[9]),
    .X(_01718_));
 sky130_fd_sc_hd__a21o_4 _31291_ (.A1(mem_addr[9]),
    .A2(_01712_),
    .B1(_01718_),
    .X(_00415_));
 sky130_fd_sc_hd__buf_1 _31292_ (.A(_01705_),
    .X(_01719_));
 sky130_fd_sc_hd__buf_1 _31293_ (.A(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__buf_1 _31294_ (.A(_01713_),
    .X(_01721_));
 sky130_fd_sc_hd__and2_4 _31295_ (.A(_01721_),
    .B(mem_la_addr[10]),
    .X(_01722_));
 sky130_fd_sc_hd__a21o_4 _31296_ (.A1(mem_addr[10]),
    .A2(_01720_),
    .B1(_01722_),
    .X(_00385_));
 sky130_fd_sc_hd__and2_4 _31297_ (.A(_01721_),
    .B(mem_la_addr[11]),
    .X(_01723_));
 sky130_fd_sc_hd__a21o_4 _31298_ (.A1(mem_addr[11]),
    .A2(_01720_),
    .B1(_01723_),
    .X(_00386_));
 sky130_fd_sc_hd__and2_4 _31299_ (.A(_01721_),
    .B(mem_la_addr[12]),
    .X(_01724_));
 sky130_fd_sc_hd__a21o_4 _31300_ (.A1(mem_addr[12]),
    .A2(_01720_),
    .B1(_01724_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_4 _31301_ (.A(_01721_),
    .B(mem_la_addr[13]),
    .X(_01725_));
 sky130_fd_sc_hd__a21o_4 _31302_ (.A1(mem_addr[13]),
    .A2(_01720_),
    .B1(_01725_),
    .X(_00388_));
 sky130_fd_sc_hd__buf_1 _31303_ (.A(_01719_),
    .X(_01726_));
 sky130_fd_sc_hd__buf_1 _31304_ (.A(_01713_),
    .X(_01727_));
 sky130_fd_sc_hd__and2_4 _31305_ (.A(_01727_),
    .B(mem_la_addr[14]),
    .X(_01728_));
 sky130_fd_sc_hd__a21o_4 _31306_ (.A1(mem_addr[14]),
    .A2(_01726_),
    .B1(_01728_),
    .X(_00389_));
 sky130_fd_sc_hd__and2_4 _31307_ (.A(_01727_),
    .B(mem_la_addr[15]),
    .X(_01729_));
 sky130_fd_sc_hd__a21o_4 _31308_ (.A1(mem_addr[15]),
    .A2(_01726_),
    .B1(_01729_),
    .X(_00390_));
 sky130_fd_sc_hd__and2_4 _31309_ (.A(_01727_),
    .B(mem_la_addr[16]),
    .X(_01730_));
 sky130_fd_sc_hd__a21o_4 _31310_ (.A1(mem_addr[16]),
    .A2(_01726_),
    .B1(_01730_),
    .X(_00391_));
 sky130_fd_sc_hd__and2_4 _31311_ (.A(_01727_),
    .B(mem_la_addr[17]),
    .X(_01731_));
 sky130_fd_sc_hd__a21o_4 _31312_ (.A1(mem_addr[17]),
    .A2(_01726_),
    .B1(_01731_),
    .X(_00392_));
 sky130_fd_sc_hd__buf_1 _31313_ (.A(_01719_),
    .X(_01732_));
 sky130_fd_sc_hd__buf_1 _31314_ (.A(_01713_),
    .X(_01733_));
 sky130_fd_sc_hd__and2_4 _31315_ (.A(_01733_),
    .B(mem_la_addr[18]),
    .X(_01734_));
 sky130_fd_sc_hd__a21o_4 _31316_ (.A1(mem_addr[18]),
    .A2(_01732_),
    .B1(_01734_),
    .X(_00393_));
 sky130_fd_sc_hd__and2_4 _31317_ (.A(_01733_),
    .B(mem_la_addr[19]),
    .X(_01735_));
 sky130_fd_sc_hd__a21o_4 _31318_ (.A1(mem_addr[19]),
    .A2(_01732_),
    .B1(_01735_),
    .X(_00394_));
 sky130_fd_sc_hd__and2_4 _31319_ (.A(_01733_),
    .B(mem_la_addr[20]),
    .X(_01736_));
 sky130_fd_sc_hd__a21o_4 _31320_ (.A1(mem_addr[20]),
    .A2(_01732_),
    .B1(_01736_),
    .X(_00396_));
 sky130_fd_sc_hd__and2_4 _31321_ (.A(_01733_),
    .B(mem_la_addr[21]),
    .X(_01737_));
 sky130_fd_sc_hd__a21o_4 _31322_ (.A1(mem_addr[21]),
    .A2(_01732_),
    .B1(_01737_),
    .X(_00397_));
 sky130_fd_sc_hd__buf_1 _31323_ (.A(_01719_),
    .X(_01738_));
 sky130_fd_sc_hd__buf_1 _31324_ (.A(_24201_),
    .X(_01739_));
 sky130_fd_sc_hd__and2_4 _31325_ (.A(_01739_),
    .B(mem_la_addr[22]),
    .X(_01740_));
 sky130_fd_sc_hd__a21o_4 _31326_ (.A1(mem_addr[22]),
    .A2(_01738_),
    .B1(_01740_),
    .X(_00398_));
 sky130_fd_sc_hd__and2_4 _31327_ (.A(_01739_),
    .B(mem_la_addr[23]),
    .X(_01741_));
 sky130_fd_sc_hd__a21o_4 _31328_ (.A1(mem_addr[23]),
    .A2(_01738_),
    .B1(_01741_),
    .X(_00399_));
 sky130_fd_sc_hd__and2_4 _31329_ (.A(_01739_),
    .B(mem_la_addr[24]),
    .X(_01742_));
 sky130_fd_sc_hd__a21o_4 _31330_ (.A1(mem_addr[24]),
    .A2(_01738_),
    .B1(_01742_),
    .X(_00400_));
 sky130_fd_sc_hd__and2_4 _31331_ (.A(_01739_),
    .B(mem_la_addr[25]),
    .X(_01743_));
 sky130_fd_sc_hd__a21o_4 _31332_ (.A1(mem_addr[25]),
    .A2(_01738_),
    .B1(_01743_),
    .X(_00401_));
 sky130_fd_sc_hd__buf_1 _31333_ (.A(_01705_),
    .X(_01744_));
 sky130_fd_sc_hd__buf_1 _31334_ (.A(_24201_),
    .X(_01745_));
 sky130_fd_sc_hd__and2_4 _31335_ (.A(_01745_),
    .B(mem_la_addr[26]),
    .X(_01746_));
 sky130_fd_sc_hd__a21o_4 _31336_ (.A1(mem_addr[26]),
    .A2(_01744_),
    .B1(_01746_),
    .X(_00402_));
 sky130_fd_sc_hd__and2_4 _31337_ (.A(_01745_),
    .B(mem_la_addr[27]),
    .X(_01747_));
 sky130_fd_sc_hd__a21o_4 _31338_ (.A1(mem_addr[27]),
    .A2(_01744_),
    .B1(_01747_),
    .X(_00403_));
 sky130_fd_sc_hd__and2_4 _31339_ (.A(_01745_),
    .B(mem_la_addr[28]),
    .X(_01748_));
 sky130_fd_sc_hd__a21o_4 _31340_ (.A1(mem_addr[28]),
    .A2(_01744_),
    .B1(_01748_),
    .X(_00404_));
 sky130_fd_sc_hd__and2_4 _31341_ (.A(_01745_),
    .B(mem_la_addr[29]),
    .X(_01749_));
 sky130_fd_sc_hd__a21o_4 _31342_ (.A1(mem_addr[29]),
    .A2(_01744_),
    .B1(_01749_),
    .X(_00405_));
 sky130_fd_sc_hd__and2_4 _31343_ (.A(_24202_),
    .B(mem_la_addr[30]),
    .X(_01750_));
 sky130_fd_sc_hd__a21o_4 _31344_ (.A1(mem_addr[30]),
    .A2(_01706_),
    .B1(_01750_),
    .X(_00407_));
 sky130_fd_sc_hd__and2_4 _31345_ (.A(_24202_),
    .B(mem_la_addr[31]),
    .X(_01751_));
 sky130_fd_sc_hd__a21o_4 _31346_ (.A1(mem_addr[31]),
    .A2(_01706_),
    .B1(_01751_),
    .X(_00408_));
 sky130_fd_sc_hd__nand3_4 _31347_ (.A(_18383_),
    .B(_24183_),
    .C(_18895_),
    .Y(_01752_));
 sky130_fd_sc_hd__and4_4 _31348_ (.A(_01573_),
    .B(_24182_),
    .C(_18834_),
    .D(_18895_),
    .X(_01753_));
 sky130_fd_sc_hd__a21o_4 _31349_ (.A1(mem_instr),
    .A2(_01752_),
    .B1(_01753_),
    .X(_00420_));
 sky130_vsdinv _31350_ (.A(_23737_),
    .Y(_01754_));
 sky130_fd_sc_hd__a21o_4 _31351_ (.A1(_18897_),
    .A2(_18254_),
    .B1(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__a21o_4 _31352_ (.A1(_24222_),
    .A2(_01755_),
    .B1(_24180_),
    .X(_01756_));
 sky130_fd_sc_hd__or2_4 _31353_ (.A(_24023_),
    .B(_01754_),
    .X(_01757_));
 sky130_fd_sc_hd__a21oi_4 _31354_ (.A1(_01756_),
    .A2(_01757_),
    .B1(_23679_),
    .Y(_00423_));
 sky130_vsdinv _31355_ (.A(\latched_rd[4] ),
    .Y(_01758_));
 sky130_fd_sc_hd__nor3_4 _31356_ (.A(_19089_),
    .B(_19094_),
    .C(_01758_),
    .Y(_01759_));
 sky130_vsdinv _31357_ (.A(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__buf_1 _31358_ (.A(_22695_),
    .X(_01761_));
 sky130_fd_sc_hd__a41oi_4 _31359_ (.A1(_19128_),
    .A2(_22093_),
    .A3(_21908_),
    .A4(_01761_),
    .B1(_18261_),
    .Y(_01762_));
 sky130_fd_sc_hd__buf_1 _31360_ (.A(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__nor3_4 _31361_ (.A(\latched_rd[2] ),
    .B(\latched_rd[3] ),
    .C(\latched_rd[4] ),
    .Y(_01764_));
 sky130_fd_sc_hd__nand3_4 _31362_ (.A(_01764_),
    .B(_19067_),
    .C(_19085_),
    .Y(_01765_));
 sky130_fd_sc_hd__buf_1 _31363_ (.A(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__nand2_4 _31364_ (.A(_01763_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__buf_1 _31365_ (.A(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__nor4_4 _31366_ (.A(_19069_),
    .B(_19087_),
    .C(_01760_),
    .D(_01768_),
    .Y(_01769_));
 sky130_vsdinv _31367_ (.A(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__buf_1 _31368_ (.A(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__buf_1 _31369_ (.A(_01771_),
    .X(_01772_));
 sky130_fd_sc_hd__buf_1 _31370_ (.A(_01760_),
    .X(_01773_));
 sky130_fd_sc_hd__nor2_4 _31371_ (.A(_22875_),
    .B(_01761_),
    .Y(_01774_));
 sky130_fd_sc_hd__o21a_4 _31372_ (.A1(_22845_),
    .A2(\reg_out[0] ),
    .B1(_01774_),
    .X(_01775_));
 sky130_fd_sc_hd__o21ai_4 _31373_ (.A1(_22844_),
    .A2(\alu_out_q[0] ),
    .B1(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__buf_1 _31374_ (.A(_01774_),
    .X(_01777_));
 sky130_vsdinv _31375_ (.A(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand3_4 _31376_ (.A(_01778_),
    .B(_21361_),
    .C(_18468_),
    .Y(_01779_));
 sky130_fd_sc_hd__o21ai_4 _31377_ (.A1(_19117_),
    .A2(\reg_next_pc[0] ),
    .B1(_18466_),
    .Y(_01780_));
 sky130_fd_sc_hd__and4_4 _31378_ (.A(_01776_),
    .B(_23455_),
    .C(_01779_),
    .D(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__buf_1 _31379_ (.A(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__buf_1 _31380_ (.A(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_1 _31381_ (.A(_01763_),
    .X(_01784_));
 sky130_fd_sc_hd__buf_1 _31382_ (.A(\latched_rd[0] ),
    .X(_01785_));
 sky130_fd_sc_hd__buf_1 _31383_ (.A(\latched_rd[1] ),
    .X(_01786_));
 sky130_fd_sc_hd__buf_1 _31384_ (.A(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__buf_1 _31385_ (.A(_01765_),
    .X(_01788_));
 sky130_fd_sc_hd__and4_4 _31386_ (.A(_01784_),
    .B(_01785_),
    .C(_01787_),
    .D(_01788_),
    .X(_01789_));
 sky130_vsdinv _31387_ (.A(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor3_4 _31388_ (.A(_01773_),
    .B(_01783_),
    .C(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__a21o_4 _31389_ (.A1(\cpuregs[19][0] ),
    .A2(_01772_),
    .B1(_01791_),
    .X(_01057_));
 sky130_fd_sc_hd__or2_4 _31390_ (.A(_01778_),
    .B(_21941_),
    .X(_01792_));
 sky130_fd_sc_hd__o21a_4 _31391_ (.A1(_22875_),
    .A2(_01761_),
    .B1(_18467_),
    .X(_01793_));
 sky130_fd_sc_hd__buf_1 _31392_ (.A(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__buf_1 _31393_ (.A(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__nand2_4 _31394_ (.A(_18304_),
    .B(_19117_),
    .Y(_01796_));
 sky130_vsdinv _31395_ (.A(\reg_pc[1] ),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_4 _31396_ (.A(_01797_),
    .B(_19118_),
    .Y(_01798_));
 sky130_fd_sc_hd__nand3_4 _31397_ (.A(_01795_),
    .B(_01796_),
    .C(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__buf_1 _31398_ (.A(_19076_),
    .X(_01800_));
 sky130_fd_sc_hd__nand2_4 _31399_ (.A(_01800_),
    .B(\reg_next_pc[1] ),
    .Y(_01801_));
 sky130_fd_sc_hd__nand4_4 _31400_ (.A(_23465_),
    .B(_01792_),
    .C(_01799_),
    .D(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__buf_1 _31401_ (.A(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__and2_4 _31402_ (.A(_01769_),
    .B(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__a21o_4 _31403_ (.A1(\cpuregs[19][1] ),
    .A2(_01772_),
    .B1(_01804_),
    .X(_01068_));
 sky130_fd_sc_hd__buf_1 _31404_ (.A(_01770_),
    .X(_01805_));
 sky130_fd_sc_hd__buf_1 _31405_ (.A(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__xor2_4 _31406_ (.A(_19117_),
    .B(_21404_),
    .X(_01807_));
 sky130_vsdinv _31407_ (.A(_01793_),
    .Y(_01808_));
 sky130_fd_sc_hd__buf_1 _31408_ (.A(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__a21oi_4 _31409_ (.A1(_01807_),
    .A2(_01796_),
    .B1(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__o21ai_4 _31410_ (.A1(_01796_),
    .A2(_01807_),
    .B1(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__buf_1 _31411_ (.A(_01777_),
    .X(_01812_));
 sky130_fd_sc_hd__buf_1 _31412_ (.A(_01812_),
    .X(_01813_));
 sky130_fd_sc_hd__nand2_4 _31413_ (.A(_21964_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nand2_4 _31414_ (.A(_01800_),
    .B(\reg_next_pc[2] ),
    .Y(_01815_));
 sky130_fd_sc_hd__and4_4 _31415_ (.A(_01811_),
    .B(_23472_),
    .C(_01814_),
    .D(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__buf_1 _31416_ (.A(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__nor2_4 _31417_ (.A(_01806_),
    .B(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__a21o_4 _31418_ (.A1(\cpuregs[19][2] ),
    .A2(_01772_),
    .B1(_01818_),
    .X(_01079_));
 sky130_fd_sc_hd__a21boi_4 _31419_ (.A1(_01797_),
    .A2(latched_compr),
    .B1_N(_21404_),
    .Y(_01819_));
 sky130_fd_sc_hd__buf_1 _31420_ (.A(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__buf_1 _31421_ (.A(_01794_),
    .X(_01821_));
 sky130_fd_sc_hd__o21ai_4 _31422_ (.A1(_21417_),
    .A2(_01820_),
    .B1(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21o_4 _31423_ (.A1(_21418_),
    .A2(_01820_),
    .B1(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__buf_1 _31424_ (.A(_01777_),
    .X(_01824_));
 sky130_fd_sc_hd__buf_1 _31425_ (.A(_01824_),
    .X(_01825_));
 sky130_fd_sc_hd__nand2_4 _31426_ (.A(_22046_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__nand2_4 _31427_ (.A(_19077_),
    .B(\reg_next_pc[3] ),
    .Y(_01827_));
 sky130_fd_sc_hd__and4_4 _31428_ (.A(_01823_),
    .B(_23477_),
    .C(_01826_),
    .D(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__buf_1 _31429_ (.A(_01828_),
    .X(_01829_));
 sky130_fd_sc_hd__nor2_4 _31430_ (.A(_01806_),
    .B(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__a21o_4 _31431_ (.A1(\cpuregs[19][3] ),
    .A2(_01772_),
    .B1(_01830_),
    .X(_01082_));
 sky130_fd_sc_hd__buf_1 _31432_ (.A(_01771_),
    .X(_01831_));
 sky130_fd_sc_hd__buf_1 _31433_ (.A(_23487_),
    .X(_01832_));
 sky130_fd_sc_hd__buf_1 _31434_ (.A(_01808_),
    .X(_01833_));
 sky130_fd_sc_hd__a21oi_4 _31435_ (.A1(_01820_),
    .A2(_21417_),
    .B1(_21441_),
    .Y(_01834_));
 sky130_fd_sc_hd__and3_4 _31436_ (.A(_01820_),
    .B(_21417_),
    .C(_21441_),
    .X(_01835_));
 sky130_fd_sc_hd__or3_4 _31437_ (.A(_01833_),
    .B(_01834_),
    .C(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__buf_1 _31438_ (.A(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__buf_1 _31439_ (.A(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__nand2_4 _31440_ (.A(_22089_),
    .B(_01813_),
    .Y(_01839_));
 sky130_fd_sc_hd__buf_1 _31441_ (.A(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__buf_1 _31442_ (.A(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__nand2_4 _31443_ (.A(_01800_),
    .B(\reg_next_pc[4] ),
    .Y(_01842_));
 sky130_fd_sc_hd__buf_1 _31444_ (.A(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__buf_1 _31445_ (.A(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__a41oi_4 _31446_ (.A1(_01832_),
    .A2(_01838_),
    .A3(_01841_),
    .A4(_01844_),
    .B1(_01806_),
    .Y(_01845_));
 sky130_fd_sc_hd__a21o_4 _31447_ (.A1(\cpuregs[19][4] ),
    .A2(_01831_),
    .B1(_01845_),
    .X(_01083_));
 sky130_fd_sc_hd__buf_1 _31448_ (.A(_23494_),
    .X(_01846_));
 sky130_fd_sc_hd__buf_1 _31449_ (.A(_01794_),
    .X(_01847_));
 sky130_fd_sc_hd__o21ai_4 _31450_ (.A1(_21457_),
    .A2(_01835_),
    .B1(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__a21o_4 _31451_ (.A1(_21458_),
    .A2(_01835_),
    .B1(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__buf_1 _31452_ (.A(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__buf_1 _31453_ (.A(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__nand2_4 _31454_ (.A(_22133_),
    .B(_01813_),
    .Y(_01852_));
 sky130_fd_sc_hd__buf_1 _31455_ (.A(_01852_),
    .X(_01853_));
 sky130_fd_sc_hd__buf_1 _31456_ (.A(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__buf_1 _31457_ (.A(_19076_),
    .X(_01855_));
 sky130_fd_sc_hd__nand2_4 _31458_ (.A(_01855_),
    .B(\reg_next_pc[5] ),
    .Y(_01856_));
 sky130_fd_sc_hd__buf_1 _31459_ (.A(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__buf_1 _31460_ (.A(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__a41oi_4 _31461_ (.A1(_01846_),
    .A2(_01851_),
    .A3(_01854_),
    .A4(_01858_),
    .B1(_01806_),
    .Y(_01859_));
 sky130_fd_sc_hd__a21o_4 _31462_ (.A1(\cpuregs[19][5] ),
    .A2(_01831_),
    .B1(_01859_),
    .X(_01084_));
 sky130_fd_sc_hd__buf_1 _31463_ (.A(_23504_),
    .X(_01860_));
 sky130_fd_sc_hd__and4_4 _31464_ (.A(_01819_),
    .B(\reg_pc[3] ),
    .C(\reg_pc[4] ),
    .D(_21457_),
    .X(_01861_));
 sky130_fd_sc_hd__buf_1 _31465_ (.A(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__o21ai_4 _31466_ (.A1(_21475_),
    .A2(_01862_),
    .B1(_01847_),
    .Y(_01863_));
 sky130_fd_sc_hd__a21o_4 _31467_ (.A1(_21475_),
    .A2(_01862_),
    .B1(_01863_),
    .X(_01864_));
 sky130_fd_sc_hd__buf_1 _31468_ (.A(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__buf_1 _31469_ (.A(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__nand2_4 _31470_ (.A(_22157_),
    .B(_01813_),
    .Y(_01867_));
 sky130_fd_sc_hd__buf_1 _31471_ (.A(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__buf_1 _31472_ (.A(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_4 _31473_ (.A(_01855_),
    .B(\reg_next_pc[6] ),
    .Y(_01870_));
 sky130_fd_sc_hd__buf_1 _31474_ (.A(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__buf_1 _31475_ (.A(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__buf_1 _31476_ (.A(_01770_),
    .X(_01873_));
 sky130_fd_sc_hd__buf_1 _31477_ (.A(_01873_),
    .X(_01874_));
 sky130_fd_sc_hd__a41oi_4 _31478_ (.A1(_01860_),
    .A2(_01866_),
    .A3(_01869_),
    .A4(_01872_),
    .B1(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21o_4 _31479_ (.A1(\cpuregs[19][6] ),
    .A2(_01831_),
    .B1(_01875_),
    .X(_01085_));
 sky130_fd_sc_hd__buf_1 _31480_ (.A(_23510_),
    .X(_01876_));
 sky130_fd_sc_hd__a21oi_4 _31481_ (.A1(_01862_),
    .A2(_21474_),
    .B1(_21489_),
    .Y(_01877_));
 sky130_fd_sc_hd__and3_4 _31482_ (.A(_01861_),
    .B(_21474_),
    .C(_21489_),
    .X(_01878_));
 sky130_fd_sc_hd__buf_1 _31483_ (.A(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__or3_4 _31484_ (.A(_01833_),
    .B(_01877_),
    .C(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__buf_1 _31485_ (.A(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__buf_1 _31486_ (.A(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_1 _31487_ (.A(_01812_),
    .X(_01883_));
 sky130_fd_sc_hd__nand2_4 _31488_ (.A(_22186_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__buf_1 _31489_ (.A(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__buf_1 _31490_ (.A(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__nand2_4 _31491_ (.A(_01855_),
    .B(\reg_next_pc[7] ),
    .Y(_01887_));
 sky130_fd_sc_hd__buf_1 _31492_ (.A(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__buf_1 _31493_ (.A(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__a41oi_4 _31494_ (.A1(_01876_),
    .A2(_01882_),
    .A3(_01886_),
    .A4(_01889_),
    .B1(_01874_),
    .Y(_01890_));
 sky130_fd_sc_hd__a21o_4 _31495_ (.A1(\cpuregs[19][7] ),
    .A2(_01831_),
    .B1(_01890_),
    .X(_01086_));
 sky130_fd_sc_hd__buf_1 _31496_ (.A(_01771_),
    .X(_01891_));
 sky130_fd_sc_hd__buf_1 _31497_ (.A(_23519_),
    .X(_01892_));
 sky130_fd_sc_hd__a41oi_4 _31498_ (.A1(_21475_),
    .A2(_01862_),
    .A3(_21490_),
    .A4(_21522_),
    .B1(_01833_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21ai_4 _31499_ (.A1(_21523_),
    .A2(_01879_),
    .B1(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__buf_1 _31500_ (.A(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__buf_1 _31501_ (.A(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__nand2_4 _31502_ (.A(_22218_),
    .B(_01883_),
    .Y(_01897_));
 sky130_fd_sc_hd__buf_1 _31503_ (.A(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__buf_1 _31504_ (.A(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__nand2_4 _31505_ (.A(_01855_),
    .B(\reg_next_pc[8] ),
    .Y(_01900_));
 sky130_fd_sc_hd__buf_1 _31506_ (.A(_01900_),
    .X(_01901_));
 sky130_fd_sc_hd__buf_1 _31507_ (.A(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__a41oi_4 _31508_ (.A1(_01892_),
    .A2(_01896_),
    .A3(_01899_),
    .A4(_01902_),
    .B1(_01874_),
    .Y(_01903_));
 sky130_fd_sc_hd__a21o_4 _31509_ (.A1(\cpuregs[19][8] ),
    .A2(_01891_),
    .B1(_01903_),
    .X(_01087_));
 sky130_fd_sc_hd__buf_1 _31510_ (.A(_23526_),
    .X(_01904_));
 sky130_fd_sc_hd__and4_4 _31511_ (.A(_01861_),
    .B(_21474_),
    .C(_21489_),
    .D(\reg_pc[8] ),
    .X(_01905_));
 sky130_fd_sc_hd__o21ai_4 _31512_ (.A1(_21541_),
    .A2(_01905_),
    .B1(_01821_),
    .Y(_01906_));
 sky130_fd_sc_hd__a21o_4 _31513_ (.A1(_21541_),
    .A2(_01905_),
    .B1(_01906_),
    .X(_01907_));
 sky130_fd_sc_hd__buf_1 _31514_ (.A(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__buf_1 _31515_ (.A(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_4 _31516_ (.A(_22250_),
    .B(_01883_),
    .Y(_01910_));
 sky130_fd_sc_hd__buf_1 _31517_ (.A(_01910_),
    .X(_01911_));
 sky130_fd_sc_hd__buf_1 _31518_ (.A(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__buf_1 _31519_ (.A(_18466_),
    .X(_01913_));
 sky130_fd_sc_hd__buf_1 _31520_ (.A(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_4 _31521_ (.A(_01914_),
    .B(\reg_next_pc[9] ),
    .Y(_01915_));
 sky130_fd_sc_hd__buf_1 _31522_ (.A(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__buf_1 _31523_ (.A(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__a41oi_4 _31524_ (.A1(_01904_),
    .A2(_01909_),
    .A3(_01912_),
    .A4(_01917_),
    .B1(_01874_),
    .Y(_01918_));
 sky130_fd_sc_hd__a21o_4 _31525_ (.A1(\cpuregs[19][9] ),
    .A2(_01891_),
    .B1(_01918_),
    .X(_01088_));
 sky130_fd_sc_hd__buf_1 _31526_ (.A(_23536_),
    .X(_01919_));
 sky130_fd_sc_hd__and2_4 _31527_ (.A(_01905_),
    .B(_21540_),
    .X(_01920_));
 sky130_fd_sc_hd__a41oi_4 _31528_ (.A1(_21522_),
    .A2(_01879_),
    .A3(_21540_),
    .A4(_21558_),
    .B1(_01808_),
    .Y(_01921_));
 sky130_fd_sc_hd__o21ai_4 _31529_ (.A1(_21559_),
    .A2(_01920_),
    .B1(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__buf_1 _31530_ (.A(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__buf_1 _31531_ (.A(_01923_),
    .X(_01924_));
 sky130_fd_sc_hd__nand2_4 _31532_ (.A(_22282_),
    .B(_01883_),
    .Y(_01925_));
 sky130_fd_sc_hd__buf_1 _31533_ (.A(_01925_),
    .X(_01926_));
 sky130_fd_sc_hd__buf_1 _31534_ (.A(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__nand2_4 _31535_ (.A(_01914_),
    .B(\reg_next_pc[10] ),
    .Y(_01928_));
 sky130_fd_sc_hd__buf_1 _31536_ (.A(_01928_),
    .X(_01929_));
 sky130_fd_sc_hd__buf_1 _31537_ (.A(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__buf_1 _31538_ (.A(_01873_),
    .X(_01931_));
 sky130_fd_sc_hd__a41oi_4 _31539_ (.A1(_01919_),
    .A2(_01924_),
    .A3(_01927_),
    .A4(_01930_),
    .B1(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__a21o_4 _31540_ (.A1(\cpuregs[19][10] ),
    .A2(_01891_),
    .B1(_01932_),
    .X(_01058_));
 sky130_fd_sc_hd__buf_1 _31541_ (.A(_23542_),
    .X(_01933_));
 sky130_fd_sc_hd__and4_4 _31542_ (.A(_01905_),
    .B(\reg_pc[9] ),
    .C(_21558_),
    .D(_21574_),
    .X(_01934_));
 sky130_fd_sc_hd__buf_1 _31543_ (.A(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__a41oi_4 _31544_ (.A1(_21522_),
    .A2(_01879_),
    .A3(_21540_),
    .A4(_21558_),
    .B1(_21574_),
    .Y(_01936_));
 sky130_fd_sc_hd__or3_4 _31545_ (.A(_01833_),
    .B(_01935_),
    .C(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__buf_1 _31546_ (.A(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__buf_1 _31547_ (.A(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__buf_1 _31548_ (.A(_01812_),
    .X(_01940_));
 sky130_fd_sc_hd__nand2_4 _31549_ (.A(_22318_),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__buf_1 _31550_ (.A(_01941_),
    .X(_01942_));
 sky130_fd_sc_hd__buf_1 _31551_ (.A(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__nand2_4 _31552_ (.A(_01914_),
    .B(\reg_next_pc[11] ),
    .Y(_01944_));
 sky130_fd_sc_hd__buf_1 _31553_ (.A(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__buf_1 _31554_ (.A(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__a41oi_4 _31555_ (.A1(_01933_),
    .A2(_01939_),
    .A3(_01943_),
    .A4(_01946_),
    .B1(_01931_),
    .Y(_01947_));
 sky130_fd_sc_hd__a21o_4 _31556_ (.A1(\cpuregs[19][11] ),
    .A2(_01891_),
    .B1(_01947_),
    .X(_01059_));
 sky130_fd_sc_hd__buf_1 _31557_ (.A(_01770_),
    .X(_01948_));
 sky130_fd_sc_hd__buf_1 _31558_ (.A(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__buf_1 _31559_ (.A(_23550_),
    .X(_01950_));
 sky130_fd_sc_hd__o21ai_4 _31560_ (.A1(_21586_),
    .A2(_01935_),
    .B1(_01821_),
    .Y(_01951_));
 sky130_fd_sc_hd__a21o_4 _31561_ (.A1(_21587_),
    .A2(_01935_),
    .B1(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__buf_1 _31562_ (.A(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__buf_1 _31563_ (.A(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__nand2_4 _31564_ (.A(_22346_),
    .B(_01940_),
    .Y(_01955_));
 sky130_fd_sc_hd__buf_1 _31565_ (.A(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__buf_1 _31566_ (.A(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__nand2_4 _31567_ (.A(_01914_),
    .B(\reg_next_pc[12] ),
    .Y(_01958_));
 sky130_fd_sc_hd__buf_1 _31568_ (.A(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__buf_1 _31569_ (.A(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__a41oi_4 _31570_ (.A1(_01950_),
    .A2(_01954_),
    .A3(_01957_),
    .A4(_01960_),
    .B1(_01931_),
    .Y(_01961_));
 sky130_fd_sc_hd__a21o_4 _31571_ (.A1(\cpuregs[19][12] ),
    .A2(_01949_),
    .B1(_01961_),
    .X(_01060_));
 sky130_fd_sc_hd__buf_1 _31572_ (.A(_23557_),
    .X(_01962_));
 sky130_fd_sc_hd__and3_4 _31573_ (.A(_01934_),
    .B(_21586_),
    .C(_21617_),
    .X(_01963_));
 sky130_vsdinv _31574_ (.A(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__a21o_4 _31575_ (.A1(_01935_),
    .A2(_21586_),
    .B1(_21617_),
    .X(_01965_));
 sky130_fd_sc_hd__nand3_4 _31576_ (.A(_01964_),
    .B(_01795_),
    .C(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__buf_1 _31577_ (.A(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__buf_1 _31578_ (.A(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__nand2_4 _31579_ (.A(_22379_),
    .B(_01940_),
    .Y(_01969_));
 sky130_fd_sc_hd__buf_1 _31580_ (.A(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__buf_1 _31581_ (.A(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__buf_1 _31582_ (.A(_01913_),
    .X(_01972_));
 sky130_fd_sc_hd__nand2_4 _31583_ (.A(_01972_),
    .B(\reg_next_pc[13] ),
    .Y(_01973_));
 sky130_fd_sc_hd__buf_1 _31584_ (.A(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__buf_1 _31585_ (.A(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__a41oi_4 _31586_ (.A1(_01962_),
    .A2(_01968_),
    .A3(_01971_),
    .A4(_01975_),
    .B1(_01931_),
    .Y(_01976_));
 sky130_fd_sc_hd__a21o_4 _31587_ (.A1(\cpuregs[19][13] ),
    .A2(_01949_),
    .B1(_01976_),
    .X(_01061_));
 sky130_fd_sc_hd__buf_1 _31588_ (.A(_23567_),
    .X(_01977_));
 sky130_fd_sc_hd__o21a_4 _31589_ (.A1(_21635_),
    .A2(_01963_),
    .B1(_01821_),
    .X(_01978_));
 sky130_fd_sc_hd__and4_4 _31590_ (.A(_01934_),
    .B(\reg_pc[12] ),
    .C(\reg_pc[13] ),
    .D(_21635_),
    .X(_01979_));
 sky130_fd_sc_hd__buf_1 _31591_ (.A(_01979_),
    .X(_01980_));
 sky130_vsdinv _31592_ (.A(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__nand2_4 _31593_ (.A(_01978_),
    .B(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__buf_1 _31594_ (.A(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__buf_1 _31595_ (.A(_01983_),
    .X(_01984_));
 sky130_fd_sc_hd__nand2_4 _31596_ (.A(_22403_),
    .B(_01940_),
    .Y(_01985_));
 sky130_fd_sc_hd__buf_1 _31597_ (.A(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__buf_1 _31598_ (.A(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__nand2_4 _31599_ (.A(_01972_),
    .B(\reg_next_pc[14] ),
    .Y(_01988_));
 sky130_fd_sc_hd__buf_1 _31600_ (.A(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__buf_1 _31601_ (.A(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__buf_1 _31602_ (.A(_01873_),
    .X(_01991_));
 sky130_fd_sc_hd__a41oi_4 _31603_ (.A1(_01977_),
    .A2(_01984_),
    .A3(_01987_),
    .A4(_01990_),
    .B1(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__a21o_4 _31604_ (.A1(\cpuregs[19][14] ),
    .A2(_01949_),
    .B1(_01992_),
    .X(_01062_));
 sky130_fd_sc_hd__buf_1 _31605_ (.A(_23573_),
    .X(_01993_));
 sky130_fd_sc_hd__and2_4 _31606_ (.A(_01980_),
    .B(_21650_),
    .X(_01994_));
 sky130_vsdinv _31607_ (.A(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__buf_1 _31608_ (.A(_01793_),
    .X(_01996_));
 sky130_fd_sc_hd__o21a_4 _31609_ (.A1(_21650_),
    .A2(_01980_),
    .B1(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_4 _31610_ (.A(_01995_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__buf_1 _31611_ (.A(_01998_),
    .X(_01999_));
 sky130_fd_sc_hd__buf_1 _31612_ (.A(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__buf_1 _31613_ (.A(_01812_),
    .X(_02001_));
 sky130_fd_sc_hd__nand2_4 _31614_ (.A(_22436_),
    .B(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__buf_1 _31615_ (.A(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__buf_1 _31616_ (.A(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__nand2_4 _31617_ (.A(_01972_),
    .B(\reg_next_pc[15] ),
    .Y(_02005_));
 sky130_fd_sc_hd__buf_1 _31618_ (.A(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__buf_1 _31619_ (.A(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__a41oi_4 _31620_ (.A1(_01993_),
    .A2(_02000_),
    .A3(_02004_),
    .A4(_02007_),
    .B1(_01991_),
    .Y(_02008_));
 sky130_fd_sc_hd__a21o_4 _31621_ (.A1(\cpuregs[19][15] ),
    .A2(_01949_),
    .B1(_02008_),
    .X(_01063_));
 sky130_fd_sc_hd__buf_1 _31622_ (.A(_01948_),
    .X(_02009_));
 sky130_fd_sc_hd__buf_1 _31623_ (.A(_23582_),
    .X(_02010_));
 sky130_fd_sc_hd__buf_1 _31624_ (.A(_01793_),
    .X(_02011_));
 sky130_fd_sc_hd__o21a_4 _31625_ (.A1(_21665_),
    .A2(_01994_),
    .B1(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__and3_4 _31626_ (.A(_01980_),
    .B(_21649_),
    .C(_21664_),
    .X(_02013_));
 sky130_vsdinv _31627_ (.A(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__nand2_4 _31628_ (.A(_02012_),
    .B(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__buf_1 _31629_ (.A(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__buf_1 _31630_ (.A(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__nand2_4 _31631_ (.A(_22465_),
    .B(_02001_),
    .Y(_02018_));
 sky130_fd_sc_hd__buf_1 _31632_ (.A(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__buf_1 _31633_ (.A(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__nand2_4 _31634_ (.A(_01972_),
    .B(\reg_next_pc[16] ),
    .Y(_02021_));
 sky130_fd_sc_hd__buf_1 _31635_ (.A(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__buf_1 _31636_ (.A(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__a41oi_4 _31637_ (.A1(_02010_),
    .A2(_02017_),
    .A3(_02020_),
    .A4(_02023_),
    .B1(_01991_),
    .Y(_02024_));
 sky130_fd_sc_hd__a21o_4 _31638_ (.A1(\cpuregs[19][16] ),
    .A2(_02009_),
    .B1(_02024_),
    .X(_01064_));
 sky130_fd_sc_hd__buf_1 _31639_ (.A(_23590_),
    .X(_02025_));
 sky130_fd_sc_hd__o21a_4 _31640_ (.A1(_21674_),
    .A2(_02013_),
    .B1(_02011_),
    .X(_02026_));
 sky130_fd_sc_hd__and4_4 _31641_ (.A(_01979_),
    .B(_21649_),
    .C(_21664_),
    .D(_21674_),
    .X(_02027_));
 sky130_fd_sc_hd__buf_1 _31642_ (.A(_02027_),
    .X(_02028_));
 sky130_vsdinv _31643_ (.A(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand2_4 _31644_ (.A(_02026_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__buf_1 _31645_ (.A(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__buf_1 _31646_ (.A(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__nand2_4 _31647_ (.A(_22500_),
    .B(_02001_),
    .Y(_02033_));
 sky130_fd_sc_hd__buf_1 _31648_ (.A(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__buf_1 _31649_ (.A(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__buf_1 _31650_ (.A(_01913_),
    .X(_02036_));
 sky130_fd_sc_hd__nand2_4 _31651_ (.A(_02036_),
    .B(\reg_next_pc[17] ),
    .Y(_02037_));
 sky130_fd_sc_hd__buf_1 _31652_ (.A(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__buf_1 _31653_ (.A(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__a41oi_4 _31654_ (.A1(_02025_),
    .A2(_02032_),
    .A3(_02035_),
    .A4(_02039_),
    .B1(_01991_),
    .Y(_02040_));
 sky130_fd_sc_hd__a21o_4 _31655_ (.A1(\cpuregs[19][17] ),
    .A2(_02009_),
    .B1(_02040_),
    .X(_01065_));
 sky130_fd_sc_hd__buf_1 _31656_ (.A(_23599_),
    .X(_02041_));
 sky130_fd_sc_hd__a21oi_4 _31657_ (.A1(_02028_),
    .A2(_21701_),
    .B1(_01809_),
    .Y(_02042_));
 sky130_fd_sc_hd__o21ai_4 _31658_ (.A1(_21701_),
    .A2(_02028_),
    .B1(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__buf_1 _31659_ (.A(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__buf_1 _31660_ (.A(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__buf_1 _31661_ (.A(_01824_),
    .X(_02046_));
 sky130_fd_sc_hd__nand2_4 _31662_ (.A(_22524_),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__buf_1 _31663_ (.A(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__buf_1 _31664_ (.A(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__nand2_4 _31665_ (.A(_19077_),
    .B(\reg_next_pc[18] ),
    .Y(_02050_));
 sky130_fd_sc_hd__buf_1 _31666_ (.A(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__buf_1 _31667_ (.A(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__buf_1 _31668_ (.A(_01805_),
    .X(_02053_));
 sky130_fd_sc_hd__a41oi_4 _31669_ (.A1(_02041_),
    .A2(_02045_),
    .A3(_02049_),
    .A4(_02052_),
    .B1(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__a21o_4 _31670_ (.A1(\cpuregs[19][18] ),
    .A2(_02009_),
    .B1(_02054_),
    .X(_01066_));
 sky130_fd_sc_hd__buf_1 _31671_ (.A(_23605_),
    .X(_02055_));
 sky130_fd_sc_hd__and2_4 _31672_ (.A(_02028_),
    .B(_21700_),
    .X(_02056_));
 sky130_fd_sc_hd__o21a_4 _31673_ (.A1(_21717_),
    .A2(_02056_),
    .B1(_02011_),
    .X(_02057_));
 sky130_fd_sc_hd__and3_4 _31674_ (.A(_02027_),
    .B(_21700_),
    .C(_21716_),
    .X(_02058_));
 sky130_vsdinv _31675_ (.A(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__nand2_4 _31676_ (.A(_02057_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__buf_1 _31677_ (.A(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__buf_1 _31678_ (.A(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__nand2_4 _31679_ (.A(_22552_),
    .B(_02001_),
    .Y(_02063_));
 sky130_fd_sc_hd__buf_1 _31680_ (.A(_02063_),
    .X(_02064_));
 sky130_fd_sc_hd__buf_1 _31681_ (.A(_02064_),
    .X(_02065_));
 sky130_fd_sc_hd__nand2_4 _31682_ (.A(_02036_),
    .B(\reg_next_pc[19] ),
    .Y(_02066_));
 sky130_fd_sc_hd__buf_1 _31683_ (.A(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__buf_1 _31684_ (.A(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__a41oi_4 _31685_ (.A1(_02055_),
    .A2(_02062_),
    .A3(_02065_),
    .A4(_02068_),
    .B1(_02053_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21o_4 _31686_ (.A1(\cpuregs[19][19] ),
    .A2(_02009_),
    .B1(_02069_),
    .X(_01067_));
 sky130_fd_sc_hd__buf_1 _31687_ (.A(_01948_),
    .X(_02070_));
 sky130_fd_sc_hd__buf_1 _31688_ (.A(_23613_),
    .X(_02071_));
 sky130_fd_sc_hd__o21a_4 _31689_ (.A1(_21735_),
    .A2(_02058_),
    .B1(_02011_),
    .X(_02072_));
 sky130_fd_sc_hd__and4_4 _31690_ (.A(_02027_),
    .B(_21700_),
    .C(_21716_),
    .D(_21735_),
    .X(_02073_));
 sky130_fd_sc_hd__buf_1 _31691_ (.A(_02073_),
    .X(_02074_));
 sky130_vsdinv _31692_ (.A(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_4 _31693_ (.A(_02072_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__buf_1 _31694_ (.A(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__buf_1 _31695_ (.A(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__buf_1 _31696_ (.A(_01777_),
    .X(_02079_));
 sky130_fd_sc_hd__nand2_4 _31697_ (.A(_22575_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__buf_1 _31698_ (.A(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__buf_1 _31699_ (.A(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__nand2_4 _31700_ (.A(_02036_),
    .B(\reg_next_pc[20] ),
    .Y(_02083_));
 sky130_fd_sc_hd__buf_1 _31701_ (.A(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__buf_1 _31702_ (.A(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__a41oi_4 _31703_ (.A1(_02071_),
    .A2(_02078_),
    .A3(_02082_),
    .A4(_02085_),
    .B1(_02053_),
    .Y(_02086_));
 sky130_fd_sc_hd__a21o_4 _31704_ (.A1(\cpuregs[19][20] ),
    .A2(_02070_),
    .B1(_02086_),
    .X(_01069_));
 sky130_fd_sc_hd__buf_1 _31705_ (.A(_23620_),
    .X(_02087_));
 sky130_fd_sc_hd__and2_4 _31706_ (.A(_02074_),
    .B(_21742_),
    .X(_02088_));
 sky130_vsdinv _31707_ (.A(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__o21a_4 _31708_ (.A1(_21743_),
    .A2(_02074_),
    .B1(_01794_),
    .X(_02090_));
 sky130_fd_sc_hd__nand2_4 _31709_ (.A(_02089_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__buf_1 _31710_ (.A(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__buf_1 _31711_ (.A(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__nand2_4 _31712_ (.A(_22610_),
    .B(_02079_),
    .Y(_02094_));
 sky130_fd_sc_hd__buf_1 _31713_ (.A(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__buf_1 _31714_ (.A(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__nand2_4 _31715_ (.A(_02036_),
    .B(\reg_next_pc[21] ),
    .Y(_02097_));
 sky130_fd_sc_hd__buf_1 _31716_ (.A(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__buf_1 _31717_ (.A(_02098_),
    .X(_02099_));
 sky130_fd_sc_hd__a41oi_4 _31718_ (.A1(_02087_),
    .A2(_02093_),
    .A3(_02096_),
    .A4(_02099_),
    .B1(_02053_),
    .Y(_02100_));
 sky130_fd_sc_hd__a21o_4 _31719_ (.A1(\cpuregs[19][21] ),
    .A2(_02070_),
    .B1(_02100_),
    .X(_01070_));
 sky130_fd_sc_hd__buf_1 _31720_ (.A(_23628_),
    .X(_02101_));
 sky130_fd_sc_hd__o21a_4 _31721_ (.A1(_21762_),
    .A2(_02088_),
    .B1(_01795_),
    .X(_02102_));
 sky130_fd_sc_hd__nand3_4 _31722_ (.A(_02073_),
    .B(_21742_),
    .C(\reg_pc[22] ),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_4 _31723_ (.A(_02102_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__buf_1 _31724_ (.A(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__buf_1 _31725_ (.A(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__nand2_4 _31726_ (.A(_22636_),
    .B(_02046_),
    .Y(_02107_));
 sky130_fd_sc_hd__buf_1 _31727_ (.A(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__buf_1 _31728_ (.A(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__buf_1 _31729_ (.A(_19076_),
    .X(_02110_));
 sky130_fd_sc_hd__nand2_4 _31730_ (.A(_02110_),
    .B(\reg_next_pc[22] ),
    .Y(_02111_));
 sky130_fd_sc_hd__buf_1 _31731_ (.A(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__buf_1 _31732_ (.A(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__buf_1 _31733_ (.A(_01805_),
    .X(_02114_));
 sky130_fd_sc_hd__a41oi_4 _31734_ (.A1(_02101_),
    .A2(_02106_),
    .A3(_02109_),
    .A4(_02113_),
    .B1(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__a21o_4 _31735_ (.A1(\cpuregs[19][22] ),
    .A2(_02070_),
    .B1(_02115_),
    .X(_01071_));
 sky130_fd_sc_hd__buf_1 _31736_ (.A(_23633_),
    .X(_02116_));
 sky130_fd_sc_hd__and4_4 _31737_ (.A(_02074_),
    .B(_21742_),
    .C(_21762_),
    .D(_21772_),
    .X(_02117_));
 sky130_vsdinv _31738_ (.A(_02117_),
    .Y(_02118_));
 sky130_vsdinv _31739_ (.A(\reg_pc[23] ),
    .Y(_02119_));
 sky130_fd_sc_hd__a21oi_4 _31740_ (.A1(_02103_),
    .A2(_02119_),
    .B1(_01809_),
    .Y(_02120_));
 sky130_fd_sc_hd__nand2_4 _31741_ (.A(_02118_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__buf_1 _31742_ (.A(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__buf_1 _31743_ (.A(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__nand2_4 _31744_ (.A(_22672_),
    .B(_02079_),
    .Y(_02124_));
 sky130_fd_sc_hd__buf_1 _31745_ (.A(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__buf_1 _31746_ (.A(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__buf_1 _31747_ (.A(_01913_),
    .X(_02127_));
 sky130_fd_sc_hd__nand2_4 _31748_ (.A(_02127_),
    .B(\reg_next_pc[23] ),
    .Y(_02128_));
 sky130_fd_sc_hd__buf_1 _31749_ (.A(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__buf_1 _31750_ (.A(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__a41oi_4 _31751_ (.A1(_02116_),
    .A2(_02123_),
    .A3(_02126_),
    .A4(_02130_),
    .B1(_02114_),
    .Y(_02131_));
 sky130_fd_sc_hd__a21o_4 _31752_ (.A1(\cpuregs[19][23] ),
    .A2(_02070_),
    .B1(_02131_),
    .X(_01072_));
 sky130_fd_sc_hd__buf_1 _31753_ (.A(_01948_),
    .X(_02132_));
 sky130_fd_sc_hd__buf_1 _31754_ (.A(_23641_),
    .X(_02133_));
 sky130_fd_sc_hd__o21a_4 _31755_ (.A1(_21788_),
    .A2(_02117_),
    .B1(_01996_),
    .X(_02134_));
 sky130_vsdinv _31756_ (.A(\reg_pc[24] ),
    .Y(_02135_));
 sky130_fd_sc_hd__nor3_4 _31757_ (.A(_02119_),
    .B(_02135_),
    .C(_02103_),
    .Y(_02136_));
 sky130_vsdinv _31758_ (.A(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_4 _31759_ (.A(_02134_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__buf_1 _31760_ (.A(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__buf_1 _31761_ (.A(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__nand2_4 _31762_ (.A(_22697_),
    .B(_02079_),
    .Y(_02141_));
 sky130_fd_sc_hd__buf_1 _31763_ (.A(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__buf_1 _31764_ (.A(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__nand2_4 _31765_ (.A(_02127_),
    .B(\reg_next_pc[24] ),
    .Y(_02144_));
 sky130_fd_sc_hd__buf_1 _31766_ (.A(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__buf_1 _31767_ (.A(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__a41oi_4 _31768_ (.A1(_02133_),
    .A2(_02140_),
    .A3(_02143_),
    .A4(_02146_),
    .B1(_02114_),
    .Y(_02147_));
 sky130_fd_sc_hd__a21o_4 _31769_ (.A1(\cpuregs[19][24] ),
    .A2(_02132_),
    .B1(_02147_),
    .X(_01073_));
 sky130_fd_sc_hd__buf_1 _31770_ (.A(_23648_),
    .X(_02148_));
 sky130_fd_sc_hd__o21a_4 _31771_ (.A1(_21796_),
    .A2(_02136_),
    .B1(_01996_),
    .X(_02149_));
 sky130_vsdinv _31772_ (.A(\reg_pc[25] ),
    .Y(_02150_));
 sky130_fd_sc_hd__nor4_4 _31773_ (.A(_02119_),
    .B(_02135_),
    .C(_02150_),
    .D(_02103_),
    .Y(_02151_));
 sky130_vsdinv _31774_ (.A(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_4 _31775_ (.A(_02149_),
    .B(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__buf_1 _31776_ (.A(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__buf_1 _31777_ (.A(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__nand2_4 _31778_ (.A(_22730_),
    .B(_01824_),
    .Y(_02156_));
 sky130_fd_sc_hd__buf_1 _31779_ (.A(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_1 _31780_ (.A(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__nand2_4 _31781_ (.A(_02127_),
    .B(\reg_next_pc[25] ),
    .Y(_02159_));
 sky130_fd_sc_hd__buf_1 _31782_ (.A(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__buf_1 _31783_ (.A(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__a41oi_4 _31784_ (.A1(_02148_),
    .A2(_02155_),
    .A3(_02158_),
    .A4(_02161_),
    .B1(_02114_),
    .Y(_02162_));
 sky130_fd_sc_hd__a21o_4 _31785_ (.A1(\cpuregs[19][25] ),
    .A2(_02132_),
    .B1(_02162_),
    .X(_01074_));
 sky130_fd_sc_hd__buf_1 _31786_ (.A(_23656_),
    .X(_02163_));
 sky130_fd_sc_hd__o21a_4 _31787_ (.A1(_21817_),
    .A2(_02151_),
    .B1(_01996_),
    .X(_02164_));
 sky130_fd_sc_hd__and4_4 _31788_ (.A(_02117_),
    .B(_21788_),
    .C(_21796_),
    .D(_21816_),
    .X(_02165_));
 sky130_vsdinv _31789_ (.A(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__nand2_4 _31790_ (.A(_02164_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__buf_1 _31791_ (.A(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__buf_1 _31792_ (.A(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_4 _31793_ (.A(_22758_),
    .B(_01824_),
    .Y(_02170_));
 sky130_fd_sc_hd__buf_1 _31794_ (.A(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__buf_1 _31795_ (.A(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__nand2_4 _31796_ (.A(_02127_),
    .B(\reg_next_pc[26] ),
    .Y(_02173_));
 sky130_fd_sc_hd__buf_1 _31797_ (.A(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__buf_1 _31798_ (.A(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__buf_1 _31799_ (.A(_01805_),
    .X(_02176_));
 sky130_fd_sc_hd__a41oi_4 _31800_ (.A1(_02163_),
    .A2(_02169_),
    .A3(_02172_),
    .A4(_02175_),
    .B1(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__a21o_4 _31801_ (.A1(\cpuregs[19][26] ),
    .A2(_02132_),
    .B1(_02177_),
    .X(_01075_));
 sky130_fd_sc_hd__buf_1 _31802_ (.A(_23662_),
    .X(_02178_));
 sky130_fd_sc_hd__o21a_4 _31803_ (.A1(_21829_),
    .A2(_02165_),
    .B1(_01847_),
    .X(_02179_));
 sky130_fd_sc_hd__and4_4 _31804_ (.A(_02136_),
    .B(\reg_pc[25] ),
    .C(_21816_),
    .D(\reg_pc[27] ),
    .X(_02180_));
 sky130_vsdinv _31805_ (.A(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_4 _31806_ (.A(_02179_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__buf_1 _31807_ (.A(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__buf_1 _31808_ (.A(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__nand2_4 _31809_ (.A(_22787_),
    .B(_02046_),
    .Y(_02185_));
 sky130_fd_sc_hd__buf_1 _31810_ (.A(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__buf_1 _31811_ (.A(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__nand2_4 _31812_ (.A(_02110_),
    .B(\reg_next_pc[27] ),
    .Y(_02188_));
 sky130_fd_sc_hd__buf_1 _31813_ (.A(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__buf_1 _31814_ (.A(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__a41oi_4 _31815_ (.A1(_02178_),
    .A2(_02184_),
    .A3(_02187_),
    .A4(_02190_),
    .B1(_02176_),
    .Y(_02191_));
 sky130_fd_sc_hd__a21o_4 _31816_ (.A1(\cpuregs[19][27] ),
    .A2(_02132_),
    .B1(_02191_),
    .X(_01076_));
 sky130_fd_sc_hd__buf_1 _31817_ (.A(_01873_),
    .X(_02192_));
 sky130_fd_sc_hd__o21ai_4 _31818_ (.A1(_22093_),
    .A2(_01691_),
    .B1(_23668_),
    .Y(_02193_));
 sky130_fd_sc_hd__buf_1 _31819_ (.A(_21849_),
    .X(_02194_));
 sky130_fd_sc_hd__a41oi_4 _31820_ (.A1(_21817_),
    .A2(_02151_),
    .A3(_21828_),
    .A4(_21849_),
    .B1(_01808_),
    .Y(_02195_));
 sky130_fd_sc_hd__o21a_4 _31821_ (.A1(_02194_),
    .A2(_02180_),
    .B1(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__a211o_4 _31822_ (.A1(_22810_),
    .A2(_02046_),
    .B1(_02193_),
    .C1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__buf_1 _31823_ (.A(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__and2_4 _31824_ (.A(_02198_),
    .B(_01769_),
    .X(_02199_));
 sky130_fd_sc_hd__a21o_4 _31825_ (.A1(\cpuregs[19][28] ),
    .A2(_02192_),
    .B1(_02199_),
    .X(_01077_));
 sky130_fd_sc_hd__buf_1 _31826_ (.A(_23674_),
    .X(_02200_));
 sky130_fd_sc_hd__and4_4 _31827_ (.A(_02151_),
    .B(_21816_),
    .C(_21828_),
    .D(\reg_pc[28] ),
    .X(_02201_));
 sky130_fd_sc_hd__buf_1 _31828_ (.A(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__o21ai_4 _31829_ (.A1(_21863_),
    .A2(_02202_),
    .B1(_01795_),
    .Y(_02203_));
 sky130_fd_sc_hd__a21o_4 _31830_ (.A1(_21864_),
    .A2(_02202_),
    .B1(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__buf_1 _31831_ (.A(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__buf_1 _31832_ (.A(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__nand2_4 _31833_ (.A(_22847_),
    .B(_01825_),
    .Y(_02207_));
 sky130_fd_sc_hd__buf_1 _31834_ (.A(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__buf_1 _31835_ (.A(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__nand2_4 _31836_ (.A(_02110_),
    .B(\reg_next_pc[29] ),
    .Y(_02210_));
 sky130_fd_sc_hd__buf_1 _31837_ (.A(_02210_),
    .X(_02211_));
 sky130_fd_sc_hd__buf_1 _31838_ (.A(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__a41oi_4 _31839_ (.A1(_02200_),
    .A2(_02206_),
    .A3(_02209_),
    .A4(_02212_),
    .B1(_02176_),
    .Y(_02213_));
 sky130_fd_sc_hd__a21o_4 _31840_ (.A1(\cpuregs[19][29] ),
    .A2(_02192_),
    .B1(_02213_),
    .X(_01078_));
 sky130_fd_sc_hd__buf_1 _31841_ (.A(_23681_),
    .X(_02214_));
 sky130_fd_sc_hd__and4_4 _31842_ (.A(_02165_),
    .B(_21829_),
    .C(_02194_),
    .D(_21863_),
    .X(_02215_));
 sky130_fd_sc_hd__a41oi_4 _31843_ (.A1(_21850_),
    .A2(_02180_),
    .A3(_21863_),
    .A4(_21886_),
    .B1(_01809_),
    .Y(_02216_));
 sky130_fd_sc_hd__o21ai_4 _31844_ (.A1(_21886_),
    .A2(_02215_),
    .B1(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__buf_1 _31845_ (.A(_02217_),
    .X(_02218_));
 sky130_fd_sc_hd__buf_1 _31846_ (.A(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__nand2_4 _31847_ (.A(_22872_),
    .B(_01825_),
    .Y(_02220_));
 sky130_fd_sc_hd__buf_1 _31848_ (.A(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__buf_1 _31849_ (.A(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__nand2_4 _31850_ (.A(_02110_),
    .B(\reg_next_pc[30] ),
    .Y(_02223_));
 sky130_fd_sc_hd__buf_1 _31851_ (.A(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__buf_1 _31852_ (.A(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__a41oi_4 _31853_ (.A1(_02214_),
    .A2(_02219_),
    .A3(_02222_),
    .A4(_02225_),
    .B1(_02176_),
    .Y(_02226_));
 sky130_fd_sc_hd__a21o_4 _31854_ (.A1(\cpuregs[19][30] ),
    .A2(_02192_),
    .B1(_02226_),
    .X(_01080_));
 sky130_fd_sc_hd__buf_1 _31855_ (.A(_23686_),
    .X(_02227_));
 sky130_fd_sc_hd__and4_4 _31856_ (.A(_02180_),
    .B(_21849_),
    .C(\reg_pc[29] ),
    .D(\reg_pc[30] ),
    .X(_02228_));
 sky130_fd_sc_hd__o21a_4 _31857_ (.A1(\reg_pc[31] ),
    .A2(_02228_),
    .B1(_01847_),
    .X(_02229_));
 sky130_fd_sc_hd__nand4_4 _31858_ (.A(_21864_),
    .B(_02202_),
    .C(_21886_),
    .D(_21900_),
    .Y(_02230_));
 sky130_fd_sc_hd__nand2_4 _31859_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__buf_1 _31860_ (.A(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__buf_1 _31861_ (.A(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__nand2_4 _31862_ (.A(_22902_),
    .B(_01825_),
    .Y(_02234_));
 sky130_fd_sc_hd__buf_1 _31863_ (.A(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__buf_1 _31864_ (.A(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__nand2_4 _31865_ (.A(_01800_),
    .B(\reg_next_pc[31] ),
    .Y(_02237_));
 sky130_fd_sc_hd__buf_1 _31866_ (.A(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__buf_1 _31867_ (.A(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__a41oi_4 _31868_ (.A1(_02227_),
    .A2(_02233_),
    .A3(_02236_),
    .A4(_02239_),
    .B1(_01771_),
    .Y(_02240_));
 sky130_fd_sc_hd__a21o_4 _31869_ (.A1(\cpuregs[19][31] ),
    .A2(_02192_),
    .B1(_02240_),
    .X(_01081_));
 sky130_fd_sc_hd__buf_1 _31870_ (.A(_01762_),
    .X(_02241_));
 sky130_fd_sc_hd__nor2_4 _31871_ (.A(\latched_rd[0] ),
    .B(_19085_),
    .Y(_02242_));
 sky130_fd_sc_hd__and4_4 _31872_ (.A(_02241_),
    .B(_01759_),
    .C(_01766_),
    .D(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__buf_1 _31873_ (.A(_02243_),
    .X(_02244_));
 sky130_vsdinv _31874_ (.A(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__buf_1 _31875_ (.A(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__buf_1 _31876_ (.A(_02246_),
    .X(_02247_));
 sky130_fd_sc_hd__buf_1 _31877_ (.A(_01782_),
    .X(_02248_));
 sky130_fd_sc_hd__buf_1 _31878_ (.A(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__nor2_4 _31879_ (.A(_02249_),
    .B(_02247_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21o_4 _31880_ (.A1(\cpuregs[18][0] ),
    .A2(_02247_),
    .B1(_02250_),
    .X(_01025_));
 sky130_fd_sc_hd__buf_1 _31881_ (.A(_02244_),
    .X(_02251_));
 sky130_fd_sc_hd__buf_1 _31882_ (.A(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__buf_1 _31883_ (.A(_01802_),
    .X(_02253_));
 sky130_fd_sc_hd__buf_1 _31884_ (.A(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__buf_1 _31885_ (.A(_02244_),
    .X(_02255_));
 sky130_fd_sc_hd__buf_1 _31886_ (.A(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__nand2_4 _31887_ (.A(_02254_),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__o21ai_4 _31888_ (.A1(_19392_),
    .A2(_02252_),
    .B1(_02257_),
    .Y(_01036_));
 sky130_fd_sc_hd__buf_1 _31889_ (.A(_01811_),
    .X(_02258_));
 sky130_fd_sc_hd__buf_1 _31890_ (.A(_01814_),
    .X(_02259_));
 sky130_fd_sc_hd__buf_1 _31891_ (.A(_01815_),
    .X(_02260_));
 sky130_fd_sc_hd__a41o_4 _31892_ (.A1(_02258_),
    .A2(_23473_),
    .A3(_02259_),
    .A4(_02260_),
    .B1(_02247_),
    .X(_02261_));
 sky130_fd_sc_hd__o21ai_4 _31893_ (.A1(_19486_),
    .A2(_02252_),
    .B1(_02261_),
    .Y(_01047_));
 sky130_fd_sc_hd__buf_1 _31894_ (.A(_01823_),
    .X(_02262_));
 sky130_fd_sc_hd__buf_1 _31895_ (.A(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__buf_1 _31896_ (.A(_01826_),
    .X(_02264_));
 sky130_fd_sc_hd__buf_1 _31897_ (.A(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__buf_1 _31898_ (.A(_01827_),
    .X(_02266_));
 sky130_fd_sc_hd__buf_1 _31899_ (.A(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__a41o_4 _31900_ (.A1(_23478_),
    .A2(_02263_),
    .A3(_02265_),
    .A4(_02267_),
    .B1(_02247_),
    .X(_02268_));
 sky130_fd_sc_hd__o21ai_4 _31901_ (.A1(_19559_),
    .A2(_02252_),
    .B1(_02268_),
    .Y(_01050_));
 sky130_fd_sc_hd__buf_1 _31902_ (.A(_01836_),
    .X(_02269_));
 sky130_fd_sc_hd__buf_1 _31903_ (.A(_01839_),
    .X(_02270_));
 sky130_fd_sc_hd__buf_1 _31904_ (.A(_01842_),
    .X(_02271_));
 sky130_fd_sc_hd__buf_1 _31905_ (.A(_02246_),
    .X(_02272_));
 sky130_fd_sc_hd__a41o_4 _31906_ (.A1(_02269_),
    .A2(_23488_),
    .A3(_02270_),
    .A4(_02271_),
    .B1(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__o21ai_4 _31907_ (.A1(_19635_),
    .A2(_02252_),
    .B1(_02273_),
    .Y(_01051_));
 sky130_fd_sc_hd__buf_1 _31908_ (.A(_02244_),
    .X(_02274_));
 sky130_fd_sc_hd__buf_1 _31909_ (.A(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__buf_1 _31910_ (.A(_01849_),
    .X(_02276_));
 sky130_fd_sc_hd__buf_1 _31911_ (.A(_01852_),
    .X(_02277_));
 sky130_fd_sc_hd__buf_1 _31912_ (.A(_01856_),
    .X(_02278_));
 sky130_fd_sc_hd__a41o_4 _31913_ (.A1(_02276_),
    .A2(_23495_),
    .A3(_02277_),
    .A4(_02278_),
    .B1(_02272_),
    .X(_02279_));
 sky130_fd_sc_hd__o21ai_4 _31914_ (.A1(_19687_),
    .A2(_02275_),
    .B1(_02279_),
    .Y(_01052_));
 sky130_fd_sc_hd__buf_1 _31915_ (.A(_01864_),
    .X(_02280_));
 sky130_fd_sc_hd__buf_1 _31916_ (.A(_01867_),
    .X(_02281_));
 sky130_fd_sc_hd__buf_1 _31917_ (.A(_01870_),
    .X(_02282_));
 sky130_fd_sc_hd__a41o_4 _31918_ (.A1(_02280_),
    .A2(_23505_),
    .A3(_02281_),
    .A4(_02282_),
    .B1(_02272_),
    .X(_02283_));
 sky130_fd_sc_hd__o21ai_4 _31919_ (.A1(_19742_),
    .A2(_02275_),
    .B1(_02283_),
    .Y(_01053_));
 sky130_fd_sc_hd__buf_1 _31920_ (.A(_01880_),
    .X(_02284_));
 sky130_fd_sc_hd__buf_1 _31921_ (.A(_01884_),
    .X(_02285_));
 sky130_fd_sc_hd__buf_1 _31922_ (.A(_01887_),
    .X(_02286_));
 sky130_fd_sc_hd__a41o_4 _31923_ (.A1(_02284_),
    .A2(_23511_),
    .A3(_02285_),
    .A4(_02286_),
    .B1(_02272_),
    .X(_02287_));
 sky130_fd_sc_hd__o21ai_4 _31924_ (.A1(_19789_),
    .A2(_02275_),
    .B1(_02287_),
    .Y(_01054_));
 sky130_fd_sc_hd__buf_1 _31925_ (.A(_01894_),
    .X(_02288_));
 sky130_fd_sc_hd__buf_1 _31926_ (.A(_01897_),
    .X(_02289_));
 sky130_fd_sc_hd__buf_1 _31927_ (.A(_01900_),
    .X(_02290_));
 sky130_fd_sc_hd__buf_1 _31928_ (.A(_02246_),
    .X(_02291_));
 sky130_fd_sc_hd__a41o_4 _31929_ (.A1(_02288_),
    .A2(_23520_),
    .A3(_02289_),
    .A4(_02290_),
    .B1(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__o21ai_4 _31930_ (.A1(_19855_),
    .A2(_02275_),
    .B1(_02292_),
    .Y(_01055_));
 sky130_fd_sc_hd__buf_1 _31931_ (.A(_02274_),
    .X(_02293_));
 sky130_fd_sc_hd__buf_1 _31932_ (.A(_01907_),
    .X(_02294_));
 sky130_fd_sc_hd__buf_1 _31933_ (.A(_01910_),
    .X(_02295_));
 sky130_fd_sc_hd__buf_1 _31934_ (.A(_01915_),
    .X(_02296_));
 sky130_fd_sc_hd__a41o_4 _31935_ (.A1(_02294_),
    .A2(_23527_),
    .A3(_02295_),
    .A4(_02296_),
    .B1(_02291_),
    .X(_02297_));
 sky130_fd_sc_hd__o21ai_4 _31936_ (.A1(_19909_),
    .A2(_02293_),
    .B1(_02297_),
    .Y(_01056_));
 sky130_fd_sc_hd__buf_1 _31937_ (.A(_01922_),
    .X(_02298_));
 sky130_fd_sc_hd__buf_1 _31938_ (.A(_01925_),
    .X(_02299_));
 sky130_fd_sc_hd__buf_1 _31939_ (.A(_01928_),
    .X(_02300_));
 sky130_fd_sc_hd__a41o_4 _31940_ (.A1(_02298_),
    .A2(_23537_),
    .A3(_02299_),
    .A4(_02300_),
    .B1(_02291_),
    .X(_02301_));
 sky130_fd_sc_hd__o21ai_4 _31941_ (.A1(_19966_),
    .A2(_02293_),
    .B1(_02301_),
    .Y(_01026_));
 sky130_fd_sc_hd__buf_1 _31942_ (.A(_01937_),
    .X(_02302_));
 sky130_fd_sc_hd__buf_1 _31943_ (.A(_01941_),
    .X(_02303_));
 sky130_fd_sc_hd__buf_1 _31944_ (.A(_01944_),
    .X(_02304_));
 sky130_fd_sc_hd__a41o_4 _31945_ (.A1(_02302_),
    .A2(_23543_),
    .A3(_02303_),
    .A4(_02304_),
    .B1(_02291_),
    .X(_02305_));
 sky130_fd_sc_hd__o21ai_4 _31946_ (.A1(_20037_),
    .A2(_02293_),
    .B1(_02305_),
    .Y(_01027_));
 sky130_fd_sc_hd__buf_1 _31947_ (.A(_01952_),
    .X(_02306_));
 sky130_fd_sc_hd__buf_1 _31948_ (.A(_01955_),
    .X(_02307_));
 sky130_fd_sc_hd__buf_1 _31949_ (.A(_01958_),
    .X(_02308_));
 sky130_fd_sc_hd__buf_1 _31950_ (.A(_02245_),
    .X(_02309_));
 sky130_fd_sc_hd__a41o_4 _31951_ (.A1(_02306_),
    .A2(_23551_),
    .A3(_02307_),
    .A4(_02308_),
    .B1(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__o21ai_4 _31952_ (.A1(_20104_),
    .A2(_02293_),
    .B1(_02310_),
    .Y(_01028_));
 sky130_fd_sc_hd__buf_1 _31953_ (.A(_02274_),
    .X(_02311_));
 sky130_fd_sc_hd__buf_1 _31954_ (.A(_01966_),
    .X(_02312_));
 sky130_fd_sc_hd__buf_1 _31955_ (.A(_01969_),
    .X(_02313_));
 sky130_fd_sc_hd__buf_1 _31956_ (.A(_01973_),
    .X(_02314_));
 sky130_fd_sc_hd__a41o_4 _31957_ (.A1(_02312_),
    .A2(_23558_),
    .A3(_02313_),
    .A4(_02314_),
    .B1(_02309_),
    .X(_02315_));
 sky130_fd_sc_hd__o21ai_4 _31958_ (.A1(_20159_),
    .A2(_02311_),
    .B1(_02315_),
    .Y(_01029_));
 sky130_fd_sc_hd__buf_1 _31959_ (.A(_01982_),
    .X(_02316_));
 sky130_fd_sc_hd__buf_1 _31960_ (.A(_01985_),
    .X(_02317_));
 sky130_fd_sc_hd__buf_1 _31961_ (.A(_01988_),
    .X(_02318_));
 sky130_fd_sc_hd__a41o_4 _31962_ (.A1(_02316_),
    .A2(_23568_),
    .A3(_02317_),
    .A4(_02318_),
    .B1(_02309_),
    .X(_02319_));
 sky130_fd_sc_hd__o21ai_4 _31963_ (.A1(_20219_),
    .A2(_02311_),
    .B1(_02319_),
    .Y(_01030_));
 sky130_fd_sc_hd__buf_1 _31964_ (.A(_01998_),
    .X(_02320_));
 sky130_fd_sc_hd__buf_1 _31965_ (.A(_02002_),
    .X(_02321_));
 sky130_fd_sc_hd__buf_1 _31966_ (.A(_02005_),
    .X(_02322_));
 sky130_fd_sc_hd__a41o_4 _31967_ (.A1(_02320_),
    .A2(_23574_),
    .A3(_02321_),
    .A4(_02322_),
    .B1(_02309_),
    .X(_02323_));
 sky130_fd_sc_hd__o21ai_4 _31968_ (.A1(_20268_),
    .A2(_02311_),
    .B1(_02323_),
    .Y(_01031_));
 sky130_fd_sc_hd__buf_1 _31969_ (.A(_02015_),
    .X(_02324_));
 sky130_fd_sc_hd__buf_1 _31970_ (.A(_02018_),
    .X(_02325_));
 sky130_fd_sc_hd__buf_1 _31971_ (.A(_02021_),
    .X(_02326_));
 sky130_fd_sc_hd__buf_1 _31972_ (.A(_02245_),
    .X(_02327_));
 sky130_fd_sc_hd__a41o_4 _31973_ (.A1(_02324_),
    .A2(_23583_),
    .A3(_02325_),
    .A4(_02326_),
    .B1(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__o21ai_4 _31974_ (.A1(_20319_),
    .A2(_02311_),
    .B1(_02328_),
    .Y(_01032_));
 sky130_fd_sc_hd__buf_1 _31975_ (.A(_02274_),
    .X(_02329_));
 sky130_fd_sc_hd__buf_1 _31976_ (.A(_02030_),
    .X(_02330_));
 sky130_fd_sc_hd__buf_1 _31977_ (.A(_02033_),
    .X(_02331_));
 sky130_fd_sc_hd__buf_1 _31978_ (.A(_02037_),
    .X(_02332_));
 sky130_fd_sc_hd__a41o_4 _31979_ (.A1(_02330_),
    .A2(_23591_),
    .A3(_02331_),
    .A4(_02332_),
    .B1(_02327_),
    .X(_02333_));
 sky130_fd_sc_hd__o21ai_4 _31980_ (.A1(_20366_),
    .A2(_02329_),
    .B1(_02333_),
    .Y(_01033_));
 sky130_fd_sc_hd__nand4_4 _31981_ (.A(_23598_),
    .B(_02043_),
    .C(_02047_),
    .D(_02050_),
    .Y(_02334_));
 sky130_fd_sc_hd__buf_1 _31982_ (.A(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__buf_1 _31983_ (.A(_02255_),
    .X(_02336_));
 sky130_fd_sc_hd__nand2_4 _31984_ (.A(_02335_),
    .B(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__o21ai_4 _31985_ (.A1(_20421_),
    .A2(_02329_),
    .B1(_02337_),
    .Y(_01034_));
 sky130_fd_sc_hd__buf_1 _31986_ (.A(_02060_),
    .X(_02338_));
 sky130_fd_sc_hd__buf_1 _31987_ (.A(_02063_),
    .X(_02339_));
 sky130_fd_sc_hd__buf_1 _31988_ (.A(_02066_),
    .X(_02340_));
 sky130_fd_sc_hd__a41o_4 _31989_ (.A1(_02338_),
    .A2(_23606_),
    .A3(_02339_),
    .A4(_02340_),
    .B1(_02327_),
    .X(_02341_));
 sky130_fd_sc_hd__o21ai_4 _31990_ (.A1(_20471_),
    .A2(_02329_),
    .B1(_02341_),
    .Y(_01035_));
 sky130_fd_sc_hd__buf_1 _31991_ (.A(_02076_),
    .X(_02342_));
 sky130_fd_sc_hd__buf_1 _31992_ (.A(_02080_),
    .X(_02343_));
 sky130_fd_sc_hd__buf_1 _31993_ (.A(_02083_),
    .X(_02344_));
 sky130_fd_sc_hd__a41o_4 _31994_ (.A1(_02342_),
    .A2(_23614_),
    .A3(_02343_),
    .A4(_02344_),
    .B1(_02327_),
    .X(_02345_));
 sky130_fd_sc_hd__o21ai_4 _31995_ (.A1(_20517_),
    .A2(_02329_),
    .B1(_02345_),
    .Y(_01037_));
 sky130_fd_sc_hd__buf_1 _31996_ (.A(_02255_),
    .X(_02346_));
 sky130_fd_sc_hd__buf_1 _31997_ (.A(_02091_),
    .X(_02347_));
 sky130_fd_sc_hd__buf_1 _31998_ (.A(_02094_),
    .X(_02348_));
 sky130_fd_sc_hd__buf_1 _31999_ (.A(_02097_),
    .X(_02349_));
 sky130_fd_sc_hd__buf_1 _32000_ (.A(_02245_),
    .X(_02350_));
 sky130_fd_sc_hd__a41o_4 _32001_ (.A1(_02347_),
    .A2(_23621_),
    .A3(_02348_),
    .A4(_02349_),
    .B1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__o21ai_4 _32002_ (.A1(_20566_),
    .A2(_02346_),
    .B1(_02351_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand4_4 _32003_ (.A(_23627_),
    .B(_02104_),
    .C(_02107_),
    .D(_02111_),
    .Y(_02352_));
 sky130_fd_sc_hd__buf_1 _32004_ (.A(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__nand2_4 _32005_ (.A(_02353_),
    .B(_02336_),
    .Y(_02354_));
 sky130_fd_sc_hd__o21ai_4 _32006_ (.A1(_20608_),
    .A2(_02346_),
    .B1(_02354_),
    .Y(_01039_));
 sky130_fd_sc_hd__buf_1 _32007_ (.A(_02121_),
    .X(_02355_));
 sky130_fd_sc_hd__buf_1 _32008_ (.A(_02124_),
    .X(_02356_));
 sky130_fd_sc_hd__buf_1 _32009_ (.A(_02128_),
    .X(_02357_));
 sky130_fd_sc_hd__a41o_4 _32010_ (.A1(_02355_),
    .A2(_23634_),
    .A3(_02356_),
    .A4(_02357_),
    .B1(_02350_),
    .X(_02358_));
 sky130_fd_sc_hd__o21ai_4 _32011_ (.A1(_20650_),
    .A2(_02346_),
    .B1(_02358_),
    .Y(_01040_));
 sky130_fd_sc_hd__buf_1 _32012_ (.A(_02138_),
    .X(_02359_));
 sky130_fd_sc_hd__buf_1 _32013_ (.A(_02141_),
    .X(_02360_));
 sky130_fd_sc_hd__buf_1 _32014_ (.A(_02144_),
    .X(_02361_));
 sky130_fd_sc_hd__a41o_4 _32015_ (.A1(_02359_),
    .A2(_23642_),
    .A3(_02360_),
    .A4(_02361_),
    .B1(_02350_),
    .X(_02362_));
 sky130_fd_sc_hd__o21ai_4 _32016_ (.A1(_20696_),
    .A2(_02346_),
    .B1(_02362_),
    .Y(_01041_));
 sky130_fd_sc_hd__buf_1 _32017_ (.A(_02255_),
    .X(_02363_));
 sky130_fd_sc_hd__buf_1 _32018_ (.A(_02153_),
    .X(_02364_));
 sky130_fd_sc_hd__buf_1 _32019_ (.A(_02156_),
    .X(_02365_));
 sky130_fd_sc_hd__buf_1 _32020_ (.A(_02159_),
    .X(_02366_));
 sky130_fd_sc_hd__a41o_4 _32021_ (.A1(_02364_),
    .A2(_23649_),
    .A3(_02365_),
    .A4(_02366_),
    .B1(_02350_),
    .X(_02367_));
 sky130_fd_sc_hd__o21ai_4 _32022_ (.A1(_20743_),
    .A2(_02363_),
    .B1(_02367_),
    .Y(_01042_));
 sky130_fd_sc_hd__buf_1 _32023_ (.A(_02167_),
    .X(_02368_));
 sky130_fd_sc_hd__buf_1 _32024_ (.A(_02170_),
    .X(_02369_));
 sky130_fd_sc_hd__buf_1 _32025_ (.A(_02173_),
    .X(_02370_));
 sky130_fd_sc_hd__a41o_4 _32026_ (.A1(_02368_),
    .A2(_23657_),
    .A3(_02369_),
    .A4(_02370_),
    .B1(_02246_),
    .X(_02371_));
 sky130_fd_sc_hd__o21ai_4 _32027_ (.A1(_20786_),
    .A2(_02363_),
    .B1(_02371_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand4_4 _32028_ (.A(_23661_),
    .B(_02182_),
    .C(_02185_),
    .D(_02188_),
    .Y(_02372_));
 sky130_fd_sc_hd__buf_1 _32029_ (.A(_02372_),
    .X(_02373_));
 sky130_fd_sc_hd__nand2_4 _32030_ (.A(_02373_),
    .B(_02336_),
    .Y(_02374_));
 sky130_fd_sc_hd__o21ai_4 _32031_ (.A1(_20834_),
    .A2(_02363_),
    .B1(_02374_),
    .Y(_01044_));
 sky130_fd_sc_hd__buf_1 _32032_ (.A(_02197_),
    .X(_02375_));
 sky130_fd_sc_hd__buf_1 _32033_ (.A(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__nand2_4 _32034_ (.A(_02376_),
    .B(_02336_),
    .Y(_02377_));
 sky130_fd_sc_hd__o21ai_4 _32035_ (.A1(_20876_),
    .A2(_02363_),
    .B1(_02377_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand4_4 _32036_ (.A(_23673_),
    .B(_02204_),
    .C(_02207_),
    .D(_02210_),
    .Y(_02378_));
 sky130_fd_sc_hd__buf_1 _32037_ (.A(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__nand2_4 _32038_ (.A(_02379_),
    .B(_02251_),
    .Y(_02380_));
 sky130_fd_sc_hd__o21ai_4 _32039_ (.A1(_20923_),
    .A2(_02256_),
    .B1(_02380_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand4_4 _32040_ (.A(_23680_),
    .B(_02217_),
    .C(_02220_),
    .D(_02223_),
    .Y(_02381_));
 sky130_fd_sc_hd__buf_1 _32041_ (.A(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__nand2_4 _32042_ (.A(_02382_),
    .B(_02251_),
    .Y(_02383_));
 sky130_fd_sc_hd__o21ai_4 _32043_ (.A1(_20963_),
    .A2(_02256_),
    .B1(_02383_),
    .Y(_01048_));
 sky130_fd_sc_hd__nand4_4 _32044_ (.A(_23685_),
    .B(_02231_),
    .C(_02234_),
    .D(_02237_),
    .Y(_02384_));
 sky130_fd_sc_hd__buf_1 _32045_ (.A(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__nand2_4 _32046_ (.A(_02385_),
    .B(_02251_),
    .Y(_02386_));
 sky130_fd_sc_hd__o21ai_4 _32047_ (.A1(_21006_),
    .A2(_02256_),
    .B1(_02386_),
    .Y(_01049_));
 sky130_fd_sc_hd__nor4_4 _32048_ (.A(_19069_),
    .B(_01787_),
    .C(_01760_),
    .D(_01768_),
    .Y(_02387_));
 sky130_vsdinv _32049_ (.A(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__buf_1 _32050_ (.A(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__buf_1 _32051_ (.A(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__buf_1 _32052_ (.A(_01782_),
    .X(_02391_));
 sky130_fd_sc_hd__and4_4 _32053_ (.A(_01784_),
    .B(_01785_),
    .C(_19087_),
    .D(_01788_),
    .X(_02392_));
 sky130_vsdinv _32054_ (.A(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__nor3_4 _32055_ (.A(_01773_),
    .B(_02391_),
    .C(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__a21o_4 _32056_ (.A1(\cpuregs[17][0] ),
    .A2(_02390_),
    .B1(_02394_),
    .X(_00993_));
 sky130_fd_sc_hd__buf_1 _32057_ (.A(_01802_),
    .X(_02395_));
 sky130_fd_sc_hd__and2_4 _32058_ (.A(_02387_),
    .B(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__a21o_4 _32059_ (.A1(\cpuregs[17][1] ),
    .A2(_02390_),
    .B1(_02396_),
    .X(_01004_));
 sky130_fd_sc_hd__buf_1 _32060_ (.A(_02388_),
    .X(_02397_));
 sky130_fd_sc_hd__buf_1 _32061_ (.A(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__nor2_4 _32062_ (.A(_02398_),
    .B(_01817_),
    .Y(_02399_));
 sky130_fd_sc_hd__a21o_4 _32063_ (.A1(\cpuregs[17][2] ),
    .A2(_02390_),
    .B1(_02399_),
    .X(_01015_));
 sky130_fd_sc_hd__nor2_4 _32064_ (.A(_02398_),
    .B(_01829_),
    .Y(_02400_));
 sky130_fd_sc_hd__a21o_4 _32065_ (.A1(\cpuregs[17][3] ),
    .A2(_02390_),
    .B1(_02400_),
    .X(_01018_));
 sky130_fd_sc_hd__buf_1 _32066_ (.A(_02389_),
    .X(_02401_));
 sky130_fd_sc_hd__a41oi_4 _32067_ (.A1(_01832_),
    .A2(_01838_),
    .A3(_01841_),
    .A4(_01844_),
    .B1(_02398_),
    .Y(_02402_));
 sky130_fd_sc_hd__a21o_4 _32068_ (.A1(\cpuregs[17][4] ),
    .A2(_02401_),
    .B1(_02402_),
    .X(_01019_));
 sky130_fd_sc_hd__a41oi_4 _32069_ (.A1(_01846_),
    .A2(_01851_),
    .A3(_01854_),
    .A4(_01858_),
    .B1(_02398_),
    .Y(_02403_));
 sky130_fd_sc_hd__a21o_4 _32070_ (.A1(\cpuregs[17][5] ),
    .A2(_02401_),
    .B1(_02403_),
    .X(_01020_));
 sky130_fd_sc_hd__buf_1 _32071_ (.A(_02388_),
    .X(_02404_));
 sky130_fd_sc_hd__buf_1 _32072_ (.A(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__a41oi_4 _32073_ (.A1(_01860_),
    .A2(_01866_),
    .A3(_01869_),
    .A4(_01872_),
    .B1(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__a21o_4 _32074_ (.A1(\cpuregs[17][6] ),
    .A2(_02401_),
    .B1(_02406_),
    .X(_01021_));
 sky130_fd_sc_hd__a41oi_4 _32075_ (.A1(_01876_),
    .A2(_01882_),
    .A3(_01886_),
    .A4(_01889_),
    .B1(_02405_),
    .Y(_02407_));
 sky130_fd_sc_hd__a21o_4 _32076_ (.A1(\cpuregs[17][7] ),
    .A2(_02401_),
    .B1(_02407_),
    .X(_01022_));
 sky130_fd_sc_hd__buf_1 _32077_ (.A(_02389_),
    .X(_02408_));
 sky130_fd_sc_hd__a41oi_4 _32078_ (.A1(_01892_),
    .A2(_01896_),
    .A3(_01899_),
    .A4(_01902_),
    .B1(_02405_),
    .Y(_02409_));
 sky130_fd_sc_hd__a21o_4 _32079_ (.A1(\cpuregs[17][8] ),
    .A2(_02408_),
    .B1(_02409_),
    .X(_01023_));
 sky130_fd_sc_hd__a41oi_4 _32080_ (.A1(_01904_),
    .A2(_01909_),
    .A3(_01912_),
    .A4(_01917_),
    .B1(_02405_),
    .Y(_02410_));
 sky130_fd_sc_hd__a21o_4 _32081_ (.A1(\cpuregs[17][9] ),
    .A2(_02408_),
    .B1(_02410_),
    .X(_01024_));
 sky130_fd_sc_hd__buf_1 _32082_ (.A(_02404_),
    .X(_02411_));
 sky130_fd_sc_hd__a41oi_4 _32083_ (.A1(_01919_),
    .A2(_01924_),
    .A3(_01927_),
    .A4(_01930_),
    .B1(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__a21o_4 _32084_ (.A1(\cpuregs[17][10] ),
    .A2(_02408_),
    .B1(_02412_),
    .X(_00994_));
 sky130_fd_sc_hd__a41oi_4 _32085_ (.A1(_01933_),
    .A2(_01939_),
    .A3(_01943_),
    .A4(_01946_),
    .B1(_02411_),
    .Y(_02413_));
 sky130_fd_sc_hd__a21o_4 _32086_ (.A1(\cpuregs[17][11] ),
    .A2(_02408_),
    .B1(_02413_),
    .X(_00995_));
 sky130_fd_sc_hd__buf_1 _32087_ (.A(_02388_),
    .X(_02414_));
 sky130_fd_sc_hd__buf_1 _32088_ (.A(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__a41oi_4 _32089_ (.A1(_01950_),
    .A2(_01954_),
    .A3(_01957_),
    .A4(_01960_),
    .B1(_02411_),
    .Y(_02416_));
 sky130_fd_sc_hd__a21o_4 _32090_ (.A1(\cpuregs[17][12] ),
    .A2(_02415_),
    .B1(_02416_),
    .X(_00996_));
 sky130_fd_sc_hd__a41oi_4 _32091_ (.A1(_01962_),
    .A2(_01968_),
    .A3(_01971_),
    .A4(_01975_),
    .B1(_02411_),
    .Y(_02417_));
 sky130_fd_sc_hd__a21o_4 _32092_ (.A1(\cpuregs[17][13] ),
    .A2(_02415_),
    .B1(_02417_),
    .X(_00997_));
 sky130_fd_sc_hd__buf_1 _32093_ (.A(_02404_),
    .X(_02418_));
 sky130_fd_sc_hd__a41oi_4 _32094_ (.A1(_01977_),
    .A2(_01984_),
    .A3(_01987_),
    .A4(_01990_),
    .B1(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21o_4 _32095_ (.A1(\cpuregs[17][14] ),
    .A2(_02415_),
    .B1(_02419_),
    .X(_00998_));
 sky130_fd_sc_hd__a41oi_4 _32096_ (.A1(_01993_),
    .A2(_02000_),
    .A3(_02004_),
    .A4(_02007_),
    .B1(_02418_),
    .Y(_02420_));
 sky130_fd_sc_hd__a21o_4 _32097_ (.A1(\cpuregs[17][15] ),
    .A2(_02415_),
    .B1(_02420_),
    .X(_00999_));
 sky130_fd_sc_hd__buf_1 _32098_ (.A(_02414_),
    .X(_02421_));
 sky130_fd_sc_hd__a41oi_4 _32099_ (.A1(_02010_),
    .A2(_02017_),
    .A3(_02020_),
    .A4(_02023_),
    .B1(_02418_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21o_4 _32100_ (.A1(\cpuregs[17][16] ),
    .A2(_02421_),
    .B1(_02422_),
    .X(_01000_));
 sky130_fd_sc_hd__a41oi_4 _32101_ (.A1(_02025_),
    .A2(_02032_),
    .A3(_02035_),
    .A4(_02039_),
    .B1(_02418_),
    .Y(_02423_));
 sky130_fd_sc_hd__a21o_4 _32102_ (.A1(\cpuregs[17][17] ),
    .A2(_02421_),
    .B1(_02423_),
    .X(_01001_));
 sky130_fd_sc_hd__buf_1 _32103_ (.A(_02397_),
    .X(_02424_));
 sky130_fd_sc_hd__a41oi_4 _32104_ (.A1(_02041_),
    .A2(_02045_),
    .A3(_02049_),
    .A4(_02052_),
    .B1(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__a21o_4 _32105_ (.A1(\cpuregs[17][18] ),
    .A2(_02421_),
    .B1(_02425_),
    .X(_01002_));
 sky130_fd_sc_hd__a41oi_4 _32106_ (.A1(_02055_),
    .A2(_02062_),
    .A3(_02065_),
    .A4(_02068_),
    .B1(_02424_),
    .Y(_02426_));
 sky130_fd_sc_hd__a21o_4 _32107_ (.A1(\cpuregs[17][19] ),
    .A2(_02421_),
    .B1(_02426_),
    .X(_01003_));
 sky130_fd_sc_hd__buf_1 _32108_ (.A(_02414_),
    .X(_02427_));
 sky130_fd_sc_hd__a41oi_4 _32109_ (.A1(_02071_),
    .A2(_02078_),
    .A3(_02082_),
    .A4(_02085_),
    .B1(_02424_),
    .Y(_02428_));
 sky130_fd_sc_hd__a21o_4 _32110_ (.A1(\cpuregs[17][20] ),
    .A2(_02427_),
    .B1(_02428_),
    .X(_01005_));
 sky130_fd_sc_hd__a41oi_4 _32111_ (.A1(_02087_),
    .A2(_02093_),
    .A3(_02096_),
    .A4(_02099_),
    .B1(_02424_),
    .Y(_02429_));
 sky130_fd_sc_hd__a21o_4 _32112_ (.A1(\cpuregs[17][21] ),
    .A2(_02427_),
    .B1(_02429_),
    .X(_01006_));
 sky130_fd_sc_hd__buf_1 _32113_ (.A(_02397_),
    .X(_02430_));
 sky130_fd_sc_hd__a41oi_4 _32114_ (.A1(_02101_),
    .A2(_02106_),
    .A3(_02109_),
    .A4(_02113_),
    .B1(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__a21o_4 _32115_ (.A1(\cpuregs[17][22] ),
    .A2(_02427_),
    .B1(_02431_),
    .X(_01007_));
 sky130_fd_sc_hd__a41oi_4 _32116_ (.A1(_02116_),
    .A2(_02123_),
    .A3(_02126_),
    .A4(_02130_),
    .B1(_02430_),
    .Y(_02432_));
 sky130_fd_sc_hd__a21o_4 _32117_ (.A1(\cpuregs[17][23] ),
    .A2(_02427_),
    .B1(_02432_),
    .X(_01008_));
 sky130_fd_sc_hd__buf_1 _32118_ (.A(_02414_),
    .X(_02433_));
 sky130_fd_sc_hd__a41oi_4 _32119_ (.A1(_02133_),
    .A2(_02140_),
    .A3(_02143_),
    .A4(_02146_),
    .B1(_02430_),
    .Y(_02434_));
 sky130_fd_sc_hd__a21o_4 _32120_ (.A1(\cpuregs[17][24] ),
    .A2(_02433_),
    .B1(_02434_),
    .X(_01009_));
 sky130_fd_sc_hd__a41oi_4 _32121_ (.A1(_02148_),
    .A2(_02155_),
    .A3(_02158_),
    .A4(_02161_),
    .B1(_02430_),
    .Y(_02435_));
 sky130_fd_sc_hd__a21o_4 _32122_ (.A1(\cpuregs[17][25] ),
    .A2(_02433_),
    .B1(_02435_),
    .X(_01010_));
 sky130_fd_sc_hd__buf_1 _32123_ (.A(_02397_),
    .X(_02436_));
 sky130_fd_sc_hd__a41oi_4 _32124_ (.A1(_02163_),
    .A2(_02169_),
    .A3(_02172_),
    .A4(_02175_),
    .B1(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__a21o_4 _32125_ (.A1(\cpuregs[17][26] ),
    .A2(_02433_),
    .B1(_02437_),
    .X(_01011_));
 sky130_fd_sc_hd__a41oi_4 _32126_ (.A1(_02178_),
    .A2(_02184_),
    .A3(_02187_),
    .A4(_02190_),
    .B1(_02436_),
    .Y(_02438_));
 sky130_fd_sc_hd__a21o_4 _32127_ (.A1(\cpuregs[17][27] ),
    .A2(_02433_),
    .B1(_02438_),
    .X(_01012_));
 sky130_fd_sc_hd__buf_1 _32128_ (.A(_02404_),
    .X(_02439_));
 sky130_fd_sc_hd__and2_4 _32129_ (.A(_02198_),
    .B(_02387_),
    .X(_02440_));
 sky130_fd_sc_hd__a21o_4 _32130_ (.A1(\cpuregs[17][28] ),
    .A2(_02439_),
    .B1(_02440_),
    .X(_01013_));
 sky130_fd_sc_hd__a41oi_4 _32131_ (.A1(_02200_),
    .A2(_02206_),
    .A3(_02209_),
    .A4(_02212_),
    .B1(_02436_),
    .Y(_02441_));
 sky130_fd_sc_hd__a21o_4 _32132_ (.A1(\cpuregs[17][29] ),
    .A2(_02439_),
    .B1(_02441_),
    .X(_01014_));
 sky130_fd_sc_hd__a41oi_4 _32133_ (.A1(_02214_),
    .A2(_02219_),
    .A3(_02222_),
    .A4(_02225_),
    .B1(_02436_),
    .Y(_02442_));
 sky130_fd_sc_hd__a21o_4 _32134_ (.A1(\cpuregs[17][30] ),
    .A2(_02439_),
    .B1(_02442_),
    .X(_01016_));
 sky130_fd_sc_hd__a41oi_4 _32135_ (.A1(_02227_),
    .A2(_02233_),
    .A3(_02236_),
    .A4(_02239_),
    .B1(_02389_),
    .Y(_02443_));
 sky130_fd_sc_hd__a21o_4 _32136_ (.A1(\cpuregs[17][31] ),
    .A2(_02439_),
    .B1(_02443_),
    .X(_01017_));
 sky130_fd_sc_hd__nand4_4 _32137_ (.A(_19067_),
    .B(_01763_),
    .C(_19085_),
    .D(_01766_),
    .Y(_02444_));
 sky130_fd_sc_hd__buf_1 _32138_ (.A(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__nor2_4 _32139_ (.A(_01773_),
    .B(_02445_),
    .Y(_02446_));
 sky130_vsdinv _32140_ (.A(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__buf_1 _32141_ (.A(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__buf_1 _32142_ (.A(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__buf_1 _32143_ (.A(_02445_),
    .X(_02450_));
 sky130_fd_sc_hd__buf_1 _32144_ (.A(_01782_),
    .X(_02451_));
 sky130_fd_sc_hd__nor3_4 _32145_ (.A(_01773_),
    .B(_02450_),
    .C(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__a21o_4 _32146_ (.A1(\cpuregs[16][0] ),
    .A2(_02449_),
    .B1(_02452_),
    .X(_00961_));
 sky130_fd_sc_hd__buf_1 _32147_ (.A(_02446_),
    .X(_02453_));
 sky130_fd_sc_hd__buf_1 _32148_ (.A(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__buf_1 _32149_ (.A(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__buf_1 _32150_ (.A(_02453_),
    .X(_02456_));
 sky130_fd_sc_hd__nand2_4 _32151_ (.A(_02254_),
    .B(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__o21ai_4 _32152_ (.A1(_19403_),
    .A2(_02455_),
    .B1(_02457_),
    .Y(_00972_));
 sky130_fd_sc_hd__buf_1 _32153_ (.A(_23472_),
    .X(_02458_));
 sky130_fd_sc_hd__buf_1 _32154_ (.A(_01811_),
    .X(_02459_));
 sky130_fd_sc_hd__buf_1 _32155_ (.A(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__buf_1 _32156_ (.A(_01814_),
    .X(_02461_));
 sky130_fd_sc_hd__buf_1 _32157_ (.A(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__buf_1 _32158_ (.A(_01815_),
    .X(_02463_));
 sky130_fd_sc_hd__buf_1 _32159_ (.A(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__buf_1 _32160_ (.A(_02448_),
    .X(_02465_));
 sky130_fd_sc_hd__a41oi_4 _32161_ (.A1(_02458_),
    .A2(_02460_),
    .A3(_02462_),
    .A4(_02464_),
    .B1(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__a21o_4 _32162_ (.A1(\cpuregs[16][2] ),
    .A2(_02449_),
    .B1(_02466_),
    .X(_00983_));
 sky130_fd_sc_hd__nor2_4 _32163_ (.A(_02449_),
    .B(_01829_),
    .Y(_02467_));
 sky130_fd_sc_hd__a21o_4 _32164_ (.A1(\cpuregs[16][3] ),
    .A2(_02449_),
    .B1(_02467_),
    .X(_00986_));
 sky130_fd_sc_hd__buf_1 _32165_ (.A(_23487_),
    .X(_02468_));
 sky130_fd_sc_hd__a41o_4 _32166_ (.A1(_02269_),
    .A2(_02468_),
    .A3(_02270_),
    .A4(_02271_),
    .B1(_02465_),
    .X(_02469_));
 sky130_fd_sc_hd__o21ai_4 _32167_ (.A1(_19642_),
    .A2(_02455_),
    .B1(_02469_),
    .Y(_00987_));
 sky130_fd_sc_hd__buf_1 _32168_ (.A(_23494_),
    .X(_02470_));
 sky130_fd_sc_hd__a41o_4 _32169_ (.A1(_02276_),
    .A2(_02470_),
    .A3(_02277_),
    .A4(_02278_),
    .B1(_02465_),
    .X(_02471_));
 sky130_fd_sc_hd__o21ai_4 _32170_ (.A1(_19690_),
    .A2(_02455_),
    .B1(_02471_),
    .Y(_00988_));
 sky130_fd_sc_hd__buf_1 _32171_ (.A(_23504_),
    .X(_02472_));
 sky130_fd_sc_hd__a41o_4 _32172_ (.A1(_02280_),
    .A2(_02472_),
    .A3(_02281_),
    .A4(_02282_),
    .B1(_02465_),
    .X(_02473_));
 sky130_fd_sc_hd__o21ai_4 _32173_ (.A1(_19746_),
    .A2(_02455_),
    .B1(_02473_),
    .Y(_00989_));
 sky130_fd_sc_hd__buf_1 _32174_ (.A(_02454_),
    .X(_02474_));
 sky130_fd_sc_hd__buf_1 _32175_ (.A(_23510_),
    .X(_02475_));
 sky130_fd_sc_hd__buf_1 _32176_ (.A(_02447_),
    .X(_02476_));
 sky130_fd_sc_hd__buf_1 _32177_ (.A(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__a41o_4 _32178_ (.A1(_02284_),
    .A2(_02475_),
    .A3(_02285_),
    .A4(_02286_),
    .B1(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__o21ai_4 _32179_ (.A1(_19793_),
    .A2(_02474_),
    .B1(_02478_),
    .Y(_00990_));
 sky130_fd_sc_hd__buf_1 _32180_ (.A(_23519_),
    .X(_02479_));
 sky130_fd_sc_hd__a41o_4 _32181_ (.A1(_02288_),
    .A2(_02479_),
    .A3(_02289_),
    .A4(_02290_),
    .B1(_02477_),
    .X(_02480_));
 sky130_fd_sc_hd__o21ai_4 _32182_ (.A1(_19859_),
    .A2(_02474_),
    .B1(_02480_),
    .Y(_00991_));
 sky130_fd_sc_hd__buf_1 _32183_ (.A(_23526_),
    .X(_02481_));
 sky130_fd_sc_hd__a41o_4 _32184_ (.A1(_02294_),
    .A2(_02481_),
    .A3(_02295_),
    .A4(_02296_),
    .B1(_02477_),
    .X(_02482_));
 sky130_fd_sc_hd__o21ai_4 _32185_ (.A1(_19914_),
    .A2(_02474_),
    .B1(_02482_),
    .Y(_00992_));
 sky130_fd_sc_hd__buf_1 _32186_ (.A(_23536_),
    .X(_02483_));
 sky130_fd_sc_hd__a41o_4 _32187_ (.A1(_02298_),
    .A2(_02483_),
    .A3(_02299_),
    .A4(_02300_),
    .B1(_02477_),
    .X(_02484_));
 sky130_fd_sc_hd__o21ai_4 _32188_ (.A1(_19970_),
    .A2(_02474_),
    .B1(_02484_),
    .Y(_00962_));
 sky130_fd_sc_hd__buf_1 _32189_ (.A(_02454_),
    .X(_02485_));
 sky130_fd_sc_hd__buf_1 _32190_ (.A(_23542_),
    .X(_02486_));
 sky130_fd_sc_hd__buf_1 _32191_ (.A(_02476_),
    .X(_02487_));
 sky130_fd_sc_hd__a41o_4 _32192_ (.A1(_02302_),
    .A2(_02486_),
    .A3(_02303_),
    .A4(_02304_),
    .B1(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__o21ai_4 _32193_ (.A1(_20043_),
    .A2(_02485_),
    .B1(_02488_),
    .Y(_00963_));
 sky130_fd_sc_hd__buf_1 _32194_ (.A(_23550_),
    .X(_02489_));
 sky130_fd_sc_hd__a41o_4 _32195_ (.A1(_02306_),
    .A2(_02489_),
    .A3(_02307_),
    .A4(_02308_),
    .B1(_02487_),
    .X(_02490_));
 sky130_fd_sc_hd__o21ai_4 _32196_ (.A1(_20107_),
    .A2(_02485_),
    .B1(_02490_),
    .Y(_00964_));
 sky130_fd_sc_hd__buf_1 _32197_ (.A(_23557_),
    .X(_02491_));
 sky130_fd_sc_hd__a41o_4 _32198_ (.A1(_02312_),
    .A2(_02491_),
    .A3(_02313_),
    .A4(_02314_),
    .B1(_02487_),
    .X(_02492_));
 sky130_fd_sc_hd__o21ai_4 _32199_ (.A1(_20164_),
    .A2(_02485_),
    .B1(_02492_),
    .Y(_00965_));
 sky130_fd_sc_hd__buf_1 _32200_ (.A(_23567_),
    .X(_02493_));
 sky130_fd_sc_hd__a41o_4 _32201_ (.A1(_02316_),
    .A2(_02493_),
    .A3(_02317_),
    .A4(_02318_),
    .B1(_02487_),
    .X(_02494_));
 sky130_fd_sc_hd__o21ai_4 _32202_ (.A1(_20222_),
    .A2(_02485_),
    .B1(_02494_),
    .Y(_00966_));
 sky130_fd_sc_hd__buf_1 _32203_ (.A(_02453_),
    .X(_02495_));
 sky130_fd_sc_hd__buf_1 _32204_ (.A(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__buf_1 _32205_ (.A(_23573_),
    .X(_02497_));
 sky130_fd_sc_hd__buf_1 _32206_ (.A(_02476_),
    .X(_02498_));
 sky130_fd_sc_hd__a41o_4 _32207_ (.A1(_02320_),
    .A2(_02497_),
    .A3(_02321_),
    .A4(_02322_),
    .B1(_02498_),
    .X(_02499_));
 sky130_fd_sc_hd__o21ai_4 _32208_ (.A1(_20271_),
    .A2(_02496_),
    .B1(_02499_),
    .Y(_00967_));
 sky130_fd_sc_hd__buf_1 _32209_ (.A(_23582_),
    .X(_02500_));
 sky130_fd_sc_hd__a41o_4 _32210_ (.A1(_02324_),
    .A2(_02500_),
    .A3(_02325_),
    .A4(_02326_),
    .B1(_02498_),
    .X(_02501_));
 sky130_fd_sc_hd__o21ai_4 _32211_ (.A1(_20322_),
    .A2(_02496_),
    .B1(_02501_),
    .Y(_00968_));
 sky130_fd_sc_hd__buf_1 _32212_ (.A(_23590_),
    .X(_02502_));
 sky130_fd_sc_hd__a41o_4 _32213_ (.A1(_02330_),
    .A2(_02502_),
    .A3(_02331_),
    .A4(_02332_),
    .B1(_02498_),
    .X(_02503_));
 sky130_fd_sc_hd__o21ai_4 _32214_ (.A1(_20370_),
    .A2(_02496_),
    .B1(_02503_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_4 _32215_ (.A(_02335_),
    .B(_02456_),
    .Y(_02504_));
 sky130_fd_sc_hd__o21ai_4 _32216_ (.A1(_20424_),
    .A2(_02496_),
    .B1(_02504_),
    .Y(_00970_));
 sky130_fd_sc_hd__buf_1 _32217_ (.A(_02495_),
    .X(_02505_));
 sky130_fd_sc_hd__buf_1 _32218_ (.A(_23605_),
    .X(_02506_));
 sky130_fd_sc_hd__a41o_4 _32219_ (.A1(_02338_),
    .A2(_02506_),
    .A3(_02339_),
    .A4(_02340_),
    .B1(_02498_),
    .X(_02507_));
 sky130_fd_sc_hd__o21ai_4 _32220_ (.A1(_20474_),
    .A2(_02505_),
    .B1(_02507_),
    .Y(_00971_));
 sky130_fd_sc_hd__buf_1 _32221_ (.A(_23613_),
    .X(_02508_));
 sky130_fd_sc_hd__buf_1 _32222_ (.A(_02476_),
    .X(_02509_));
 sky130_fd_sc_hd__a41o_4 _32223_ (.A1(_02342_),
    .A2(_02508_),
    .A3(_02343_),
    .A4(_02344_),
    .B1(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__o21ai_4 _32224_ (.A1(_20521_),
    .A2(_02505_),
    .B1(_02510_),
    .Y(_00973_));
 sky130_fd_sc_hd__buf_1 _32225_ (.A(_23620_),
    .X(_02511_));
 sky130_fd_sc_hd__a41o_4 _32226_ (.A1(_02347_),
    .A2(_02511_),
    .A3(_02348_),
    .A4(_02349_),
    .B1(_02509_),
    .X(_02512_));
 sky130_fd_sc_hd__o21ai_4 _32227_ (.A1(_20569_),
    .A2(_02505_),
    .B1(_02512_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand2_4 _32228_ (.A(_02353_),
    .B(_02456_),
    .Y(_02513_));
 sky130_fd_sc_hd__o21ai_4 _32229_ (.A1(_20612_),
    .A2(_02505_),
    .B1(_02513_),
    .Y(_00975_));
 sky130_fd_sc_hd__buf_1 _32230_ (.A(_02495_),
    .X(_02514_));
 sky130_fd_sc_hd__buf_1 _32231_ (.A(_23633_),
    .X(_02515_));
 sky130_fd_sc_hd__a41o_4 _32232_ (.A1(_02355_),
    .A2(_02515_),
    .A3(_02356_),
    .A4(_02357_),
    .B1(_02509_),
    .X(_02516_));
 sky130_fd_sc_hd__o21ai_4 _32233_ (.A1(_20653_),
    .A2(_02514_),
    .B1(_02516_),
    .Y(_00976_));
 sky130_fd_sc_hd__buf_1 _32234_ (.A(_23641_),
    .X(_02517_));
 sky130_fd_sc_hd__a41o_4 _32235_ (.A1(_02359_),
    .A2(_02517_),
    .A3(_02360_),
    .A4(_02361_),
    .B1(_02509_),
    .X(_02518_));
 sky130_fd_sc_hd__o21ai_4 _32236_ (.A1(_20699_),
    .A2(_02514_),
    .B1(_02518_),
    .Y(_00977_));
 sky130_fd_sc_hd__buf_1 _32237_ (.A(_23648_),
    .X(_02519_));
 sky130_fd_sc_hd__a41o_4 _32238_ (.A1(_02364_),
    .A2(_02519_),
    .A3(_02365_),
    .A4(_02366_),
    .B1(_02448_),
    .X(_02520_));
 sky130_fd_sc_hd__o21ai_4 _32239_ (.A1(_20746_),
    .A2(_02514_),
    .B1(_02520_),
    .Y(_00978_));
 sky130_fd_sc_hd__buf_1 _32240_ (.A(_23656_),
    .X(_02521_));
 sky130_fd_sc_hd__a41o_4 _32241_ (.A1(_02368_),
    .A2(_02521_),
    .A3(_02369_),
    .A4(_02370_),
    .B1(_02448_),
    .X(_02522_));
 sky130_fd_sc_hd__o21ai_4 _32242_ (.A1(_20789_),
    .A2(_02514_),
    .B1(_02522_),
    .Y(_00979_));
 sky130_fd_sc_hd__buf_1 _32243_ (.A(_02495_),
    .X(_02523_));
 sky130_fd_sc_hd__buf_1 _32244_ (.A(_02453_),
    .X(_02524_));
 sky130_fd_sc_hd__nand2_4 _32245_ (.A(_02373_),
    .B(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__o21ai_4 _32246_ (.A1(_20837_),
    .A2(_02523_),
    .B1(_02525_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_4 _32247_ (.A(_02376_),
    .B(_02524_),
    .Y(_02526_));
 sky130_fd_sc_hd__o21ai_4 _32248_ (.A1(_20879_),
    .A2(_02523_),
    .B1(_02526_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_4 _32249_ (.A(_02379_),
    .B(_02524_),
    .Y(_02527_));
 sky130_fd_sc_hd__o21ai_4 _32250_ (.A1(_20926_),
    .A2(_02523_),
    .B1(_02527_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_4 _32251_ (.A(_02382_),
    .B(_02524_),
    .Y(_02528_));
 sky130_fd_sc_hd__o21ai_4 _32252_ (.A1(_20966_),
    .A2(_02523_),
    .B1(_02528_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_4 _32253_ (.A(_02385_),
    .B(_02454_),
    .Y(_02529_));
 sky130_fd_sc_hd__o21ai_4 _32254_ (.A1(_21009_),
    .A2(_02456_),
    .B1(_02529_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand3_4 _32255_ (.A(_01758_),
    .B(_19089_),
    .C(_19094_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor4_4 _32256_ (.A(_19069_),
    .B(_19087_),
    .C(_02530_),
    .D(_01768_),
    .Y(_02531_));
 sky130_vsdinv _32257_ (.A(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__buf_1 _32258_ (.A(_02532_),
    .X(_02533_));
 sky130_fd_sc_hd__buf_1 _32259_ (.A(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__buf_1 _32260_ (.A(_02530_),
    .X(_02535_));
 sky130_fd_sc_hd__nor3_4 _32261_ (.A(_02535_),
    .B(_02391_),
    .C(_01790_),
    .Y(_02536_));
 sky130_fd_sc_hd__a21o_4 _32262_ (.A1(\cpuregs[15][0] ),
    .A2(_02534_),
    .B1(_02536_),
    .X(_00929_));
 sky130_fd_sc_hd__and2_4 _32263_ (.A(_02531_),
    .B(_02395_),
    .X(_02537_));
 sky130_fd_sc_hd__a21o_4 _32264_ (.A1(\cpuregs[15][1] ),
    .A2(_02534_),
    .B1(_02537_),
    .X(_00940_));
 sky130_fd_sc_hd__buf_1 _32265_ (.A(_02532_),
    .X(_02538_));
 sky130_fd_sc_hd__buf_1 _32266_ (.A(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__nor2_4 _32267_ (.A(_02539_),
    .B(_01817_),
    .Y(_02540_));
 sky130_fd_sc_hd__a21o_4 _32268_ (.A1(\cpuregs[15][2] ),
    .A2(_02534_),
    .B1(_02540_),
    .X(_00951_));
 sky130_fd_sc_hd__nor2_4 _32269_ (.A(_02539_),
    .B(_01829_),
    .Y(_02541_));
 sky130_fd_sc_hd__a21o_4 _32270_ (.A1(\cpuregs[15][3] ),
    .A2(_02534_),
    .B1(_02541_),
    .X(_00954_));
 sky130_fd_sc_hd__buf_1 _32271_ (.A(_02533_),
    .X(_02542_));
 sky130_fd_sc_hd__a41oi_4 _32272_ (.A1(_01832_),
    .A2(_01838_),
    .A3(_01841_),
    .A4(_01844_),
    .B1(_02539_),
    .Y(_02543_));
 sky130_fd_sc_hd__a21o_4 _32273_ (.A1(\cpuregs[15][4] ),
    .A2(_02542_),
    .B1(_02543_),
    .X(_00955_));
 sky130_fd_sc_hd__a41oi_4 _32274_ (.A1(_01846_),
    .A2(_01851_),
    .A3(_01854_),
    .A4(_01858_),
    .B1(_02539_),
    .Y(_02544_));
 sky130_fd_sc_hd__a21o_4 _32275_ (.A1(\cpuregs[15][5] ),
    .A2(_02542_),
    .B1(_02544_),
    .X(_00956_));
 sky130_fd_sc_hd__buf_1 _32276_ (.A(_02532_),
    .X(_02545_));
 sky130_fd_sc_hd__buf_1 _32277_ (.A(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__a41oi_4 _32278_ (.A1(_01860_),
    .A2(_01866_),
    .A3(_01869_),
    .A4(_01872_),
    .B1(_02546_),
    .Y(_02547_));
 sky130_fd_sc_hd__a21o_4 _32279_ (.A1(\cpuregs[15][6] ),
    .A2(_02542_),
    .B1(_02547_),
    .X(_00957_));
 sky130_fd_sc_hd__a41oi_4 _32280_ (.A1(_01876_),
    .A2(_01882_),
    .A3(_01886_),
    .A4(_01889_),
    .B1(_02546_),
    .Y(_02548_));
 sky130_fd_sc_hd__a21o_4 _32281_ (.A1(\cpuregs[15][7] ),
    .A2(_02542_),
    .B1(_02548_),
    .X(_00958_));
 sky130_fd_sc_hd__buf_1 _32282_ (.A(_02533_),
    .X(_02549_));
 sky130_fd_sc_hd__a41oi_4 _32283_ (.A1(_01892_),
    .A2(_01896_),
    .A3(_01899_),
    .A4(_01902_),
    .B1(_02546_),
    .Y(_02550_));
 sky130_fd_sc_hd__a21o_4 _32284_ (.A1(\cpuregs[15][8] ),
    .A2(_02549_),
    .B1(_02550_),
    .X(_00959_));
 sky130_fd_sc_hd__a41oi_4 _32285_ (.A1(_01904_),
    .A2(_01909_),
    .A3(_01912_),
    .A4(_01917_),
    .B1(_02546_),
    .Y(_02551_));
 sky130_fd_sc_hd__a21o_4 _32286_ (.A1(\cpuregs[15][9] ),
    .A2(_02549_),
    .B1(_02551_),
    .X(_00960_));
 sky130_fd_sc_hd__buf_1 _32287_ (.A(_02545_),
    .X(_02552_));
 sky130_fd_sc_hd__a41oi_4 _32288_ (.A1(_01919_),
    .A2(_01924_),
    .A3(_01927_),
    .A4(_01930_),
    .B1(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__a21o_4 _32289_ (.A1(\cpuregs[15][10] ),
    .A2(_02549_),
    .B1(_02553_),
    .X(_00930_));
 sky130_fd_sc_hd__a41oi_4 _32290_ (.A1(_01933_),
    .A2(_01939_),
    .A3(_01943_),
    .A4(_01946_),
    .B1(_02552_),
    .Y(_02554_));
 sky130_fd_sc_hd__a21o_4 _32291_ (.A1(\cpuregs[15][11] ),
    .A2(_02549_),
    .B1(_02554_),
    .X(_00931_));
 sky130_fd_sc_hd__buf_1 _32292_ (.A(_02532_),
    .X(_02555_));
 sky130_fd_sc_hd__buf_1 _32293_ (.A(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__a41oi_4 _32294_ (.A1(_01950_),
    .A2(_01954_),
    .A3(_01957_),
    .A4(_01960_),
    .B1(_02552_),
    .Y(_02557_));
 sky130_fd_sc_hd__a21o_4 _32295_ (.A1(\cpuregs[15][12] ),
    .A2(_02556_),
    .B1(_02557_),
    .X(_00932_));
 sky130_fd_sc_hd__a41oi_4 _32296_ (.A1(_01962_),
    .A2(_01968_),
    .A3(_01971_),
    .A4(_01975_),
    .B1(_02552_),
    .Y(_02558_));
 sky130_fd_sc_hd__a21o_4 _32297_ (.A1(\cpuregs[15][13] ),
    .A2(_02556_),
    .B1(_02558_),
    .X(_00933_));
 sky130_fd_sc_hd__buf_1 _32298_ (.A(_02545_),
    .X(_02559_));
 sky130_fd_sc_hd__a41oi_4 _32299_ (.A1(_01977_),
    .A2(_01984_),
    .A3(_01987_),
    .A4(_01990_),
    .B1(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__a21o_4 _32300_ (.A1(\cpuregs[15][14] ),
    .A2(_02556_),
    .B1(_02560_),
    .X(_00934_));
 sky130_fd_sc_hd__a41oi_4 _32301_ (.A1(_01993_),
    .A2(_02000_),
    .A3(_02004_),
    .A4(_02007_),
    .B1(_02559_),
    .Y(_02561_));
 sky130_fd_sc_hd__a21o_4 _32302_ (.A1(\cpuregs[15][15] ),
    .A2(_02556_),
    .B1(_02561_),
    .X(_00935_));
 sky130_fd_sc_hd__buf_1 _32303_ (.A(_02555_),
    .X(_02562_));
 sky130_fd_sc_hd__a41oi_4 _32304_ (.A1(_02010_),
    .A2(_02017_),
    .A3(_02020_),
    .A4(_02023_),
    .B1(_02559_),
    .Y(_02563_));
 sky130_fd_sc_hd__a21o_4 _32305_ (.A1(\cpuregs[15][16] ),
    .A2(_02562_),
    .B1(_02563_),
    .X(_00936_));
 sky130_fd_sc_hd__a41oi_4 _32306_ (.A1(_02025_),
    .A2(_02032_),
    .A3(_02035_),
    .A4(_02039_),
    .B1(_02559_),
    .Y(_02564_));
 sky130_fd_sc_hd__a21o_4 _32307_ (.A1(\cpuregs[15][17] ),
    .A2(_02562_),
    .B1(_02564_),
    .X(_00937_));
 sky130_fd_sc_hd__buf_1 _32308_ (.A(_02538_),
    .X(_02565_));
 sky130_fd_sc_hd__a41oi_4 _32309_ (.A1(_02041_),
    .A2(_02045_),
    .A3(_02049_),
    .A4(_02052_),
    .B1(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21o_4 _32310_ (.A1(\cpuregs[15][18] ),
    .A2(_02562_),
    .B1(_02566_),
    .X(_00938_));
 sky130_fd_sc_hd__a41oi_4 _32311_ (.A1(_02055_),
    .A2(_02062_),
    .A3(_02065_),
    .A4(_02068_),
    .B1(_02565_),
    .Y(_02567_));
 sky130_fd_sc_hd__a21o_4 _32312_ (.A1(\cpuregs[15][19] ),
    .A2(_02562_),
    .B1(_02567_),
    .X(_00939_));
 sky130_fd_sc_hd__buf_1 _32313_ (.A(_02555_),
    .X(_02568_));
 sky130_fd_sc_hd__a41oi_4 _32314_ (.A1(_02071_),
    .A2(_02078_),
    .A3(_02082_),
    .A4(_02085_),
    .B1(_02565_),
    .Y(_02569_));
 sky130_fd_sc_hd__a21o_4 _32315_ (.A1(\cpuregs[15][20] ),
    .A2(_02568_),
    .B1(_02569_),
    .X(_00941_));
 sky130_fd_sc_hd__a41oi_4 _32316_ (.A1(_02087_),
    .A2(_02093_),
    .A3(_02096_),
    .A4(_02099_),
    .B1(_02565_),
    .Y(_02570_));
 sky130_fd_sc_hd__a21o_4 _32317_ (.A1(\cpuregs[15][21] ),
    .A2(_02568_),
    .B1(_02570_),
    .X(_00942_));
 sky130_fd_sc_hd__buf_1 _32318_ (.A(_02538_),
    .X(_02571_));
 sky130_fd_sc_hd__a41oi_4 _32319_ (.A1(_02101_),
    .A2(_02106_),
    .A3(_02109_),
    .A4(_02113_),
    .B1(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__a21o_4 _32320_ (.A1(\cpuregs[15][22] ),
    .A2(_02568_),
    .B1(_02572_),
    .X(_00943_));
 sky130_fd_sc_hd__a41oi_4 _32321_ (.A1(_02116_),
    .A2(_02123_),
    .A3(_02126_),
    .A4(_02130_),
    .B1(_02571_),
    .Y(_02573_));
 sky130_fd_sc_hd__a21o_4 _32322_ (.A1(\cpuregs[15][23] ),
    .A2(_02568_),
    .B1(_02573_),
    .X(_00944_));
 sky130_fd_sc_hd__buf_1 _32323_ (.A(_02555_),
    .X(_02574_));
 sky130_fd_sc_hd__a41oi_4 _32324_ (.A1(_02133_),
    .A2(_02140_),
    .A3(_02143_),
    .A4(_02146_),
    .B1(_02571_),
    .Y(_02575_));
 sky130_fd_sc_hd__a21o_4 _32325_ (.A1(\cpuregs[15][24] ),
    .A2(_02574_),
    .B1(_02575_),
    .X(_00945_));
 sky130_fd_sc_hd__a41oi_4 _32326_ (.A1(_02148_),
    .A2(_02155_),
    .A3(_02158_),
    .A4(_02161_),
    .B1(_02571_),
    .Y(_02576_));
 sky130_fd_sc_hd__a21o_4 _32327_ (.A1(\cpuregs[15][25] ),
    .A2(_02574_),
    .B1(_02576_),
    .X(_00946_));
 sky130_fd_sc_hd__buf_1 _32328_ (.A(_02538_),
    .X(_02577_));
 sky130_fd_sc_hd__a41oi_4 _32329_ (.A1(_02163_),
    .A2(_02169_),
    .A3(_02172_),
    .A4(_02175_),
    .B1(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__a21o_4 _32330_ (.A1(\cpuregs[15][26] ),
    .A2(_02574_),
    .B1(_02578_),
    .X(_00947_));
 sky130_fd_sc_hd__a41oi_4 _32331_ (.A1(_02178_),
    .A2(_02184_),
    .A3(_02187_),
    .A4(_02190_),
    .B1(_02577_),
    .Y(_02579_));
 sky130_fd_sc_hd__a21o_4 _32332_ (.A1(\cpuregs[15][27] ),
    .A2(_02574_),
    .B1(_02579_),
    .X(_00948_));
 sky130_fd_sc_hd__buf_1 _32333_ (.A(_02545_),
    .X(_02580_));
 sky130_fd_sc_hd__and2_4 _32334_ (.A(_02198_),
    .B(_02531_),
    .X(_02581_));
 sky130_fd_sc_hd__a21o_4 _32335_ (.A1(\cpuregs[15][28] ),
    .A2(_02580_),
    .B1(_02581_),
    .X(_00949_));
 sky130_fd_sc_hd__a41oi_4 _32336_ (.A1(_02200_),
    .A2(_02206_),
    .A3(_02209_),
    .A4(_02212_),
    .B1(_02577_),
    .Y(_02582_));
 sky130_fd_sc_hd__a21o_4 _32337_ (.A1(\cpuregs[15][29] ),
    .A2(_02580_),
    .B1(_02582_),
    .X(_00950_));
 sky130_fd_sc_hd__a41oi_4 _32338_ (.A1(_02214_),
    .A2(_02219_),
    .A3(_02222_),
    .A4(_02225_),
    .B1(_02577_),
    .Y(_02583_));
 sky130_fd_sc_hd__a21o_4 _32339_ (.A1(\cpuregs[15][30] ),
    .A2(_02580_),
    .B1(_02583_),
    .X(_00952_));
 sky130_fd_sc_hd__a41oi_4 _32340_ (.A1(_02227_),
    .A2(_02233_),
    .A3(_02236_),
    .A4(_02239_),
    .B1(_02533_),
    .Y(_02584_));
 sky130_fd_sc_hd__a21o_4 _32341_ (.A1(\cpuregs[15][31] ),
    .A2(_02580_),
    .B1(_02584_),
    .X(_00953_));
 sky130_vsdinv _32342_ (.A(_02530_),
    .Y(_02585_));
 sky130_fd_sc_hd__and4_4 _32343_ (.A(_02241_),
    .B(_01788_),
    .C(_02242_),
    .D(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__buf_1 _32344_ (.A(_02586_),
    .X(_02587_));
 sky130_vsdinv _32345_ (.A(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__buf_1 _32346_ (.A(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__buf_1 _32347_ (.A(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__nor2_4 _32348_ (.A(_02249_),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__a21o_4 _32349_ (.A1(\cpuregs[14][0] ),
    .A2(_02590_),
    .B1(_02591_),
    .X(_00897_));
 sky130_fd_sc_hd__buf_1 _32350_ (.A(_02587_),
    .X(_02592_));
 sky130_fd_sc_hd__buf_1 _32351_ (.A(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__buf_1 _32352_ (.A(_02587_),
    .X(_02594_));
 sky130_fd_sc_hd__buf_1 _32353_ (.A(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__nand2_4 _32354_ (.A(_02254_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__o21ai_4 _32355_ (.A1(_19288_),
    .A2(_02593_),
    .B1(_02596_),
    .Y(_00908_));
 sky130_fd_sc_hd__buf_1 _32356_ (.A(_23472_),
    .X(_02597_));
 sky130_fd_sc_hd__a41o_4 _32357_ (.A1(_02258_),
    .A2(_02597_),
    .A3(_02259_),
    .A4(_02260_),
    .B1(_02590_),
    .X(_02598_));
 sky130_fd_sc_hd__o21ai_4 _32358_ (.A1(_19435_),
    .A2(_02593_),
    .B1(_02598_),
    .Y(_00919_));
 sky130_fd_sc_hd__buf_1 _32359_ (.A(_23477_),
    .X(_02599_));
 sky130_fd_sc_hd__a41o_4 _32360_ (.A1(_02599_),
    .A2(_02263_),
    .A3(_02265_),
    .A4(_02267_),
    .B1(_02590_),
    .X(_02600_));
 sky130_fd_sc_hd__o21ai_4 _32361_ (.A1(_19502_),
    .A2(_02593_),
    .B1(_02600_),
    .Y(_00922_));
 sky130_fd_sc_hd__buf_1 _32362_ (.A(_01836_),
    .X(_02601_));
 sky130_fd_sc_hd__buf_1 _32363_ (.A(_01839_),
    .X(_02602_));
 sky130_fd_sc_hd__buf_1 _32364_ (.A(_01842_),
    .X(_02603_));
 sky130_fd_sc_hd__buf_1 _32365_ (.A(_02589_),
    .X(_02604_));
 sky130_fd_sc_hd__a41o_4 _32366_ (.A1(_02601_),
    .A2(_02468_),
    .A3(_02602_),
    .A4(_02603_),
    .B1(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__o21ai_4 _32367_ (.A1(_19572_),
    .A2(_02593_),
    .B1(_02605_),
    .Y(_00923_));
 sky130_fd_sc_hd__buf_1 _32368_ (.A(_02587_),
    .X(_02606_));
 sky130_fd_sc_hd__buf_1 _32369_ (.A(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__buf_1 _32370_ (.A(_01849_),
    .X(_02608_));
 sky130_fd_sc_hd__buf_1 _32371_ (.A(_01852_),
    .X(_02609_));
 sky130_fd_sc_hd__buf_1 _32372_ (.A(_01856_),
    .X(_02610_));
 sky130_fd_sc_hd__a41o_4 _32373_ (.A1(_02608_),
    .A2(_02470_),
    .A3(_02609_),
    .A4(_02610_),
    .B1(_02604_),
    .X(_02611_));
 sky130_fd_sc_hd__o21ai_4 _32374_ (.A1(_19654_),
    .A2(_02607_),
    .B1(_02611_),
    .Y(_00924_));
 sky130_fd_sc_hd__buf_1 _32375_ (.A(_01864_),
    .X(_02612_));
 sky130_fd_sc_hd__buf_1 _32376_ (.A(_01867_),
    .X(_02613_));
 sky130_fd_sc_hd__buf_1 _32377_ (.A(_01870_),
    .X(_02614_));
 sky130_fd_sc_hd__a41o_4 _32378_ (.A1(_02612_),
    .A2(_02472_),
    .A3(_02613_),
    .A4(_02614_),
    .B1(_02604_),
    .X(_02615_));
 sky130_fd_sc_hd__o21ai_4 _32379_ (.A1(_19699_),
    .A2(_02607_),
    .B1(_02615_),
    .Y(_00925_));
 sky130_fd_sc_hd__buf_1 _32380_ (.A(_01880_),
    .X(_02616_));
 sky130_fd_sc_hd__buf_1 _32381_ (.A(_01884_),
    .X(_02617_));
 sky130_fd_sc_hd__buf_1 _32382_ (.A(_01887_),
    .X(_02618_));
 sky130_fd_sc_hd__a41o_4 _32383_ (.A1(_02616_),
    .A2(_02475_),
    .A3(_02617_),
    .A4(_02618_),
    .B1(_02604_),
    .X(_02619_));
 sky130_fd_sc_hd__o21ai_4 _32384_ (.A1(_19754_),
    .A2(_02607_),
    .B1(_02619_),
    .Y(_00926_));
 sky130_fd_sc_hd__buf_1 _32385_ (.A(_01894_),
    .X(_02620_));
 sky130_fd_sc_hd__buf_1 _32386_ (.A(_01897_),
    .X(_02621_));
 sky130_fd_sc_hd__buf_1 _32387_ (.A(_01900_),
    .X(_02622_));
 sky130_fd_sc_hd__buf_1 _32388_ (.A(_02589_),
    .X(_02623_));
 sky130_fd_sc_hd__a41o_4 _32389_ (.A1(_02620_),
    .A2(_02479_),
    .A3(_02621_),
    .A4(_02622_),
    .B1(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__o21ai_4 _32390_ (.A1(_19806_),
    .A2(_02607_),
    .B1(_02624_),
    .Y(_00927_));
 sky130_fd_sc_hd__buf_1 _32391_ (.A(_02606_),
    .X(_02625_));
 sky130_fd_sc_hd__buf_1 _32392_ (.A(_01907_),
    .X(_02626_));
 sky130_fd_sc_hd__buf_1 _32393_ (.A(_01910_),
    .X(_02627_));
 sky130_fd_sc_hd__buf_1 _32394_ (.A(_01915_),
    .X(_02628_));
 sky130_fd_sc_hd__a41o_4 _32395_ (.A1(_02626_),
    .A2(_02481_),
    .A3(_02627_),
    .A4(_02628_),
    .B1(_02623_),
    .X(_02629_));
 sky130_fd_sc_hd__o21ai_4 _32396_ (.A1(_19869_),
    .A2(_02625_),
    .B1(_02629_),
    .Y(_00928_));
 sky130_fd_sc_hd__buf_1 _32397_ (.A(_01922_),
    .X(_02630_));
 sky130_fd_sc_hd__buf_1 _32398_ (.A(_01925_),
    .X(_02631_));
 sky130_fd_sc_hd__buf_1 _32399_ (.A(_01928_),
    .X(_02632_));
 sky130_fd_sc_hd__a41o_4 _32400_ (.A1(_02630_),
    .A2(_02483_),
    .A3(_02631_),
    .A4(_02632_),
    .B1(_02623_),
    .X(_02633_));
 sky130_fd_sc_hd__o21ai_4 _32401_ (.A1(_19950_),
    .A2(_02625_),
    .B1(_02633_),
    .Y(_00898_));
 sky130_fd_sc_hd__buf_1 _32402_ (.A(_01937_),
    .X(_02634_));
 sky130_fd_sc_hd__buf_1 _32403_ (.A(_01941_),
    .X(_02635_));
 sky130_fd_sc_hd__buf_1 _32404_ (.A(_01944_),
    .X(_02636_));
 sky130_fd_sc_hd__a41o_4 _32405_ (.A1(_02634_),
    .A2(_02486_),
    .A3(_02635_),
    .A4(_02636_),
    .B1(_02623_),
    .X(_02637_));
 sky130_fd_sc_hd__o21ai_4 _32406_ (.A1(_19984_),
    .A2(_02625_),
    .B1(_02637_),
    .Y(_00899_));
 sky130_fd_sc_hd__buf_1 _32407_ (.A(_01952_),
    .X(_02638_));
 sky130_fd_sc_hd__buf_1 _32408_ (.A(_01955_),
    .X(_02639_));
 sky130_fd_sc_hd__buf_1 _32409_ (.A(_01958_),
    .X(_02640_));
 sky130_fd_sc_hd__buf_1 _32410_ (.A(_02588_),
    .X(_02641_));
 sky130_fd_sc_hd__a41o_4 _32411_ (.A1(_02638_),
    .A2(_02489_),
    .A3(_02639_),
    .A4(_02640_),
    .B1(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__o21ai_4 _32412_ (.A1(_20059_),
    .A2(_02625_),
    .B1(_02642_),
    .Y(_00900_));
 sky130_fd_sc_hd__buf_1 _32413_ (.A(_02606_),
    .X(_02643_));
 sky130_fd_sc_hd__buf_1 _32414_ (.A(_01966_),
    .X(_02644_));
 sky130_fd_sc_hd__buf_1 _32415_ (.A(_01969_),
    .X(_02645_));
 sky130_fd_sc_hd__buf_1 _32416_ (.A(_01973_),
    .X(_02646_));
 sky130_fd_sc_hd__a41o_4 _32417_ (.A1(_02644_),
    .A2(_02491_),
    .A3(_02645_),
    .A4(_02646_),
    .B1(_02641_),
    .X(_02647_));
 sky130_fd_sc_hd__o21ai_4 _32418_ (.A1(_20116_),
    .A2(_02643_),
    .B1(_02647_),
    .Y(_00901_));
 sky130_fd_sc_hd__buf_1 _32419_ (.A(_01982_),
    .X(_02648_));
 sky130_fd_sc_hd__buf_1 _32420_ (.A(_01985_),
    .X(_02649_));
 sky130_fd_sc_hd__buf_1 _32421_ (.A(_01988_),
    .X(_02650_));
 sky130_fd_sc_hd__a41o_4 _32422_ (.A1(_02648_),
    .A2(_02493_),
    .A3(_02649_),
    .A4(_02650_),
    .B1(_02641_),
    .X(_02651_));
 sky130_fd_sc_hd__o21ai_4 _32423_ (.A1(_20180_),
    .A2(_02643_),
    .B1(_02651_),
    .Y(_00902_));
 sky130_fd_sc_hd__buf_1 _32424_ (.A(_01998_),
    .X(_02652_));
 sky130_fd_sc_hd__buf_1 _32425_ (.A(_02002_),
    .X(_02653_));
 sky130_fd_sc_hd__buf_1 _32426_ (.A(_02005_),
    .X(_02654_));
 sky130_fd_sc_hd__a41o_4 _32427_ (.A1(_02652_),
    .A2(_02497_),
    .A3(_02653_),
    .A4(_02654_),
    .B1(_02641_),
    .X(_02655_));
 sky130_fd_sc_hd__o21ai_4 _32428_ (.A1(_20236_),
    .A2(_02643_),
    .B1(_02655_),
    .Y(_00903_));
 sky130_fd_sc_hd__buf_1 _32429_ (.A(_02015_),
    .X(_02656_));
 sky130_fd_sc_hd__buf_1 _32430_ (.A(_02018_),
    .X(_02657_));
 sky130_fd_sc_hd__buf_1 _32431_ (.A(_02021_),
    .X(_02658_));
 sky130_fd_sc_hd__buf_1 _32432_ (.A(_02588_),
    .X(_02659_));
 sky130_fd_sc_hd__a41o_4 _32433_ (.A1(_02656_),
    .A2(_02500_),
    .A3(_02657_),
    .A4(_02658_),
    .B1(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__o21ai_4 _32434_ (.A1(_20281_),
    .A2(_02643_),
    .B1(_02660_),
    .Y(_00904_));
 sky130_fd_sc_hd__buf_1 _32435_ (.A(_02606_),
    .X(_02661_));
 sky130_fd_sc_hd__buf_1 _32436_ (.A(_02030_),
    .X(_02662_));
 sky130_fd_sc_hd__buf_1 _32437_ (.A(_02033_),
    .X(_02663_));
 sky130_fd_sc_hd__buf_1 _32438_ (.A(_02037_),
    .X(_02664_));
 sky130_fd_sc_hd__a41o_4 _32439_ (.A1(_02662_),
    .A2(_02502_),
    .A3(_02663_),
    .A4(_02664_),
    .B1(_02659_),
    .X(_02665_));
 sky130_fd_sc_hd__o21ai_4 _32440_ (.A1(_20335_),
    .A2(_02661_),
    .B1(_02665_),
    .Y(_00905_));
 sky130_fd_sc_hd__buf_1 _32441_ (.A(_02594_),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_4 _32442_ (.A(_02335_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__o21ai_4 _32443_ (.A1(_20391_),
    .A2(_02661_),
    .B1(_02667_),
    .Y(_00906_));
 sky130_fd_sc_hd__buf_1 _32444_ (.A(_02060_),
    .X(_02668_));
 sky130_fd_sc_hd__buf_1 _32445_ (.A(_02063_),
    .X(_02669_));
 sky130_fd_sc_hd__buf_1 _32446_ (.A(_02066_),
    .X(_02670_));
 sky130_fd_sc_hd__a41o_4 _32447_ (.A1(_02668_),
    .A2(_02506_),
    .A3(_02669_),
    .A4(_02670_),
    .B1(_02659_),
    .X(_02671_));
 sky130_fd_sc_hd__o21ai_4 _32448_ (.A1(_20439_),
    .A2(_02661_),
    .B1(_02671_),
    .Y(_00907_));
 sky130_fd_sc_hd__buf_1 _32449_ (.A(_02076_),
    .X(_02672_));
 sky130_fd_sc_hd__buf_1 _32450_ (.A(_02080_),
    .X(_02673_));
 sky130_fd_sc_hd__buf_1 _32451_ (.A(_02083_),
    .X(_02674_));
 sky130_fd_sc_hd__a41o_4 _32452_ (.A1(_02672_),
    .A2(_02508_),
    .A3(_02673_),
    .A4(_02674_),
    .B1(_02659_),
    .X(_02675_));
 sky130_fd_sc_hd__o21ai_4 _32453_ (.A1(_20481_),
    .A2(_02661_),
    .B1(_02675_),
    .Y(_00909_));
 sky130_fd_sc_hd__buf_1 _32454_ (.A(_02594_),
    .X(_02676_));
 sky130_fd_sc_hd__buf_1 _32455_ (.A(_02091_),
    .X(_02677_));
 sky130_fd_sc_hd__buf_1 _32456_ (.A(_02094_),
    .X(_02678_));
 sky130_fd_sc_hd__buf_1 _32457_ (.A(_02097_),
    .X(_02679_));
 sky130_fd_sc_hd__buf_1 _32458_ (.A(_02588_),
    .X(_02680_));
 sky130_fd_sc_hd__a41o_4 _32459_ (.A1(_02677_),
    .A2(_02511_),
    .A3(_02678_),
    .A4(_02679_),
    .B1(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__o21ai_4 _32460_ (.A1(_20536_),
    .A2(_02676_),
    .B1(_02681_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand2_4 _32461_ (.A(_02353_),
    .B(_02666_),
    .Y(_02682_));
 sky130_fd_sc_hd__o21ai_4 _32462_ (.A1(_20592_),
    .A2(_02676_),
    .B1(_02682_),
    .Y(_00911_));
 sky130_fd_sc_hd__buf_1 _32463_ (.A(_02121_),
    .X(_02683_));
 sky130_fd_sc_hd__buf_1 _32464_ (.A(_02124_),
    .X(_02684_));
 sky130_fd_sc_hd__buf_1 _32465_ (.A(_02128_),
    .X(_02685_));
 sky130_fd_sc_hd__a41o_4 _32466_ (.A1(_02683_),
    .A2(_02515_),
    .A3(_02684_),
    .A4(_02685_),
    .B1(_02680_),
    .X(_02686_));
 sky130_fd_sc_hd__o21ai_4 _32467_ (.A1(_20619_),
    .A2(_02676_),
    .B1(_02686_),
    .Y(_00912_));
 sky130_fd_sc_hd__buf_1 _32468_ (.A(_02138_),
    .X(_02687_));
 sky130_fd_sc_hd__buf_1 _32469_ (.A(_02141_),
    .X(_02688_));
 sky130_fd_sc_hd__buf_1 _32470_ (.A(_02144_),
    .X(_02689_));
 sky130_fd_sc_hd__a41o_4 _32471_ (.A1(_02687_),
    .A2(_02517_),
    .A3(_02688_),
    .A4(_02689_),
    .B1(_02680_),
    .X(_02690_));
 sky130_fd_sc_hd__o21ai_4 _32472_ (.A1(_20664_),
    .A2(_02676_),
    .B1(_02690_),
    .Y(_00913_));
 sky130_fd_sc_hd__buf_1 _32473_ (.A(_02594_),
    .X(_02691_));
 sky130_fd_sc_hd__buf_1 _32474_ (.A(_02153_),
    .X(_02692_));
 sky130_fd_sc_hd__buf_1 _32475_ (.A(_02156_),
    .X(_02693_));
 sky130_fd_sc_hd__buf_1 _32476_ (.A(_02159_),
    .X(_02694_));
 sky130_fd_sc_hd__a41o_4 _32477_ (.A1(_02692_),
    .A2(_02519_),
    .A3(_02693_),
    .A4(_02694_),
    .B1(_02680_),
    .X(_02695_));
 sky130_fd_sc_hd__o21ai_4 _32478_ (.A1(_20712_),
    .A2(_02691_),
    .B1(_02695_),
    .Y(_00914_));
 sky130_fd_sc_hd__buf_1 _32479_ (.A(_02167_),
    .X(_02696_));
 sky130_fd_sc_hd__buf_1 _32480_ (.A(_02170_),
    .X(_02697_));
 sky130_fd_sc_hd__buf_1 _32481_ (.A(_02173_),
    .X(_02698_));
 sky130_fd_sc_hd__a41o_4 _32482_ (.A1(_02696_),
    .A2(_02521_),
    .A3(_02697_),
    .A4(_02698_),
    .B1(_02589_),
    .X(_02699_));
 sky130_fd_sc_hd__o21ai_4 _32483_ (.A1(_20755_),
    .A2(_02691_),
    .B1(_02699_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand2_4 _32484_ (.A(_02373_),
    .B(_02666_),
    .Y(_02700_));
 sky130_fd_sc_hd__o21ai_4 _32485_ (.A1(_20818_),
    .A2(_02691_),
    .B1(_02700_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand2_4 _32486_ (.A(_02376_),
    .B(_02666_),
    .Y(_02701_));
 sky130_fd_sc_hd__o21ai_4 _32487_ (.A1(_20844_),
    .A2(_02691_),
    .B1(_02701_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_4 _32488_ (.A(_02379_),
    .B(_02592_),
    .Y(_02702_));
 sky130_fd_sc_hd__o21ai_4 _32489_ (.A1(_20893_),
    .A2(_02595_),
    .B1(_02702_),
    .Y(_00918_));
 sky130_fd_sc_hd__nand2_4 _32490_ (.A(_02382_),
    .B(_02592_),
    .Y(_02703_));
 sky130_fd_sc_hd__o21ai_4 _32491_ (.A1(_20933_),
    .A2(_02595_),
    .B1(_02703_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand2_4 _32492_ (.A(_02385_),
    .B(_02592_),
    .Y(_02704_));
 sky130_fd_sc_hd__o21ai_4 _32493_ (.A1(_20976_),
    .A2(_02595_),
    .B1(_02704_),
    .Y(_00921_));
 sky130_fd_sc_hd__buf_1 _32494_ (.A(_19068_),
    .X(_02705_));
 sky130_fd_sc_hd__nor3_4 _32495_ (.A(_19089_),
    .B(_19098_),
    .C(_19095_),
    .Y(_02706_));
 sky130_vsdinv _32496_ (.A(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__nor4_4 _32497_ (.A(_02705_),
    .B(_19086_),
    .C(_02707_),
    .D(_01768_),
    .Y(_02708_));
 sky130_vsdinv _32498_ (.A(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__buf_1 _32499_ (.A(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__buf_1 _32500_ (.A(_02710_),
    .X(_02711_));
 sky130_fd_sc_hd__buf_1 _32501_ (.A(_02707_),
    .X(_02712_));
 sky130_fd_sc_hd__nor3_4 _32502_ (.A(_02712_),
    .B(_02391_),
    .C(_01790_),
    .Y(_02713_));
 sky130_fd_sc_hd__a21o_4 _32503_ (.A1(\cpuregs[11][0] ),
    .A2(_02711_),
    .B1(_02713_),
    .X(_00801_));
 sky130_fd_sc_hd__and2_4 _32504_ (.A(_02708_),
    .B(_02395_),
    .X(_02714_));
 sky130_fd_sc_hd__a21o_4 _32505_ (.A1(\cpuregs[11][1] ),
    .A2(_02711_),
    .B1(_02714_),
    .X(_00812_));
 sky130_fd_sc_hd__buf_1 _32506_ (.A(_02709_),
    .X(_02715_));
 sky130_fd_sc_hd__buf_1 _32507_ (.A(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__nor2_4 _32508_ (.A(_02716_),
    .B(_01817_),
    .Y(_02717_));
 sky130_fd_sc_hd__a21o_4 _32509_ (.A1(\cpuregs[11][2] ),
    .A2(_02711_),
    .B1(_02717_),
    .X(_00823_));
 sky130_fd_sc_hd__buf_1 _32510_ (.A(_01828_),
    .X(_02718_));
 sky130_fd_sc_hd__nor2_4 _32511_ (.A(_02716_),
    .B(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__a21o_4 _32512_ (.A1(\cpuregs[11][3] ),
    .A2(_02711_),
    .B1(_02719_),
    .X(_00826_));
 sky130_fd_sc_hd__buf_1 _32513_ (.A(_02710_),
    .X(_02720_));
 sky130_fd_sc_hd__a41oi_4 _32514_ (.A1(_01832_),
    .A2(_01838_),
    .A3(_01841_),
    .A4(_01844_),
    .B1(_02716_),
    .Y(_02721_));
 sky130_fd_sc_hd__a21o_4 _32515_ (.A1(\cpuregs[11][4] ),
    .A2(_02720_),
    .B1(_02721_),
    .X(_00827_));
 sky130_fd_sc_hd__a41oi_4 _32516_ (.A1(_01846_),
    .A2(_01851_),
    .A3(_01854_),
    .A4(_01858_),
    .B1(_02716_),
    .Y(_02722_));
 sky130_fd_sc_hd__a21o_4 _32517_ (.A1(\cpuregs[11][5] ),
    .A2(_02720_),
    .B1(_02722_),
    .X(_00828_));
 sky130_fd_sc_hd__buf_1 _32518_ (.A(_02709_),
    .X(_02723_));
 sky130_fd_sc_hd__buf_1 _32519_ (.A(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__a41oi_4 _32520_ (.A1(_01860_),
    .A2(_01866_),
    .A3(_01869_),
    .A4(_01872_),
    .B1(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__a21o_4 _32521_ (.A1(\cpuregs[11][6] ),
    .A2(_02720_),
    .B1(_02725_),
    .X(_00829_));
 sky130_fd_sc_hd__a41oi_4 _32522_ (.A1(_01876_),
    .A2(_01882_),
    .A3(_01886_),
    .A4(_01889_),
    .B1(_02724_),
    .Y(_02726_));
 sky130_fd_sc_hd__a21o_4 _32523_ (.A1(\cpuregs[11][7] ),
    .A2(_02720_),
    .B1(_02726_),
    .X(_00830_));
 sky130_fd_sc_hd__buf_1 _32524_ (.A(_02710_),
    .X(_02727_));
 sky130_fd_sc_hd__a41oi_4 _32525_ (.A1(_01892_),
    .A2(_01896_),
    .A3(_01899_),
    .A4(_01902_),
    .B1(_02724_),
    .Y(_02728_));
 sky130_fd_sc_hd__a21o_4 _32526_ (.A1(\cpuregs[11][8] ),
    .A2(_02727_),
    .B1(_02728_),
    .X(_00831_));
 sky130_fd_sc_hd__a41oi_4 _32527_ (.A1(_01904_),
    .A2(_01909_),
    .A3(_01912_),
    .A4(_01917_),
    .B1(_02724_),
    .Y(_02729_));
 sky130_fd_sc_hd__a21o_4 _32528_ (.A1(\cpuregs[11][9] ),
    .A2(_02727_),
    .B1(_02729_),
    .X(_00832_));
 sky130_fd_sc_hd__buf_1 _32529_ (.A(_02723_),
    .X(_02730_));
 sky130_fd_sc_hd__a41oi_4 _32530_ (.A1(_01919_),
    .A2(_01924_),
    .A3(_01927_),
    .A4(_01930_),
    .B1(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__a21o_4 _32531_ (.A1(\cpuregs[11][10] ),
    .A2(_02727_),
    .B1(_02731_),
    .X(_00802_));
 sky130_fd_sc_hd__a41oi_4 _32532_ (.A1(_01933_),
    .A2(_01939_),
    .A3(_01943_),
    .A4(_01946_),
    .B1(_02730_),
    .Y(_02732_));
 sky130_fd_sc_hd__a21o_4 _32533_ (.A1(\cpuregs[11][11] ),
    .A2(_02727_),
    .B1(_02732_),
    .X(_00803_));
 sky130_fd_sc_hd__buf_1 _32534_ (.A(_02709_),
    .X(_02733_));
 sky130_fd_sc_hd__buf_1 _32535_ (.A(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__a41oi_4 _32536_ (.A1(_01950_),
    .A2(_01954_),
    .A3(_01957_),
    .A4(_01960_),
    .B1(_02730_),
    .Y(_02735_));
 sky130_fd_sc_hd__a21o_4 _32537_ (.A1(\cpuregs[11][12] ),
    .A2(_02734_),
    .B1(_02735_),
    .X(_00804_));
 sky130_fd_sc_hd__a41oi_4 _32538_ (.A1(_01962_),
    .A2(_01968_),
    .A3(_01971_),
    .A4(_01975_),
    .B1(_02730_),
    .Y(_02736_));
 sky130_fd_sc_hd__a21o_4 _32539_ (.A1(\cpuregs[11][13] ),
    .A2(_02734_),
    .B1(_02736_),
    .X(_00805_));
 sky130_fd_sc_hd__buf_1 _32540_ (.A(_02723_),
    .X(_02737_));
 sky130_fd_sc_hd__a41oi_4 _32541_ (.A1(_01977_),
    .A2(_01984_),
    .A3(_01987_),
    .A4(_01990_),
    .B1(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__a21o_4 _32542_ (.A1(\cpuregs[11][14] ),
    .A2(_02734_),
    .B1(_02738_),
    .X(_00806_));
 sky130_fd_sc_hd__a41oi_4 _32543_ (.A1(_01993_),
    .A2(_02000_),
    .A3(_02004_),
    .A4(_02007_),
    .B1(_02737_),
    .Y(_02739_));
 sky130_fd_sc_hd__a21o_4 _32544_ (.A1(\cpuregs[11][15] ),
    .A2(_02734_),
    .B1(_02739_),
    .X(_00807_));
 sky130_fd_sc_hd__buf_1 _32545_ (.A(_02733_),
    .X(_02740_));
 sky130_fd_sc_hd__a41oi_4 _32546_ (.A1(_02010_),
    .A2(_02017_),
    .A3(_02020_),
    .A4(_02023_),
    .B1(_02737_),
    .Y(_02741_));
 sky130_fd_sc_hd__a21o_4 _32547_ (.A1(\cpuregs[11][16] ),
    .A2(_02740_),
    .B1(_02741_),
    .X(_00808_));
 sky130_fd_sc_hd__a41oi_4 _32548_ (.A1(_02025_),
    .A2(_02032_),
    .A3(_02035_),
    .A4(_02039_),
    .B1(_02737_),
    .Y(_02742_));
 sky130_fd_sc_hd__a21o_4 _32549_ (.A1(\cpuregs[11][17] ),
    .A2(_02740_),
    .B1(_02742_),
    .X(_00809_));
 sky130_fd_sc_hd__buf_1 _32550_ (.A(_02715_),
    .X(_02743_));
 sky130_fd_sc_hd__a41oi_4 _32551_ (.A1(_02041_),
    .A2(_02045_),
    .A3(_02049_),
    .A4(_02052_),
    .B1(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__a21o_4 _32552_ (.A1(\cpuregs[11][18] ),
    .A2(_02740_),
    .B1(_02744_),
    .X(_00810_));
 sky130_fd_sc_hd__a41oi_4 _32553_ (.A1(_02055_),
    .A2(_02062_),
    .A3(_02065_),
    .A4(_02068_),
    .B1(_02743_),
    .Y(_02745_));
 sky130_fd_sc_hd__a21o_4 _32554_ (.A1(\cpuregs[11][19] ),
    .A2(_02740_),
    .B1(_02745_),
    .X(_00811_));
 sky130_fd_sc_hd__buf_1 _32555_ (.A(_02733_),
    .X(_02746_));
 sky130_fd_sc_hd__a41oi_4 _32556_ (.A1(_02071_),
    .A2(_02078_),
    .A3(_02082_),
    .A4(_02085_),
    .B1(_02743_),
    .Y(_02747_));
 sky130_fd_sc_hd__a21o_4 _32557_ (.A1(\cpuregs[11][20] ),
    .A2(_02746_),
    .B1(_02747_),
    .X(_00813_));
 sky130_fd_sc_hd__a41oi_4 _32558_ (.A1(_02087_),
    .A2(_02093_),
    .A3(_02096_),
    .A4(_02099_),
    .B1(_02743_),
    .Y(_02748_));
 sky130_fd_sc_hd__a21o_4 _32559_ (.A1(\cpuregs[11][21] ),
    .A2(_02746_),
    .B1(_02748_),
    .X(_00814_));
 sky130_fd_sc_hd__buf_1 _32560_ (.A(_02715_),
    .X(_02749_));
 sky130_fd_sc_hd__a41oi_4 _32561_ (.A1(_02101_),
    .A2(_02106_),
    .A3(_02109_),
    .A4(_02113_),
    .B1(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__a21o_4 _32562_ (.A1(\cpuregs[11][22] ),
    .A2(_02746_),
    .B1(_02750_),
    .X(_00815_));
 sky130_fd_sc_hd__a41oi_4 _32563_ (.A1(_02116_),
    .A2(_02123_),
    .A3(_02126_),
    .A4(_02130_),
    .B1(_02749_),
    .Y(_02751_));
 sky130_fd_sc_hd__a21o_4 _32564_ (.A1(\cpuregs[11][23] ),
    .A2(_02746_),
    .B1(_02751_),
    .X(_00816_));
 sky130_fd_sc_hd__buf_1 _32565_ (.A(_02733_),
    .X(_02752_));
 sky130_fd_sc_hd__a41oi_4 _32566_ (.A1(_02133_),
    .A2(_02140_),
    .A3(_02143_),
    .A4(_02146_),
    .B1(_02749_),
    .Y(_02753_));
 sky130_fd_sc_hd__a21o_4 _32567_ (.A1(\cpuregs[11][24] ),
    .A2(_02752_),
    .B1(_02753_),
    .X(_00817_));
 sky130_fd_sc_hd__a41oi_4 _32568_ (.A1(_02148_),
    .A2(_02155_),
    .A3(_02158_),
    .A4(_02161_),
    .B1(_02749_),
    .Y(_02754_));
 sky130_fd_sc_hd__a21o_4 _32569_ (.A1(\cpuregs[11][25] ),
    .A2(_02752_),
    .B1(_02754_),
    .X(_00818_));
 sky130_fd_sc_hd__buf_1 _32570_ (.A(_02715_),
    .X(_02755_));
 sky130_fd_sc_hd__a41oi_4 _32571_ (.A1(_02163_),
    .A2(_02169_),
    .A3(_02172_),
    .A4(_02175_),
    .B1(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__a21o_4 _32572_ (.A1(\cpuregs[11][26] ),
    .A2(_02752_),
    .B1(_02756_),
    .X(_00819_));
 sky130_fd_sc_hd__a41oi_4 _32573_ (.A1(_02178_),
    .A2(_02184_),
    .A3(_02187_),
    .A4(_02190_),
    .B1(_02755_),
    .Y(_02757_));
 sky130_fd_sc_hd__a21o_4 _32574_ (.A1(\cpuregs[11][27] ),
    .A2(_02752_),
    .B1(_02757_),
    .X(_00820_));
 sky130_fd_sc_hd__buf_1 _32575_ (.A(_02723_),
    .X(_02758_));
 sky130_fd_sc_hd__buf_1 _32576_ (.A(_02197_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_4 _32577_ (.A(_02759_),
    .B(_02708_),
    .X(_02760_));
 sky130_fd_sc_hd__a21o_4 _32578_ (.A1(\cpuregs[11][28] ),
    .A2(_02758_),
    .B1(_02760_),
    .X(_00821_));
 sky130_fd_sc_hd__a41oi_4 _32579_ (.A1(_02200_),
    .A2(_02206_),
    .A3(_02209_),
    .A4(_02212_),
    .B1(_02755_),
    .Y(_02761_));
 sky130_fd_sc_hd__a21o_4 _32580_ (.A1(\cpuregs[11][29] ),
    .A2(_02758_),
    .B1(_02761_),
    .X(_00822_));
 sky130_fd_sc_hd__a41oi_4 _32581_ (.A1(_02214_),
    .A2(_02219_),
    .A3(_02222_),
    .A4(_02225_),
    .B1(_02755_),
    .Y(_02762_));
 sky130_fd_sc_hd__a21o_4 _32582_ (.A1(\cpuregs[11][30] ),
    .A2(_02758_),
    .B1(_02762_),
    .X(_00824_));
 sky130_fd_sc_hd__a41oi_4 _32583_ (.A1(_02227_),
    .A2(_02233_),
    .A3(_02236_),
    .A4(_02239_),
    .B1(_02710_),
    .Y(_02763_));
 sky130_fd_sc_hd__a21o_4 _32584_ (.A1(\cpuregs[11][31] ),
    .A2(_02758_),
    .B1(_02763_),
    .X(_00825_));
 sky130_fd_sc_hd__and4_4 _32585_ (.A(_02241_),
    .B(_01788_),
    .C(_02242_),
    .D(_02706_),
    .X(_02764_));
 sky130_fd_sc_hd__buf_1 _32586_ (.A(_02764_),
    .X(_02765_));
 sky130_vsdinv _32587_ (.A(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__buf_1 _32588_ (.A(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__buf_1 _32589_ (.A(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__nor2_4 _32590_ (.A(_02249_),
    .B(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__a21o_4 _32591_ (.A1(\cpuregs[10][0] ),
    .A2(_02768_),
    .B1(_02769_),
    .X(_00769_));
 sky130_fd_sc_hd__buf_1 _32592_ (.A(_02765_),
    .X(_02770_));
 sky130_fd_sc_hd__buf_1 _32593_ (.A(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__buf_1 _32594_ (.A(_02765_),
    .X(_02772_));
 sky130_fd_sc_hd__buf_1 _32595_ (.A(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_4 _32596_ (.A(_02254_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__o21ai_4 _32597_ (.A1(_19321_),
    .A2(_02771_),
    .B1(_02774_),
    .Y(_00780_));
 sky130_fd_sc_hd__a41o_4 _32598_ (.A1(_02459_),
    .A2(_02597_),
    .A3(_02461_),
    .A4(_02463_),
    .B1(_02768_),
    .X(_02775_));
 sky130_fd_sc_hd__o21ai_4 _32599_ (.A1(_19443_),
    .A2(_02771_),
    .B1(_02775_),
    .Y(_00791_));
 sky130_fd_sc_hd__a41o_4 _32600_ (.A1(_02599_),
    .A2(_02262_),
    .A3(_02264_),
    .A4(_02266_),
    .B1(_02768_),
    .X(_02776_));
 sky130_fd_sc_hd__o21ai_4 _32601_ (.A1(_19514_),
    .A2(_02771_),
    .B1(_02776_),
    .Y(_00794_));
 sky130_fd_sc_hd__buf_1 _32602_ (.A(_02767_),
    .X(_02777_));
 sky130_fd_sc_hd__a41o_4 _32603_ (.A1(_02601_),
    .A2(_02468_),
    .A3(_02602_),
    .A4(_02603_),
    .B1(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__o21ai_4 _32604_ (.A1(_19595_),
    .A2(_02771_),
    .B1(_02778_),
    .Y(_00795_));
 sky130_fd_sc_hd__buf_1 _32605_ (.A(_02765_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_1 _32606_ (.A(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__a41o_4 _32607_ (.A1(_02608_),
    .A2(_02470_),
    .A3(_02609_),
    .A4(_02610_),
    .B1(_02777_),
    .X(_02781_));
 sky130_fd_sc_hd__o21ai_4 _32608_ (.A1(_19666_),
    .A2(_02780_),
    .B1(_02781_),
    .Y(_00796_));
 sky130_fd_sc_hd__a41o_4 _32609_ (.A1(_02612_),
    .A2(_02472_),
    .A3(_02613_),
    .A4(_02614_),
    .B1(_02777_),
    .X(_02782_));
 sky130_fd_sc_hd__o21ai_4 _32610_ (.A1(_19712_),
    .A2(_02780_),
    .B1(_02782_),
    .Y(_00797_));
 sky130_fd_sc_hd__a41o_4 _32611_ (.A1(_02616_),
    .A2(_02475_),
    .A3(_02617_),
    .A4(_02618_),
    .B1(_02777_),
    .X(_02783_));
 sky130_fd_sc_hd__o21ai_4 _32612_ (.A1(_19765_),
    .A2(_02780_),
    .B1(_02783_),
    .Y(_00798_));
 sky130_fd_sc_hd__buf_1 _32613_ (.A(_02767_),
    .X(_02784_));
 sky130_fd_sc_hd__a41o_4 _32614_ (.A1(_02620_),
    .A2(_02479_),
    .A3(_02621_),
    .A4(_02622_),
    .B1(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__o21ai_4 _32615_ (.A1(_19823_),
    .A2(_02780_),
    .B1(_02785_),
    .Y(_00799_));
 sky130_fd_sc_hd__buf_1 _32616_ (.A(_02779_),
    .X(_02786_));
 sky130_fd_sc_hd__a41o_4 _32617_ (.A1(_02626_),
    .A2(_02481_),
    .A3(_02627_),
    .A4(_02628_),
    .B1(_02784_),
    .X(_02787_));
 sky130_fd_sc_hd__o21ai_4 _32618_ (.A1(_19881_),
    .A2(_02786_),
    .B1(_02787_),
    .Y(_00800_));
 sky130_fd_sc_hd__a41o_4 _32619_ (.A1(_02630_),
    .A2(_02483_),
    .A3(_02631_),
    .A4(_02632_),
    .B1(_02784_),
    .X(_02788_));
 sky130_fd_sc_hd__o21ai_4 _32620_ (.A1(_19960_),
    .A2(_02786_),
    .B1(_02788_),
    .Y(_00770_));
 sky130_fd_sc_hd__a41o_4 _32621_ (.A1(_02634_),
    .A2(_02486_),
    .A3(_02635_),
    .A4(_02636_),
    .B1(_02784_),
    .X(_02789_));
 sky130_fd_sc_hd__o21ai_4 _32622_ (.A1(_19998_),
    .A2(_02786_),
    .B1(_02789_),
    .Y(_00771_));
 sky130_fd_sc_hd__buf_1 _32623_ (.A(_02766_),
    .X(_02790_));
 sky130_fd_sc_hd__a41o_4 _32624_ (.A1(_02638_),
    .A2(_02489_),
    .A3(_02639_),
    .A4(_02640_),
    .B1(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__o21ai_4 _32625_ (.A1(_20072_),
    .A2(_02786_),
    .B1(_02791_),
    .Y(_00772_));
 sky130_fd_sc_hd__buf_1 _32626_ (.A(_02779_),
    .X(_02792_));
 sky130_fd_sc_hd__a41o_4 _32627_ (.A1(_02644_),
    .A2(_02491_),
    .A3(_02645_),
    .A4(_02646_),
    .B1(_02790_),
    .X(_02793_));
 sky130_fd_sc_hd__o21ai_4 _32628_ (.A1(_20129_),
    .A2(_02792_),
    .B1(_02793_),
    .Y(_00773_));
 sky130_fd_sc_hd__a41o_4 _32629_ (.A1(_02648_),
    .A2(_02493_),
    .A3(_02649_),
    .A4(_02650_),
    .B1(_02790_),
    .X(_02794_));
 sky130_fd_sc_hd__o21ai_4 _32630_ (.A1(_20193_),
    .A2(_02792_),
    .B1(_02794_),
    .Y(_00774_));
 sky130_fd_sc_hd__a41o_4 _32631_ (.A1(_02652_),
    .A2(_02497_),
    .A3(_02653_),
    .A4(_02654_),
    .B1(_02790_),
    .X(_02795_));
 sky130_fd_sc_hd__o21ai_4 _32632_ (.A1(_20246_),
    .A2(_02792_),
    .B1(_02795_),
    .Y(_00775_));
 sky130_fd_sc_hd__buf_1 _32633_ (.A(_02766_),
    .X(_02796_));
 sky130_fd_sc_hd__a41o_4 _32634_ (.A1(_02656_),
    .A2(_02500_),
    .A3(_02657_),
    .A4(_02658_),
    .B1(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__o21ai_4 _32635_ (.A1(_20292_),
    .A2(_02792_),
    .B1(_02797_),
    .Y(_00776_));
 sky130_fd_sc_hd__buf_1 _32636_ (.A(_02779_),
    .X(_02798_));
 sky130_fd_sc_hd__a41o_4 _32637_ (.A1(_02662_),
    .A2(_02502_),
    .A3(_02663_),
    .A4(_02664_),
    .B1(_02796_),
    .X(_02799_));
 sky130_fd_sc_hd__o21ai_4 _32638_ (.A1(_20346_),
    .A2(_02798_),
    .B1(_02799_),
    .Y(_00777_));
 sky130_fd_sc_hd__buf_1 _32639_ (.A(_02772_),
    .X(_02800_));
 sky130_fd_sc_hd__nand2_4 _32640_ (.A(_02335_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__o21ai_4 _32641_ (.A1(_20401_),
    .A2(_02798_),
    .B1(_02801_),
    .Y(_00778_));
 sky130_fd_sc_hd__a41o_4 _32642_ (.A1(_02668_),
    .A2(_02506_),
    .A3(_02669_),
    .A4(_02670_),
    .B1(_02796_),
    .X(_02802_));
 sky130_fd_sc_hd__o21ai_4 _32643_ (.A1(_20451_),
    .A2(_02798_),
    .B1(_02802_),
    .Y(_00779_));
 sky130_fd_sc_hd__a41o_4 _32644_ (.A1(_02672_),
    .A2(_02508_),
    .A3(_02673_),
    .A4(_02674_),
    .B1(_02796_),
    .X(_02803_));
 sky130_fd_sc_hd__o21ai_4 _32645_ (.A1(_20493_),
    .A2(_02798_),
    .B1(_02803_),
    .Y(_00781_));
 sky130_fd_sc_hd__buf_1 _32646_ (.A(_02772_),
    .X(_02804_));
 sky130_fd_sc_hd__buf_1 _32647_ (.A(_02766_),
    .X(_02805_));
 sky130_fd_sc_hd__a41o_4 _32648_ (.A1(_02677_),
    .A2(_02511_),
    .A3(_02678_),
    .A4(_02679_),
    .B1(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__o21ai_4 _32649_ (.A1(_20546_),
    .A2(_02804_),
    .B1(_02806_),
    .Y(_00782_));
 sky130_fd_sc_hd__nand2_4 _32650_ (.A(_02353_),
    .B(_02800_),
    .Y(_02807_));
 sky130_fd_sc_hd__o21ai_4 _32651_ (.A1(_20602_),
    .A2(_02804_),
    .B1(_02807_),
    .Y(_00783_));
 sky130_fd_sc_hd__a41o_4 _32652_ (.A1(_02683_),
    .A2(_02515_),
    .A3(_02684_),
    .A4(_02685_),
    .B1(_02805_),
    .X(_02808_));
 sky130_fd_sc_hd__o21ai_4 _32653_ (.A1(_20629_),
    .A2(_02804_),
    .B1(_02808_),
    .Y(_00784_));
 sky130_fd_sc_hd__a41o_4 _32654_ (.A1(_02687_),
    .A2(_02517_),
    .A3(_02688_),
    .A4(_02689_),
    .B1(_02805_),
    .X(_02809_));
 sky130_fd_sc_hd__o21ai_4 _32655_ (.A1(_20674_),
    .A2(_02804_),
    .B1(_02809_),
    .Y(_00785_));
 sky130_fd_sc_hd__buf_1 _32656_ (.A(_02772_),
    .X(_02810_));
 sky130_fd_sc_hd__a41o_4 _32657_ (.A1(_02692_),
    .A2(_02519_),
    .A3(_02693_),
    .A4(_02694_),
    .B1(_02805_),
    .X(_02811_));
 sky130_fd_sc_hd__o21ai_4 _32658_ (.A1(_20722_),
    .A2(_02810_),
    .B1(_02811_),
    .Y(_00786_));
 sky130_fd_sc_hd__a41o_4 _32659_ (.A1(_02696_),
    .A2(_02521_),
    .A3(_02697_),
    .A4(_02698_),
    .B1(_02767_),
    .X(_02812_));
 sky130_fd_sc_hd__o21ai_4 _32660_ (.A1(_20765_),
    .A2(_02810_),
    .B1(_02812_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand2_4 _32661_ (.A(_02373_),
    .B(_02800_),
    .Y(_02813_));
 sky130_fd_sc_hd__o21ai_4 _32662_ (.A1(_20828_),
    .A2(_02810_),
    .B1(_02813_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand2_4 _32663_ (.A(_02376_),
    .B(_02800_),
    .Y(_02814_));
 sky130_fd_sc_hd__o21ai_4 _32664_ (.A1(_20854_),
    .A2(_02810_),
    .B1(_02814_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand2_4 _32665_ (.A(_02379_),
    .B(_02770_),
    .Y(_02815_));
 sky130_fd_sc_hd__o21ai_4 _32666_ (.A1(_20903_),
    .A2(_02773_),
    .B1(_02815_),
    .Y(_00790_));
 sky130_fd_sc_hd__nand2_4 _32667_ (.A(_02382_),
    .B(_02770_),
    .Y(_02816_));
 sky130_fd_sc_hd__o21ai_4 _32668_ (.A1(_20943_),
    .A2(_02773_),
    .B1(_02816_),
    .Y(_00792_));
 sky130_fd_sc_hd__nand2_4 _32669_ (.A(_02385_),
    .B(_02770_),
    .Y(_02817_));
 sky130_fd_sc_hd__o21ai_4 _32670_ (.A1(_20986_),
    .A2(_02773_),
    .B1(_02817_),
    .Y(_00793_));
 sky130_fd_sc_hd__buf_1 _32671_ (.A(_01767_),
    .X(_02818_));
 sky130_fd_sc_hd__nor4_4 _32672_ (.A(_02705_),
    .B(_01787_),
    .C(_02707_),
    .D(_02818_),
    .Y(_02819_));
 sky130_vsdinv _32673_ (.A(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__buf_1 _32674_ (.A(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__buf_1 _32675_ (.A(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__nor3_4 _32676_ (.A(_02712_),
    .B(_02391_),
    .C(_02393_),
    .Y(_02823_));
 sky130_fd_sc_hd__a21o_4 _32677_ (.A1(\cpuregs[9][0] ),
    .A2(_02822_),
    .B1(_02823_),
    .X(_01345_));
 sky130_fd_sc_hd__and2_4 _32678_ (.A(_02819_),
    .B(_02395_),
    .X(_02824_));
 sky130_fd_sc_hd__a21o_4 _32679_ (.A1(\cpuregs[9][1] ),
    .A2(_02822_),
    .B1(_02824_),
    .X(_01356_));
 sky130_fd_sc_hd__buf_1 _32680_ (.A(_02820_),
    .X(_02825_));
 sky130_fd_sc_hd__buf_1 _32681_ (.A(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__buf_1 _32682_ (.A(_01816_),
    .X(_02827_));
 sky130_fd_sc_hd__nor2_4 _32683_ (.A(_02826_),
    .B(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__a21o_4 _32684_ (.A1(\cpuregs[9][2] ),
    .A2(_02822_),
    .B1(_02828_),
    .X(_01367_));
 sky130_fd_sc_hd__nor2_4 _32685_ (.A(_02826_),
    .B(_02718_),
    .Y(_02829_));
 sky130_fd_sc_hd__a21o_4 _32686_ (.A1(\cpuregs[9][3] ),
    .A2(_02822_),
    .B1(_02829_),
    .X(_01370_));
 sky130_fd_sc_hd__buf_1 _32687_ (.A(_02821_),
    .X(_02830_));
 sky130_fd_sc_hd__buf_1 _32688_ (.A(_23487_),
    .X(_02831_));
 sky130_fd_sc_hd__buf_1 _32689_ (.A(_01836_),
    .X(_02832_));
 sky130_fd_sc_hd__buf_1 _32690_ (.A(_01839_),
    .X(_02833_));
 sky130_fd_sc_hd__buf_1 _32691_ (.A(_01842_),
    .X(_02834_));
 sky130_fd_sc_hd__a41oi_4 _32692_ (.A1(_02831_),
    .A2(_02832_),
    .A3(_02833_),
    .A4(_02834_),
    .B1(_02826_),
    .Y(_02835_));
 sky130_fd_sc_hd__a21o_4 _32693_ (.A1(\cpuregs[9][4] ),
    .A2(_02830_),
    .B1(_02835_),
    .X(_01371_));
 sky130_fd_sc_hd__buf_1 _32694_ (.A(_23494_),
    .X(_02836_));
 sky130_fd_sc_hd__buf_1 _32695_ (.A(_01849_),
    .X(_02837_));
 sky130_fd_sc_hd__buf_1 _32696_ (.A(_01852_),
    .X(_02838_));
 sky130_fd_sc_hd__buf_1 _32697_ (.A(_01856_),
    .X(_02839_));
 sky130_fd_sc_hd__a41oi_4 _32698_ (.A1(_02836_),
    .A2(_02837_),
    .A3(_02838_),
    .A4(_02839_),
    .B1(_02826_),
    .Y(_02840_));
 sky130_fd_sc_hd__a21o_4 _32699_ (.A1(\cpuregs[9][5] ),
    .A2(_02830_),
    .B1(_02840_),
    .X(_01372_));
 sky130_fd_sc_hd__buf_1 _32700_ (.A(_23504_),
    .X(_02841_));
 sky130_fd_sc_hd__buf_1 _32701_ (.A(_01864_),
    .X(_02842_));
 sky130_fd_sc_hd__buf_1 _32702_ (.A(_01867_),
    .X(_02843_));
 sky130_fd_sc_hd__buf_1 _32703_ (.A(_01870_),
    .X(_02844_));
 sky130_fd_sc_hd__buf_1 _32704_ (.A(_02820_),
    .X(_02845_));
 sky130_fd_sc_hd__buf_1 _32705_ (.A(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__a41oi_4 _32706_ (.A1(_02841_),
    .A2(_02842_),
    .A3(_02843_),
    .A4(_02844_),
    .B1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__a21o_4 _32707_ (.A1(\cpuregs[9][6] ),
    .A2(_02830_),
    .B1(_02847_),
    .X(_01373_));
 sky130_fd_sc_hd__buf_1 _32708_ (.A(_23510_),
    .X(_02848_));
 sky130_fd_sc_hd__buf_1 _32709_ (.A(_01880_),
    .X(_02849_));
 sky130_fd_sc_hd__buf_1 _32710_ (.A(_01884_),
    .X(_02850_));
 sky130_fd_sc_hd__buf_1 _32711_ (.A(_01887_),
    .X(_02851_));
 sky130_fd_sc_hd__a41oi_4 _32712_ (.A1(_02848_),
    .A2(_02849_),
    .A3(_02850_),
    .A4(_02851_),
    .B1(_02846_),
    .Y(_02852_));
 sky130_fd_sc_hd__a21o_4 _32713_ (.A1(\cpuregs[9][7] ),
    .A2(_02830_),
    .B1(_02852_),
    .X(_01374_));
 sky130_fd_sc_hd__buf_1 _32714_ (.A(_02821_),
    .X(_02853_));
 sky130_fd_sc_hd__buf_1 _32715_ (.A(_23519_),
    .X(_02854_));
 sky130_fd_sc_hd__buf_1 _32716_ (.A(_01894_),
    .X(_02855_));
 sky130_fd_sc_hd__buf_1 _32717_ (.A(_01897_),
    .X(_02856_));
 sky130_fd_sc_hd__buf_1 _32718_ (.A(_01900_),
    .X(_02857_));
 sky130_fd_sc_hd__a41oi_4 _32719_ (.A1(_02854_),
    .A2(_02855_),
    .A3(_02856_),
    .A4(_02857_),
    .B1(_02846_),
    .Y(_02858_));
 sky130_fd_sc_hd__a21o_4 _32720_ (.A1(\cpuregs[9][8] ),
    .A2(_02853_),
    .B1(_02858_),
    .X(_01375_));
 sky130_fd_sc_hd__buf_1 _32721_ (.A(_23526_),
    .X(_02859_));
 sky130_fd_sc_hd__buf_1 _32722_ (.A(_01907_),
    .X(_02860_));
 sky130_fd_sc_hd__buf_1 _32723_ (.A(_01910_),
    .X(_02861_));
 sky130_fd_sc_hd__buf_1 _32724_ (.A(_01915_),
    .X(_02862_));
 sky130_fd_sc_hd__a41oi_4 _32725_ (.A1(_02859_),
    .A2(_02860_),
    .A3(_02861_),
    .A4(_02862_),
    .B1(_02846_),
    .Y(_02863_));
 sky130_fd_sc_hd__a21o_4 _32726_ (.A1(\cpuregs[9][9] ),
    .A2(_02853_),
    .B1(_02863_),
    .X(_01376_));
 sky130_fd_sc_hd__buf_1 _32727_ (.A(_23536_),
    .X(_02864_));
 sky130_fd_sc_hd__buf_1 _32728_ (.A(_01922_),
    .X(_02865_));
 sky130_fd_sc_hd__buf_1 _32729_ (.A(_01925_),
    .X(_02866_));
 sky130_fd_sc_hd__buf_1 _32730_ (.A(_01928_),
    .X(_02867_));
 sky130_fd_sc_hd__buf_1 _32731_ (.A(_02845_),
    .X(_02868_));
 sky130_fd_sc_hd__a41oi_4 _32732_ (.A1(_02864_),
    .A2(_02865_),
    .A3(_02866_),
    .A4(_02867_),
    .B1(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__a21o_4 _32733_ (.A1(\cpuregs[9][10] ),
    .A2(_02853_),
    .B1(_02869_),
    .X(_01346_));
 sky130_fd_sc_hd__buf_1 _32734_ (.A(_23542_),
    .X(_02870_));
 sky130_fd_sc_hd__buf_1 _32735_ (.A(_01937_),
    .X(_02871_));
 sky130_fd_sc_hd__buf_1 _32736_ (.A(_01941_),
    .X(_02872_));
 sky130_fd_sc_hd__buf_1 _32737_ (.A(_01944_),
    .X(_02873_));
 sky130_fd_sc_hd__a41oi_4 _32738_ (.A1(_02870_),
    .A2(_02871_),
    .A3(_02872_),
    .A4(_02873_),
    .B1(_02868_),
    .Y(_02874_));
 sky130_fd_sc_hd__a21o_4 _32739_ (.A1(\cpuregs[9][11] ),
    .A2(_02853_),
    .B1(_02874_),
    .X(_01347_));
 sky130_fd_sc_hd__buf_1 _32740_ (.A(_02820_),
    .X(_02875_));
 sky130_fd_sc_hd__buf_1 _32741_ (.A(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__buf_1 _32742_ (.A(_23550_),
    .X(_02877_));
 sky130_fd_sc_hd__buf_1 _32743_ (.A(_01952_),
    .X(_02878_));
 sky130_fd_sc_hd__buf_1 _32744_ (.A(_01955_),
    .X(_02879_));
 sky130_fd_sc_hd__buf_1 _32745_ (.A(_01958_),
    .X(_02880_));
 sky130_fd_sc_hd__a41oi_4 _32746_ (.A1(_02877_),
    .A2(_02878_),
    .A3(_02879_),
    .A4(_02880_),
    .B1(_02868_),
    .Y(_02881_));
 sky130_fd_sc_hd__a21o_4 _32747_ (.A1(\cpuregs[9][12] ),
    .A2(_02876_),
    .B1(_02881_),
    .X(_01348_));
 sky130_fd_sc_hd__buf_1 _32748_ (.A(_23557_),
    .X(_02882_));
 sky130_fd_sc_hd__buf_1 _32749_ (.A(_01966_),
    .X(_02883_));
 sky130_fd_sc_hd__buf_1 _32750_ (.A(_01969_),
    .X(_02884_));
 sky130_fd_sc_hd__buf_1 _32751_ (.A(_01973_),
    .X(_02885_));
 sky130_fd_sc_hd__a41oi_4 _32752_ (.A1(_02882_),
    .A2(_02883_),
    .A3(_02884_),
    .A4(_02885_),
    .B1(_02868_),
    .Y(_02886_));
 sky130_fd_sc_hd__a21o_4 _32753_ (.A1(\cpuregs[9][13] ),
    .A2(_02876_),
    .B1(_02886_),
    .X(_01349_));
 sky130_fd_sc_hd__buf_1 _32754_ (.A(_23567_),
    .X(_02887_));
 sky130_fd_sc_hd__buf_1 _32755_ (.A(_01982_),
    .X(_02888_));
 sky130_fd_sc_hd__buf_1 _32756_ (.A(_01985_),
    .X(_02889_));
 sky130_fd_sc_hd__buf_1 _32757_ (.A(_01988_),
    .X(_02890_));
 sky130_fd_sc_hd__buf_1 _32758_ (.A(_02845_),
    .X(_02891_));
 sky130_fd_sc_hd__a41oi_4 _32759_ (.A1(_02887_),
    .A2(_02888_),
    .A3(_02889_),
    .A4(_02890_),
    .B1(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__a21o_4 _32760_ (.A1(\cpuregs[9][14] ),
    .A2(_02876_),
    .B1(_02892_),
    .X(_01350_));
 sky130_fd_sc_hd__buf_1 _32761_ (.A(_23573_),
    .X(_02893_));
 sky130_fd_sc_hd__buf_1 _32762_ (.A(_01998_),
    .X(_02894_));
 sky130_fd_sc_hd__buf_1 _32763_ (.A(_02002_),
    .X(_02895_));
 sky130_fd_sc_hd__buf_1 _32764_ (.A(_02005_),
    .X(_02896_));
 sky130_fd_sc_hd__a41oi_4 _32765_ (.A1(_02893_),
    .A2(_02894_),
    .A3(_02895_),
    .A4(_02896_),
    .B1(_02891_),
    .Y(_02897_));
 sky130_fd_sc_hd__a21o_4 _32766_ (.A1(\cpuregs[9][15] ),
    .A2(_02876_),
    .B1(_02897_),
    .X(_01351_));
 sky130_fd_sc_hd__buf_1 _32767_ (.A(_02875_),
    .X(_02898_));
 sky130_fd_sc_hd__buf_1 _32768_ (.A(_23582_),
    .X(_02899_));
 sky130_fd_sc_hd__buf_1 _32769_ (.A(_02015_),
    .X(_02900_));
 sky130_fd_sc_hd__buf_1 _32770_ (.A(_02018_),
    .X(_02901_));
 sky130_fd_sc_hd__buf_1 _32771_ (.A(_02021_),
    .X(_02902_));
 sky130_fd_sc_hd__a41oi_4 _32772_ (.A1(_02899_),
    .A2(_02900_),
    .A3(_02901_),
    .A4(_02902_),
    .B1(_02891_),
    .Y(_02903_));
 sky130_fd_sc_hd__a21o_4 _32773_ (.A1(\cpuregs[9][16] ),
    .A2(_02898_),
    .B1(_02903_),
    .X(_01352_));
 sky130_fd_sc_hd__buf_1 _32774_ (.A(_23590_),
    .X(_02904_));
 sky130_fd_sc_hd__buf_1 _32775_ (.A(_02030_),
    .X(_02905_));
 sky130_fd_sc_hd__buf_1 _32776_ (.A(_02033_),
    .X(_02906_));
 sky130_fd_sc_hd__buf_1 _32777_ (.A(_02037_),
    .X(_02907_));
 sky130_fd_sc_hd__a41oi_4 _32778_ (.A1(_02904_),
    .A2(_02905_),
    .A3(_02906_),
    .A4(_02907_),
    .B1(_02891_),
    .Y(_02908_));
 sky130_fd_sc_hd__a21o_4 _32779_ (.A1(\cpuregs[9][17] ),
    .A2(_02898_),
    .B1(_02908_),
    .X(_01353_));
 sky130_fd_sc_hd__buf_1 _32780_ (.A(_23598_),
    .X(_02909_));
 sky130_fd_sc_hd__buf_1 _32781_ (.A(_02044_),
    .X(_02910_));
 sky130_fd_sc_hd__buf_1 _32782_ (.A(_02048_),
    .X(_02911_));
 sky130_fd_sc_hd__buf_1 _32783_ (.A(_02051_),
    .X(_02912_));
 sky130_fd_sc_hd__buf_1 _32784_ (.A(_02825_),
    .X(_02913_));
 sky130_fd_sc_hd__a41oi_4 _32785_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_02911_),
    .A4(_02912_),
    .B1(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__a21o_4 _32786_ (.A1(\cpuregs[9][18] ),
    .A2(_02898_),
    .B1(_02914_),
    .X(_01354_));
 sky130_fd_sc_hd__buf_1 _32787_ (.A(_23605_),
    .X(_02915_));
 sky130_fd_sc_hd__buf_1 _32788_ (.A(_02060_),
    .X(_02916_));
 sky130_fd_sc_hd__buf_1 _32789_ (.A(_02063_),
    .X(_02917_));
 sky130_fd_sc_hd__buf_1 _32790_ (.A(_02066_),
    .X(_02918_));
 sky130_fd_sc_hd__a41oi_4 _32791_ (.A1(_02915_),
    .A2(_02916_),
    .A3(_02917_),
    .A4(_02918_),
    .B1(_02913_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21o_4 _32792_ (.A1(\cpuregs[9][19] ),
    .A2(_02898_),
    .B1(_02919_),
    .X(_01355_));
 sky130_fd_sc_hd__buf_1 _32793_ (.A(_02875_),
    .X(_02920_));
 sky130_fd_sc_hd__buf_1 _32794_ (.A(_23613_),
    .X(_02921_));
 sky130_fd_sc_hd__buf_1 _32795_ (.A(_02076_),
    .X(_02922_));
 sky130_fd_sc_hd__buf_1 _32796_ (.A(_02080_),
    .X(_02923_));
 sky130_fd_sc_hd__buf_1 _32797_ (.A(_02083_),
    .X(_02924_));
 sky130_fd_sc_hd__a41oi_4 _32798_ (.A1(_02921_),
    .A2(_02922_),
    .A3(_02923_),
    .A4(_02924_),
    .B1(_02913_),
    .Y(_02925_));
 sky130_fd_sc_hd__a21o_4 _32799_ (.A1(\cpuregs[9][20] ),
    .A2(_02920_),
    .B1(_02925_),
    .X(_01357_));
 sky130_fd_sc_hd__buf_1 _32800_ (.A(_23620_),
    .X(_02926_));
 sky130_fd_sc_hd__buf_1 _32801_ (.A(_02091_),
    .X(_02927_));
 sky130_fd_sc_hd__buf_1 _32802_ (.A(_02094_),
    .X(_02928_));
 sky130_fd_sc_hd__buf_1 _32803_ (.A(_02097_),
    .X(_02929_));
 sky130_fd_sc_hd__a41oi_4 _32804_ (.A1(_02926_),
    .A2(_02927_),
    .A3(_02928_),
    .A4(_02929_),
    .B1(_02913_),
    .Y(_02930_));
 sky130_fd_sc_hd__a21o_4 _32805_ (.A1(\cpuregs[9][21] ),
    .A2(_02920_),
    .B1(_02930_),
    .X(_01358_));
 sky130_fd_sc_hd__buf_1 _32806_ (.A(_23627_),
    .X(_02931_));
 sky130_fd_sc_hd__buf_1 _32807_ (.A(_02105_),
    .X(_02932_));
 sky130_fd_sc_hd__buf_1 _32808_ (.A(_02108_),
    .X(_02933_));
 sky130_fd_sc_hd__buf_1 _32809_ (.A(_02112_),
    .X(_02934_));
 sky130_fd_sc_hd__buf_1 _32810_ (.A(_02825_),
    .X(_02935_));
 sky130_fd_sc_hd__a41oi_4 _32811_ (.A1(_02931_),
    .A2(_02932_),
    .A3(_02933_),
    .A4(_02934_),
    .B1(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__a21o_4 _32812_ (.A1(\cpuregs[9][22] ),
    .A2(_02920_),
    .B1(_02936_),
    .X(_01359_));
 sky130_fd_sc_hd__buf_1 _32813_ (.A(_23633_),
    .X(_02937_));
 sky130_fd_sc_hd__buf_1 _32814_ (.A(_02121_),
    .X(_02938_));
 sky130_fd_sc_hd__buf_1 _32815_ (.A(_02124_),
    .X(_02939_));
 sky130_fd_sc_hd__buf_1 _32816_ (.A(_02128_),
    .X(_02940_));
 sky130_fd_sc_hd__a41oi_4 _32817_ (.A1(_02937_),
    .A2(_02938_),
    .A3(_02939_),
    .A4(_02940_),
    .B1(_02935_),
    .Y(_02941_));
 sky130_fd_sc_hd__a21o_4 _32818_ (.A1(\cpuregs[9][23] ),
    .A2(_02920_),
    .B1(_02941_),
    .X(_01360_));
 sky130_fd_sc_hd__buf_1 _32819_ (.A(_02875_),
    .X(_02942_));
 sky130_fd_sc_hd__buf_1 _32820_ (.A(_23641_),
    .X(_02943_));
 sky130_fd_sc_hd__buf_1 _32821_ (.A(_02138_),
    .X(_02944_));
 sky130_fd_sc_hd__buf_1 _32822_ (.A(_02141_),
    .X(_02945_));
 sky130_fd_sc_hd__buf_1 _32823_ (.A(_02144_),
    .X(_02946_));
 sky130_fd_sc_hd__a41oi_4 _32824_ (.A1(_02943_),
    .A2(_02944_),
    .A3(_02945_),
    .A4(_02946_),
    .B1(_02935_),
    .Y(_02947_));
 sky130_fd_sc_hd__a21o_4 _32825_ (.A1(\cpuregs[9][24] ),
    .A2(_02942_),
    .B1(_02947_),
    .X(_01361_));
 sky130_fd_sc_hd__buf_1 _32826_ (.A(_23648_),
    .X(_02948_));
 sky130_fd_sc_hd__buf_1 _32827_ (.A(_02153_),
    .X(_02949_));
 sky130_fd_sc_hd__buf_1 _32828_ (.A(_02156_),
    .X(_02950_));
 sky130_fd_sc_hd__buf_1 _32829_ (.A(_02159_),
    .X(_02951_));
 sky130_fd_sc_hd__a41oi_4 _32830_ (.A1(_02948_),
    .A2(_02949_),
    .A3(_02950_),
    .A4(_02951_),
    .B1(_02935_),
    .Y(_02952_));
 sky130_fd_sc_hd__a21o_4 _32831_ (.A1(\cpuregs[9][25] ),
    .A2(_02942_),
    .B1(_02952_),
    .X(_01362_));
 sky130_fd_sc_hd__buf_1 _32832_ (.A(_23656_),
    .X(_02953_));
 sky130_fd_sc_hd__buf_1 _32833_ (.A(_02167_),
    .X(_02954_));
 sky130_fd_sc_hd__buf_1 _32834_ (.A(_02170_),
    .X(_02955_));
 sky130_fd_sc_hd__buf_1 _32835_ (.A(_02173_),
    .X(_02956_));
 sky130_fd_sc_hd__buf_1 _32836_ (.A(_02825_),
    .X(_02957_));
 sky130_fd_sc_hd__a41oi_4 _32837_ (.A1(_02953_),
    .A2(_02954_),
    .A3(_02955_),
    .A4(_02956_),
    .B1(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__a21o_4 _32838_ (.A1(\cpuregs[9][26] ),
    .A2(_02942_),
    .B1(_02958_),
    .X(_01363_));
 sky130_fd_sc_hd__buf_1 _32839_ (.A(_23661_),
    .X(_02959_));
 sky130_fd_sc_hd__buf_1 _32840_ (.A(_02183_),
    .X(_02960_));
 sky130_fd_sc_hd__buf_1 _32841_ (.A(_02186_),
    .X(_02961_));
 sky130_fd_sc_hd__buf_1 _32842_ (.A(_02189_),
    .X(_02962_));
 sky130_fd_sc_hd__a41oi_4 _32843_ (.A1(_02959_),
    .A2(_02960_),
    .A3(_02961_),
    .A4(_02962_),
    .B1(_02957_),
    .Y(_02963_));
 sky130_fd_sc_hd__a21o_4 _32844_ (.A1(\cpuregs[9][27] ),
    .A2(_02942_),
    .B1(_02963_),
    .X(_01364_));
 sky130_fd_sc_hd__buf_1 _32845_ (.A(_02845_),
    .X(_02964_));
 sky130_fd_sc_hd__and2_4 _32846_ (.A(_02759_),
    .B(_02819_),
    .X(_02965_));
 sky130_fd_sc_hd__a21o_4 _32847_ (.A1(\cpuregs[9][28] ),
    .A2(_02964_),
    .B1(_02965_),
    .X(_01365_));
 sky130_fd_sc_hd__buf_1 _32848_ (.A(_23673_),
    .X(_02966_));
 sky130_fd_sc_hd__buf_1 _32849_ (.A(_02205_),
    .X(_02967_));
 sky130_fd_sc_hd__buf_1 _32850_ (.A(_02208_),
    .X(_02968_));
 sky130_fd_sc_hd__buf_1 _32851_ (.A(_02211_),
    .X(_02969_));
 sky130_fd_sc_hd__a41oi_4 _32852_ (.A1(_02966_),
    .A2(_02967_),
    .A3(_02968_),
    .A4(_02969_),
    .B1(_02957_),
    .Y(_02970_));
 sky130_fd_sc_hd__a21o_4 _32853_ (.A1(\cpuregs[9][29] ),
    .A2(_02964_),
    .B1(_02970_),
    .X(_01366_));
 sky130_fd_sc_hd__buf_1 _32854_ (.A(_23680_),
    .X(_02971_));
 sky130_fd_sc_hd__buf_1 _32855_ (.A(_02218_),
    .X(_02972_));
 sky130_fd_sc_hd__buf_1 _32856_ (.A(_02221_),
    .X(_02973_));
 sky130_fd_sc_hd__buf_1 _32857_ (.A(_02224_),
    .X(_02974_));
 sky130_fd_sc_hd__a41oi_4 _32858_ (.A1(_02971_),
    .A2(_02972_),
    .A3(_02973_),
    .A4(_02974_),
    .B1(_02957_),
    .Y(_02975_));
 sky130_fd_sc_hd__a21o_4 _32859_ (.A1(\cpuregs[9][30] ),
    .A2(_02964_),
    .B1(_02975_),
    .X(_01368_));
 sky130_fd_sc_hd__buf_1 _32860_ (.A(_23685_),
    .X(_02976_));
 sky130_fd_sc_hd__buf_1 _32861_ (.A(_02232_),
    .X(_02977_));
 sky130_fd_sc_hd__buf_1 _32862_ (.A(_02235_),
    .X(_02978_));
 sky130_fd_sc_hd__buf_1 _32863_ (.A(_02238_),
    .X(_02979_));
 sky130_fd_sc_hd__a41oi_4 _32864_ (.A1(_02976_),
    .A2(_02977_),
    .A3(_02978_),
    .A4(_02979_),
    .B1(_02821_),
    .Y(_02980_));
 sky130_fd_sc_hd__a21o_4 _32865_ (.A1(\cpuregs[9][31] ),
    .A2(_02964_),
    .B1(_02980_),
    .X(_01369_));
 sky130_fd_sc_hd__nor2_4 _32866_ (.A(_02712_),
    .B(_02445_),
    .Y(_02981_));
 sky130_vsdinv _32867_ (.A(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__buf_1 _32868_ (.A(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_1 _32869_ (.A(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__nor3_4 _32870_ (.A(_02450_),
    .B(_02712_),
    .C(_01783_),
    .Y(_02985_));
 sky130_fd_sc_hd__a21o_4 _32871_ (.A1(\cpuregs[8][0] ),
    .A2(_02984_),
    .B1(_02985_),
    .X(_01313_));
 sky130_fd_sc_hd__buf_1 _32872_ (.A(_02981_),
    .X(_02986_));
 sky130_fd_sc_hd__buf_1 _32873_ (.A(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__buf_1 _32874_ (.A(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__buf_1 _32875_ (.A(_01802_),
    .X(_02989_));
 sky130_fd_sc_hd__buf_1 _32876_ (.A(_02986_),
    .X(_02990_));
 sky130_fd_sc_hd__nand2_4 _32877_ (.A(_02989_),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__o21ai_4 _32878_ (.A1(_19313_),
    .A2(_02988_),
    .B1(_02991_),
    .Y(_01324_));
 sky130_fd_sc_hd__buf_1 _32879_ (.A(_02983_),
    .X(_02992_));
 sky130_fd_sc_hd__a41oi_4 _32880_ (.A1(_02458_),
    .A2(_02460_),
    .A3(_02462_),
    .A4(_02464_),
    .B1(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__a21o_4 _32881_ (.A1(\cpuregs[8][2] ),
    .A2(_02984_),
    .B1(_02993_),
    .X(_01335_));
 sky130_fd_sc_hd__nor2_4 _32882_ (.A(_02984_),
    .B(_02718_),
    .Y(_02994_));
 sky130_fd_sc_hd__a21o_4 _32883_ (.A1(\cpuregs[8][3] ),
    .A2(_02984_),
    .B1(_02994_),
    .X(_01338_));
 sky130_fd_sc_hd__a41o_4 _32884_ (.A1(_02601_),
    .A2(_02468_),
    .A3(_02602_),
    .A4(_02603_),
    .B1(_02992_),
    .X(_02995_));
 sky130_fd_sc_hd__o21ai_4 _32885_ (.A1(_19589_),
    .A2(_02988_),
    .B1(_02995_),
    .Y(_01339_));
 sky130_fd_sc_hd__a41o_4 _32886_ (.A1(_02608_),
    .A2(_02470_),
    .A3(_02609_),
    .A4(_02610_),
    .B1(_02992_),
    .X(_02996_));
 sky130_fd_sc_hd__o21ai_4 _32887_ (.A1(_19663_),
    .A2(_02988_),
    .B1(_02996_),
    .Y(_01340_));
 sky130_fd_sc_hd__a41o_4 _32888_ (.A1(_02612_),
    .A2(_02472_),
    .A3(_02613_),
    .A4(_02614_),
    .B1(_02992_),
    .X(_02997_));
 sky130_fd_sc_hd__o21ai_4 _32889_ (.A1(_19708_),
    .A2(_02988_),
    .B1(_02997_),
    .Y(_01341_));
 sky130_fd_sc_hd__buf_1 _32890_ (.A(_02987_),
    .X(_02998_));
 sky130_fd_sc_hd__buf_1 _32891_ (.A(_02982_),
    .X(_02999_));
 sky130_fd_sc_hd__buf_1 _32892_ (.A(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__a41o_4 _32893_ (.A1(_02616_),
    .A2(_02475_),
    .A3(_02617_),
    .A4(_02618_),
    .B1(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__o21ai_4 _32894_ (.A1(_19762_),
    .A2(_02998_),
    .B1(_03001_),
    .Y(_01342_));
 sky130_fd_sc_hd__a41o_4 _32895_ (.A1(_02620_),
    .A2(_02479_),
    .A3(_02621_),
    .A4(_02622_),
    .B1(_03000_),
    .X(_03002_));
 sky130_fd_sc_hd__o21ai_4 _32896_ (.A1(_19818_),
    .A2(_02998_),
    .B1(_03002_),
    .Y(_01343_));
 sky130_fd_sc_hd__a41o_4 _32897_ (.A1(_02626_),
    .A2(_02481_),
    .A3(_02627_),
    .A4(_02628_),
    .B1(_03000_),
    .X(_03003_));
 sky130_fd_sc_hd__o21ai_4 _32898_ (.A1(_19877_),
    .A2(_02998_),
    .B1(_03003_),
    .Y(_01344_));
 sky130_fd_sc_hd__a41o_4 _32899_ (.A1(_02630_),
    .A2(_02483_),
    .A3(_02631_),
    .A4(_02632_),
    .B1(_03000_),
    .X(_03004_));
 sky130_fd_sc_hd__o21ai_4 _32900_ (.A1(_19957_),
    .A2(_02998_),
    .B1(_03004_),
    .Y(_01314_));
 sky130_fd_sc_hd__buf_1 _32901_ (.A(_02987_),
    .X(_03005_));
 sky130_fd_sc_hd__buf_1 _32902_ (.A(_02999_),
    .X(_03006_));
 sky130_fd_sc_hd__a41o_4 _32903_ (.A1(_02634_),
    .A2(_02486_),
    .A3(_02635_),
    .A4(_02636_),
    .B1(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__o21ai_4 _32904_ (.A1(_19995_),
    .A2(_03005_),
    .B1(_03007_),
    .Y(_01315_));
 sky130_fd_sc_hd__a41o_4 _32905_ (.A1(_02638_),
    .A2(_02489_),
    .A3(_02639_),
    .A4(_02640_),
    .B1(_03006_),
    .X(_03008_));
 sky130_fd_sc_hd__o21ai_4 _32906_ (.A1(_20069_),
    .A2(_03005_),
    .B1(_03008_),
    .Y(_01316_));
 sky130_fd_sc_hd__a41o_4 _32907_ (.A1(_02644_),
    .A2(_02491_),
    .A3(_02645_),
    .A4(_02646_),
    .B1(_03006_),
    .X(_03009_));
 sky130_fd_sc_hd__o21ai_4 _32908_ (.A1(_20125_),
    .A2(_03005_),
    .B1(_03009_),
    .Y(_01317_));
 sky130_fd_sc_hd__a41o_4 _32909_ (.A1(_02648_),
    .A2(_02493_),
    .A3(_02649_),
    .A4(_02650_),
    .B1(_03006_),
    .X(_03010_));
 sky130_fd_sc_hd__o21ai_4 _32910_ (.A1(_20189_),
    .A2(_03005_),
    .B1(_03010_),
    .Y(_01318_));
 sky130_fd_sc_hd__buf_1 _32911_ (.A(_02986_),
    .X(_03011_));
 sky130_fd_sc_hd__buf_1 _32912_ (.A(_03011_),
    .X(_03012_));
 sky130_fd_sc_hd__buf_1 _32913_ (.A(_02999_),
    .X(_03013_));
 sky130_fd_sc_hd__a41o_4 _32914_ (.A1(_02652_),
    .A2(_02497_),
    .A3(_02653_),
    .A4(_02654_),
    .B1(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__o21ai_4 _32915_ (.A1(_20243_),
    .A2(_03012_),
    .B1(_03014_),
    .Y(_01319_));
 sky130_fd_sc_hd__a41o_4 _32916_ (.A1(_02656_),
    .A2(_02500_),
    .A3(_02657_),
    .A4(_02658_),
    .B1(_03013_),
    .X(_03015_));
 sky130_fd_sc_hd__o21ai_4 _32917_ (.A1(_20288_),
    .A2(_03012_),
    .B1(_03015_),
    .Y(_01320_));
 sky130_fd_sc_hd__a41o_4 _32918_ (.A1(_02662_),
    .A2(_02502_),
    .A3(_02663_),
    .A4(_02664_),
    .B1(_03013_),
    .X(_03016_));
 sky130_fd_sc_hd__o21ai_4 _32919_ (.A1(_20343_),
    .A2(_03012_),
    .B1(_03016_),
    .Y(_01321_));
 sky130_fd_sc_hd__buf_1 _32920_ (.A(_02334_),
    .X(_03017_));
 sky130_fd_sc_hd__nand2_4 _32921_ (.A(_03017_),
    .B(_02990_),
    .Y(_03018_));
 sky130_fd_sc_hd__o21ai_4 _32922_ (.A1(_20398_),
    .A2(_03012_),
    .B1(_03018_),
    .Y(_01322_));
 sky130_fd_sc_hd__buf_1 _32923_ (.A(_03011_),
    .X(_03019_));
 sky130_fd_sc_hd__a41o_4 _32924_ (.A1(_02668_),
    .A2(_02506_),
    .A3(_02669_),
    .A4(_02670_),
    .B1(_03013_),
    .X(_03020_));
 sky130_fd_sc_hd__o21ai_4 _32925_ (.A1(_20447_),
    .A2(_03019_),
    .B1(_03020_),
    .Y(_01323_));
 sky130_fd_sc_hd__buf_1 _32926_ (.A(_02999_),
    .X(_03021_));
 sky130_fd_sc_hd__a41o_4 _32927_ (.A1(_02672_),
    .A2(_02508_),
    .A3(_02673_),
    .A4(_02674_),
    .B1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__o21ai_4 _32928_ (.A1(_20489_),
    .A2(_03019_),
    .B1(_03022_),
    .Y(_01325_));
 sky130_fd_sc_hd__a41o_4 _32929_ (.A1(_02677_),
    .A2(_02511_),
    .A3(_02678_),
    .A4(_02679_),
    .B1(_03021_),
    .X(_03023_));
 sky130_fd_sc_hd__o21ai_4 _32930_ (.A1(_20543_),
    .A2(_03019_),
    .B1(_03023_),
    .Y(_01326_));
 sky130_fd_sc_hd__buf_1 _32931_ (.A(_02352_),
    .X(_03024_));
 sky130_fd_sc_hd__nand2_4 _32932_ (.A(_03024_),
    .B(_02990_),
    .Y(_03025_));
 sky130_fd_sc_hd__o21ai_4 _32933_ (.A1(_20599_),
    .A2(_03019_),
    .B1(_03025_),
    .Y(_01327_));
 sky130_fd_sc_hd__buf_1 _32934_ (.A(_03011_),
    .X(_03026_));
 sky130_fd_sc_hd__a41o_4 _32935_ (.A1(_02683_),
    .A2(_02515_),
    .A3(_02684_),
    .A4(_02685_),
    .B1(_03021_),
    .X(_03027_));
 sky130_fd_sc_hd__o21ai_4 _32936_ (.A1(_20626_),
    .A2(_03026_),
    .B1(_03027_),
    .Y(_01328_));
 sky130_fd_sc_hd__a41o_4 _32937_ (.A1(_02687_),
    .A2(_02517_),
    .A3(_02688_),
    .A4(_02689_),
    .B1(_03021_),
    .X(_03028_));
 sky130_fd_sc_hd__o21ai_4 _32938_ (.A1(_20671_),
    .A2(_03026_),
    .B1(_03028_),
    .Y(_01329_));
 sky130_fd_sc_hd__a41o_4 _32939_ (.A1(_02692_),
    .A2(_02519_),
    .A3(_02693_),
    .A4(_02694_),
    .B1(_02983_),
    .X(_03029_));
 sky130_fd_sc_hd__o21ai_4 _32940_ (.A1(_20719_),
    .A2(_03026_),
    .B1(_03029_),
    .Y(_01330_));
 sky130_fd_sc_hd__a41o_4 _32941_ (.A1(_02696_),
    .A2(_02521_),
    .A3(_02697_),
    .A4(_02698_),
    .B1(_02983_),
    .X(_03030_));
 sky130_fd_sc_hd__o21ai_4 _32942_ (.A1(_20762_),
    .A2(_03026_),
    .B1(_03030_),
    .Y(_01331_));
 sky130_fd_sc_hd__buf_1 _32943_ (.A(_03011_),
    .X(_03031_));
 sky130_fd_sc_hd__buf_1 _32944_ (.A(_02372_),
    .X(_03032_));
 sky130_fd_sc_hd__buf_1 _32945_ (.A(_02986_),
    .X(_03033_));
 sky130_fd_sc_hd__nand2_4 _32946_ (.A(_03032_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__o21ai_4 _32947_ (.A1(_20825_),
    .A2(_03031_),
    .B1(_03034_),
    .Y(_01332_));
 sky130_fd_sc_hd__buf_1 _32948_ (.A(_02197_),
    .X(_03035_));
 sky130_fd_sc_hd__nand2_4 _32949_ (.A(_03035_),
    .B(_03033_),
    .Y(_03036_));
 sky130_fd_sc_hd__o21ai_4 _32950_ (.A1(_20851_),
    .A2(_03031_),
    .B1(_03036_),
    .Y(_01333_));
 sky130_fd_sc_hd__buf_1 _32951_ (.A(_02378_),
    .X(_03037_));
 sky130_fd_sc_hd__nand2_4 _32952_ (.A(_03037_),
    .B(_03033_),
    .Y(_03038_));
 sky130_fd_sc_hd__o21ai_4 _32953_ (.A1(_20900_),
    .A2(_03031_),
    .B1(_03038_),
    .Y(_01334_));
 sky130_fd_sc_hd__buf_1 _32954_ (.A(_02381_),
    .X(_03039_));
 sky130_fd_sc_hd__nand2_4 _32955_ (.A(_03039_),
    .B(_03033_),
    .Y(_03040_));
 sky130_fd_sc_hd__o21ai_4 _32956_ (.A1(_20940_),
    .A2(_03031_),
    .B1(_03040_),
    .Y(_01336_));
 sky130_fd_sc_hd__buf_1 _32957_ (.A(_02384_),
    .X(_03041_));
 sky130_fd_sc_hd__nand2_4 _32958_ (.A(_03041_),
    .B(_02987_),
    .Y(_03042_));
 sky130_fd_sc_hd__o21ai_4 _32959_ (.A1(_20983_),
    .A2(_02990_),
    .B1(_03042_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor3_4 _32960_ (.A(_19094_),
    .B(_19098_),
    .C(_19090_),
    .Y(_03043_));
 sky130_vsdinv _32961_ (.A(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__nor4_4 _32962_ (.A(_02705_),
    .B(_19086_),
    .C(_03044_),
    .D(_02818_),
    .Y(_03045_));
 sky130_vsdinv _32963_ (.A(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__buf_1 _32964_ (.A(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__buf_1 _32965_ (.A(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__buf_1 _32966_ (.A(_03044_),
    .X(_03049_));
 sky130_fd_sc_hd__nor3_4 _32967_ (.A(_03049_),
    .B(_02248_),
    .C(_01790_),
    .Y(_03050_));
 sky130_fd_sc_hd__a21o_4 _32968_ (.A1(\cpuregs[7][0] ),
    .A2(_03048_),
    .B1(_03050_),
    .X(_01281_));
 sky130_fd_sc_hd__and2_4 _32969_ (.A(_03045_),
    .B(_02253_),
    .X(_03051_));
 sky130_fd_sc_hd__a21o_4 _32970_ (.A1(\cpuregs[7][1] ),
    .A2(_03048_),
    .B1(_03051_),
    .X(_01292_));
 sky130_fd_sc_hd__buf_1 _32971_ (.A(_03046_),
    .X(_03052_));
 sky130_fd_sc_hd__buf_1 _32972_ (.A(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__nor2_4 _32973_ (.A(_03053_),
    .B(_02827_),
    .Y(_03054_));
 sky130_fd_sc_hd__a21o_4 _32974_ (.A1(\cpuregs[7][2] ),
    .A2(_03048_),
    .B1(_03054_),
    .X(_01303_));
 sky130_fd_sc_hd__nor2_4 _32975_ (.A(_03053_),
    .B(_02718_),
    .Y(_03055_));
 sky130_fd_sc_hd__a21o_4 _32976_ (.A1(\cpuregs[7][3] ),
    .A2(_03048_),
    .B1(_03055_),
    .X(_01306_));
 sky130_fd_sc_hd__buf_1 _32977_ (.A(_03047_),
    .X(_03056_));
 sky130_fd_sc_hd__a41oi_4 _32978_ (.A1(_02831_),
    .A2(_02832_),
    .A3(_02833_),
    .A4(_02834_),
    .B1(_03053_),
    .Y(_03057_));
 sky130_fd_sc_hd__a21o_4 _32979_ (.A1(\cpuregs[7][4] ),
    .A2(_03056_),
    .B1(_03057_),
    .X(_01307_));
 sky130_fd_sc_hd__a41oi_4 _32980_ (.A1(_02836_),
    .A2(_02837_),
    .A3(_02838_),
    .A4(_02839_),
    .B1(_03053_),
    .Y(_03058_));
 sky130_fd_sc_hd__a21o_4 _32981_ (.A1(\cpuregs[7][5] ),
    .A2(_03056_),
    .B1(_03058_),
    .X(_01308_));
 sky130_fd_sc_hd__buf_1 _32982_ (.A(_03046_),
    .X(_03059_));
 sky130_fd_sc_hd__buf_1 _32983_ (.A(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__a41oi_4 _32984_ (.A1(_02841_),
    .A2(_02842_),
    .A3(_02843_),
    .A4(_02844_),
    .B1(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__a21o_4 _32985_ (.A1(\cpuregs[7][6] ),
    .A2(_03056_),
    .B1(_03061_),
    .X(_01309_));
 sky130_fd_sc_hd__a41oi_4 _32986_ (.A1(_02848_),
    .A2(_02849_),
    .A3(_02850_),
    .A4(_02851_),
    .B1(_03060_),
    .Y(_03062_));
 sky130_fd_sc_hd__a21o_4 _32987_ (.A1(\cpuregs[7][7] ),
    .A2(_03056_),
    .B1(_03062_),
    .X(_01310_));
 sky130_fd_sc_hd__buf_1 _32988_ (.A(_03047_),
    .X(_03063_));
 sky130_fd_sc_hd__a41oi_4 _32989_ (.A1(_02854_),
    .A2(_02855_),
    .A3(_02856_),
    .A4(_02857_),
    .B1(_03060_),
    .Y(_03064_));
 sky130_fd_sc_hd__a21o_4 _32990_ (.A1(\cpuregs[7][8] ),
    .A2(_03063_),
    .B1(_03064_),
    .X(_01311_));
 sky130_fd_sc_hd__a41oi_4 _32991_ (.A1(_02859_),
    .A2(_02860_),
    .A3(_02861_),
    .A4(_02862_),
    .B1(_03060_),
    .Y(_03065_));
 sky130_fd_sc_hd__a21o_4 _32992_ (.A1(\cpuregs[7][9] ),
    .A2(_03063_),
    .B1(_03065_),
    .X(_01312_));
 sky130_fd_sc_hd__buf_1 _32993_ (.A(_03059_),
    .X(_03066_));
 sky130_fd_sc_hd__a41oi_4 _32994_ (.A1(_02864_),
    .A2(_02865_),
    .A3(_02866_),
    .A4(_02867_),
    .B1(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__a21o_4 _32995_ (.A1(\cpuregs[7][10] ),
    .A2(_03063_),
    .B1(_03067_),
    .X(_01282_));
 sky130_fd_sc_hd__a41oi_4 _32996_ (.A1(_02870_),
    .A2(_02871_),
    .A3(_02872_),
    .A4(_02873_),
    .B1(_03066_),
    .Y(_03068_));
 sky130_fd_sc_hd__a21o_4 _32997_ (.A1(\cpuregs[7][11] ),
    .A2(_03063_),
    .B1(_03068_),
    .X(_01283_));
 sky130_fd_sc_hd__buf_1 _32998_ (.A(_03046_),
    .X(_03069_));
 sky130_fd_sc_hd__buf_1 _32999_ (.A(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__a41oi_4 _33000_ (.A1(_02877_),
    .A2(_02878_),
    .A3(_02879_),
    .A4(_02880_),
    .B1(_03066_),
    .Y(_03071_));
 sky130_fd_sc_hd__a21o_4 _33001_ (.A1(\cpuregs[7][12] ),
    .A2(_03070_),
    .B1(_03071_),
    .X(_01284_));
 sky130_fd_sc_hd__a41oi_4 _33002_ (.A1(_02882_),
    .A2(_02883_),
    .A3(_02884_),
    .A4(_02885_),
    .B1(_03066_),
    .Y(_03072_));
 sky130_fd_sc_hd__a21o_4 _33003_ (.A1(\cpuregs[7][13] ),
    .A2(_03070_),
    .B1(_03072_),
    .X(_01285_));
 sky130_fd_sc_hd__buf_1 _33004_ (.A(_03059_),
    .X(_03073_));
 sky130_fd_sc_hd__a41oi_4 _33005_ (.A1(_02887_),
    .A2(_02888_),
    .A3(_02889_),
    .A4(_02890_),
    .B1(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__a21o_4 _33006_ (.A1(\cpuregs[7][14] ),
    .A2(_03070_),
    .B1(_03074_),
    .X(_01286_));
 sky130_fd_sc_hd__a41oi_4 _33007_ (.A1(_02893_),
    .A2(_02894_),
    .A3(_02895_),
    .A4(_02896_),
    .B1(_03073_),
    .Y(_03075_));
 sky130_fd_sc_hd__a21o_4 _33008_ (.A1(\cpuregs[7][15] ),
    .A2(_03070_),
    .B1(_03075_),
    .X(_01287_));
 sky130_fd_sc_hd__buf_1 _33009_ (.A(_03069_),
    .X(_03076_));
 sky130_fd_sc_hd__a41oi_4 _33010_ (.A1(_02899_),
    .A2(_02900_),
    .A3(_02901_),
    .A4(_02902_),
    .B1(_03073_),
    .Y(_03077_));
 sky130_fd_sc_hd__a21o_4 _33011_ (.A1(\cpuregs[7][16] ),
    .A2(_03076_),
    .B1(_03077_),
    .X(_01288_));
 sky130_fd_sc_hd__a41oi_4 _33012_ (.A1(_02904_),
    .A2(_02905_),
    .A3(_02906_),
    .A4(_02907_),
    .B1(_03073_),
    .Y(_03078_));
 sky130_fd_sc_hd__a21o_4 _33013_ (.A1(\cpuregs[7][17] ),
    .A2(_03076_),
    .B1(_03078_),
    .X(_01289_));
 sky130_fd_sc_hd__buf_1 _33014_ (.A(_03052_),
    .X(_03079_));
 sky130_fd_sc_hd__a41oi_4 _33015_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_02911_),
    .A4(_02912_),
    .B1(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__a21o_4 _33016_ (.A1(\cpuregs[7][18] ),
    .A2(_03076_),
    .B1(_03080_),
    .X(_01290_));
 sky130_fd_sc_hd__a41oi_4 _33017_ (.A1(_02915_),
    .A2(_02916_),
    .A3(_02917_),
    .A4(_02918_),
    .B1(_03079_),
    .Y(_03081_));
 sky130_fd_sc_hd__a21o_4 _33018_ (.A1(\cpuregs[7][19] ),
    .A2(_03076_),
    .B1(_03081_),
    .X(_01291_));
 sky130_fd_sc_hd__buf_1 _33019_ (.A(_03069_),
    .X(_03082_));
 sky130_fd_sc_hd__a41oi_4 _33020_ (.A1(_02921_),
    .A2(_02922_),
    .A3(_02923_),
    .A4(_02924_),
    .B1(_03079_),
    .Y(_03083_));
 sky130_fd_sc_hd__a21o_4 _33021_ (.A1(\cpuregs[7][20] ),
    .A2(_03082_),
    .B1(_03083_),
    .X(_01293_));
 sky130_fd_sc_hd__a41oi_4 _33022_ (.A1(_02926_),
    .A2(_02927_),
    .A3(_02928_),
    .A4(_02929_),
    .B1(_03079_),
    .Y(_03084_));
 sky130_fd_sc_hd__a21o_4 _33023_ (.A1(\cpuregs[7][21] ),
    .A2(_03082_),
    .B1(_03084_),
    .X(_01294_));
 sky130_fd_sc_hd__buf_1 _33024_ (.A(_03052_),
    .X(_03085_));
 sky130_fd_sc_hd__a41oi_4 _33025_ (.A1(_02931_),
    .A2(_02932_),
    .A3(_02933_),
    .A4(_02934_),
    .B1(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__a21o_4 _33026_ (.A1(\cpuregs[7][22] ),
    .A2(_03082_),
    .B1(_03086_),
    .X(_01295_));
 sky130_fd_sc_hd__a41oi_4 _33027_ (.A1(_02937_),
    .A2(_02938_),
    .A3(_02939_),
    .A4(_02940_),
    .B1(_03085_),
    .Y(_03087_));
 sky130_fd_sc_hd__a21o_4 _33028_ (.A1(\cpuregs[7][23] ),
    .A2(_03082_),
    .B1(_03087_),
    .X(_01296_));
 sky130_fd_sc_hd__buf_1 _33029_ (.A(_03069_),
    .X(_03088_));
 sky130_fd_sc_hd__a41oi_4 _33030_ (.A1(_02943_),
    .A2(_02944_),
    .A3(_02945_),
    .A4(_02946_),
    .B1(_03085_),
    .Y(_03089_));
 sky130_fd_sc_hd__a21o_4 _33031_ (.A1(\cpuregs[7][24] ),
    .A2(_03088_),
    .B1(_03089_),
    .X(_01297_));
 sky130_fd_sc_hd__a41oi_4 _33032_ (.A1(_02948_),
    .A2(_02949_),
    .A3(_02950_),
    .A4(_02951_),
    .B1(_03085_),
    .Y(_03090_));
 sky130_fd_sc_hd__a21o_4 _33033_ (.A1(\cpuregs[7][25] ),
    .A2(_03088_),
    .B1(_03090_),
    .X(_01298_));
 sky130_fd_sc_hd__buf_1 _33034_ (.A(_03052_),
    .X(_03091_));
 sky130_fd_sc_hd__a41oi_4 _33035_ (.A1(_02953_),
    .A2(_02954_),
    .A3(_02955_),
    .A4(_02956_),
    .B1(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__a21o_4 _33036_ (.A1(\cpuregs[7][26] ),
    .A2(_03088_),
    .B1(_03092_),
    .X(_01299_));
 sky130_fd_sc_hd__a41oi_4 _33037_ (.A1(_02959_),
    .A2(_02960_),
    .A3(_02961_),
    .A4(_02962_),
    .B1(_03091_),
    .Y(_03093_));
 sky130_fd_sc_hd__a21o_4 _33038_ (.A1(\cpuregs[7][27] ),
    .A2(_03088_),
    .B1(_03093_),
    .X(_01300_));
 sky130_fd_sc_hd__buf_1 _33039_ (.A(_03059_),
    .X(_03094_));
 sky130_fd_sc_hd__and2_4 _33040_ (.A(_02759_),
    .B(_03045_),
    .X(_03095_));
 sky130_fd_sc_hd__a21o_4 _33041_ (.A1(\cpuregs[7][28] ),
    .A2(_03094_),
    .B1(_03095_),
    .X(_01301_));
 sky130_fd_sc_hd__a41oi_4 _33042_ (.A1(_02966_),
    .A2(_02967_),
    .A3(_02968_),
    .A4(_02969_),
    .B1(_03091_),
    .Y(_03096_));
 sky130_fd_sc_hd__a21o_4 _33043_ (.A1(\cpuregs[7][29] ),
    .A2(_03094_),
    .B1(_03096_),
    .X(_01302_));
 sky130_fd_sc_hd__a41oi_4 _33044_ (.A1(_02971_),
    .A2(_02972_),
    .A3(_02973_),
    .A4(_02974_),
    .B1(_03091_),
    .Y(_03097_));
 sky130_fd_sc_hd__a21o_4 _33045_ (.A1(\cpuregs[7][30] ),
    .A2(_03094_),
    .B1(_03097_),
    .X(_01304_));
 sky130_fd_sc_hd__a41oi_4 _33046_ (.A1(_02976_),
    .A2(_02977_),
    .A3(_02978_),
    .A4(_02979_),
    .B1(_03047_),
    .Y(_03098_));
 sky130_fd_sc_hd__a21o_4 _33047_ (.A1(\cpuregs[7][31] ),
    .A2(_03094_),
    .B1(_03098_),
    .X(_01305_));
 sky130_fd_sc_hd__and4_4 _33048_ (.A(_02241_),
    .B(_01766_),
    .C(_02242_),
    .D(_03043_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_1 _33049_ (.A(_03099_),
    .X(_03100_));
 sky130_vsdinv _33050_ (.A(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__buf_1 _33051_ (.A(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_1 _33052_ (.A(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__nor2_4 _33053_ (.A(_02249_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__a21o_4 _33054_ (.A1(\cpuregs[6][0] ),
    .A2(_03103_),
    .B1(_03104_),
    .X(_01249_));
 sky130_fd_sc_hd__buf_1 _33055_ (.A(_03100_),
    .X(_03105_));
 sky130_fd_sc_hd__buf_1 _33056_ (.A(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_1 _33057_ (.A(_03100_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_1 _33058_ (.A(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__nand2_4 _33059_ (.A(_02989_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__o21ai_4 _33060_ (.A1(_19362_),
    .A2(_03106_),
    .B1(_03109_),
    .Y(_01260_));
 sky130_fd_sc_hd__a41o_4 _33061_ (.A1(_02459_),
    .A2(_02597_),
    .A3(_02461_),
    .A4(_02463_),
    .B1(_03103_),
    .X(_03110_));
 sky130_fd_sc_hd__o21ai_4 _33062_ (.A1(_19458_),
    .A2(_03106_),
    .B1(_03110_),
    .Y(_01271_));
 sky130_fd_sc_hd__a41o_4 _33063_ (.A1(_02599_),
    .A2(_02262_),
    .A3(_02264_),
    .A4(_02266_),
    .B1(_03103_),
    .X(_03111_));
 sky130_fd_sc_hd__o21ai_4 _33064_ (.A1(_19535_),
    .A2(_03106_),
    .B1(_03111_),
    .Y(_01274_));
 sky130_fd_sc_hd__buf_1 _33065_ (.A(_23486_),
    .X(_03112_));
 sky130_fd_sc_hd__buf_1 _33066_ (.A(_03102_),
    .X(_03113_));
 sky130_fd_sc_hd__a41o_4 _33067_ (.A1(_02601_),
    .A2(_03112_),
    .A3(_02602_),
    .A4(_02603_),
    .B1(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__o21ai_4 _33068_ (.A1(_19617_),
    .A2(_03106_),
    .B1(_03114_),
    .Y(_01275_));
 sky130_fd_sc_hd__buf_1 _33069_ (.A(_03100_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_1 _33070_ (.A(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_1 _33071_ (.A(_23493_),
    .X(_03117_));
 sky130_fd_sc_hd__a41o_4 _33072_ (.A1(_02608_),
    .A2(_03117_),
    .A3(_02609_),
    .A4(_02610_),
    .B1(_03113_),
    .X(_03118_));
 sky130_fd_sc_hd__o21ai_4 _33073_ (.A1(_19679_),
    .A2(_03116_),
    .B1(_03118_),
    .Y(_01276_));
 sky130_fd_sc_hd__buf_1 _33074_ (.A(_23503_),
    .X(_03119_));
 sky130_fd_sc_hd__a41o_4 _33075_ (.A1(_02612_),
    .A2(_03119_),
    .A3(_02613_),
    .A4(_02614_),
    .B1(_03113_),
    .X(_03120_));
 sky130_fd_sc_hd__o21ai_4 _33076_ (.A1(_19729_),
    .A2(_03116_),
    .B1(_03120_),
    .Y(_01277_));
 sky130_fd_sc_hd__buf_1 _33077_ (.A(_23509_),
    .X(_03121_));
 sky130_fd_sc_hd__a41o_4 _33078_ (.A1(_02616_),
    .A2(_03121_),
    .A3(_02617_),
    .A4(_02618_),
    .B1(_03113_),
    .X(_03122_));
 sky130_fd_sc_hd__o21ai_4 _33079_ (.A1(_19778_),
    .A2(_03116_),
    .B1(_03122_),
    .Y(_01278_));
 sky130_fd_sc_hd__buf_1 _33080_ (.A(_23518_),
    .X(_03123_));
 sky130_fd_sc_hd__buf_1 _33081_ (.A(_03102_),
    .X(_03124_));
 sky130_fd_sc_hd__a41o_4 _33082_ (.A1(_02620_),
    .A2(_03123_),
    .A3(_02621_),
    .A4(_02622_),
    .B1(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__o21ai_4 _33083_ (.A1(_19840_),
    .A2(_03116_),
    .B1(_03125_),
    .Y(_01279_));
 sky130_fd_sc_hd__buf_1 _33084_ (.A(_03115_),
    .X(_03126_));
 sky130_fd_sc_hd__buf_1 _33085_ (.A(_23525_),
    .X(_03127_));
 sky130_fd_sc_hd__a41o_4 _33086_ (.A1(_02626_),
    .A2(_03127_),
    .A3(_02627_),
    .A4(_02628_),
    .B1(_03124_),
    .X(_03128_));
 sky130_fd_sc_hd__o21ai_4 _33087_ (.A1(_19900_),
    .A2(_03126_),
    .B1(_03128_),
    .Y(_01280_));
 sky130_fd_sc_hd__buf_1 _33088_ (.A(_23535_),
    .X(_03129_));
 sky130_fd_sc_hd__a41o_4 _33089_ (.A1(_02630_),
    .A2(_03129_),
    .A3(_02631_),
    .A4(_02632_),
    .B1(_03124_),
    .X(_03130_));
 sky130_fd_sc_hd__o21ai_4 _33090_ (.A1(_19941_),
    .A2(_03126_),
    .B1(_03130_),
    .Y(_01250_));
 sky130_fd_sc_hd__buf_1 _33091_ (.A(_23541_),
    .X(_03131_));
 sky130_fd_sc_hd__a41o_4 _33092_ (.A1(_02634_),
    .A2(_03131_),
    .A3(_02635_),
    .A4(_02636_),
    .B1(_03124_),
    .X(_03132_));
 sky130_fd_sc_hd__o21ai_4 _33093_ (.A1(_20019_),
    .A2(_03126_),
    .B1(_03132_),
    .Y(_01251_));
 sky130_fd_sc_hd__buf_1 _33094_ (.A(_23549_),
    .X(_03133_));
 sky130_fd_sc_hd__buf_1 _33095_ (.A(_03101_),
    .X(_03134_));
 sky130_fd_sc_hd__a41o_4 _33096_ (.A1(_02638_),
    .A2(_03133_),
    .A3(_02639_),
    .A4(_02640_),
    .B1(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__o21ai_4 _33097_ (.A1(_20094_),
    .A2(_03126_),
    .B1(_03135_),
    .Y(_01252_));
 sky130_fd_sc_hd__buf_1 _33098_ (.A(_03115_),
    .X(_03136_));
 sky130_fd_sc_hd__buf_1 _33099_ (.A(_23556_),
    .X(_03137_));
 sky130_fd_sc_hd__a41o_4 _33100_ (.A1(_02644_),
    .A2(_03137_),
    .A3(_02645_),
    .A4(_02646_),
    .B1(_03134_),
    .X(_03138_));
 sky130_fd_sc_hd__o21ai_4 _33101_ (.A1(_20145_),
    .A2(_03136_),
    .B1(_03138_),
    .Y(_01253_));
 sky130_fd_sc_hd__buf_1 _33102_ (.A(_23566_),
    .X(_03139_));
 sky130_fd_sc_hd__a41o_4 _33103_ (.A1(_02648_),
    .A2(_03139_),
    .A3(_02649_),
    .A4(_02650_),
    .B1(_03134_),
    .X(_03140_));
 sky130_fd_sc_hd__o21ai_4 _33104_ (.A1(_20211_),
    .A2(_03136_),
    .B1(_03140_),
    .Y(_01254_));
 sky130_fd_sc_hd__buf_1 _33105_ (.A(_23572_),
    .X(_03141_));
 sky130_fd_sc_hd__a41o_4 _33106_ (.A1(_02652_),
    .A2(_03141_),
    .A3(_02653_),
    .A4(_02654_),
    .B1(_03134_),
    .X(_03142_));
 sky130_fd_sc_hd__o21ai_4 _33107_ (.A1(_20258_),
    .A2(_03136_),
    .B1(_03142_),
    .Y(_01255_));
 sky130_fd_sc_hd__buf_1 _33108_ (.A(_23581_),
    .X(_03143_));
 sky130_fd_sc_hd__buf_1 _33109_ (.A(_03101_),
    .X(_03144_));
 sky130_fd_sc_hd__a41o_4 _33110_ (.A1(_02656_),
    .A2(_03143_),
    .A3(_02657_),
    .A4(_02658_),
    .B1(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__o21ai_4 _33111_ (.A1(_20308_),
    .A2(_03136_),
    .B1(_03145_),
    .Y(_01256_));
 sky130_fd_sc_hd__buf_1 _33112_ (.A(_03115_),
    .X(_03146_));
 sky130_fd_sc_hd__buf_1 _33113_ (.A(_23589_),
    .X(_03147_));
 sky130_fd_sc_hd__a41o_4 _33114_ (.A1(_02662_),
    .A2(_03147_),
    .A3(_02663_),
    .A4(_02664_),
    .B1(_03144_),
    .X(_03148_));
 sky130_fd_sc_hd__o21ai_4 _33115_ (.A1(_20358_),
    .A2(_03146_),
    .B1(_03148_),
    .Y(_01257_));
 sky130_fd_sc_hd__buf_1 _33116_ (.A(_03107_),
    .X(_03149_));
 sky130_fd_sc_hd__nand2_4 _33117_ (.A(_03017_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__o21ai_4 _33118_ (.A1(_20413_),
    .A2(_03146_),
    .B1(_03150_),
    .Y(_01258_));
 sky130_fd_sc_hd__buf_1 _33119_ (.A(_23604_),
    .X(_03151_));
 sky130_fd_sc_hd__a41o_4 _33120_ (.A1(_02668_),
    .A2(_03151_),
    .A3(_02669_),
    .A4(_02670_),
    .B1(_03144_),
    .X(_03152_));
 sky130_fd_sc_hd__o21ai_4 _33121_ (.A1(_20463_),
    .A2(_03146_),
    .B1(_03152_),
    .Y(_01259_));
 sky130_fd_sc_hd__buf_1 _33122_ (.A(_23612_),
    .X(_03153_));
 sky130_fd_sc_hd__a41o_4 _33123_ (.A1(_02672_),
    .A2(_03153_),
    .A3(_02673_),
    .A4(_02674_),
    .B1(_03144_),
    .X(_03154_));
 sky130_fd_sc_hd__o21ai_4 _33124_ (.A1(_20507_),
    .A2(_03146_),
    .B1(_03154_),
    .Y(_01261_));
 sky130_fd_sc_hd__buf_1 _33125_ (.A(_03107_),
    .X(_03155_));
 sky130_fd_sc_hd__buf_1 _33126_ (.A(_23619_),
    .X(_03156_));
 sky130_fd_sc_hd__buf_1 _33127_ (.A(_03101_),
    .X(_03157_));
 sky130_fd_sc_hd__a41o_4 _33128_ (.A1(_02677_),
    .A2(_03156_),
    .A3(_02678_),
    .A4(_02679_),
    .B1(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__o21ai_4 _33129_ (.A1(_20558_),
    .A2(_03155_),
    .B1(_03158_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_4 _33130_ (.A(_03024_),
    .B(_03149_),
    .Y(_03159_));
 sky130_fd_sc_hd__o21ai_4 _33131_ (.A1(_20584_),
    .A2(_03155_),
    .B1(_03159_),
    .Y(_01263_));
 sky130_fd_sc_hd__buf_1 _33132_ (.A(_23632_),
    .X(_03160_));
 sky130_fd_sc_hd__a41o_4 _33133_ (.A1(_02683_),
    .A2(_03160_),
    .A3(_02684_),
    .A4(_02685_),
    .B1(_03157_),
    .X(_03161_));
 sky130_fd_sc_hd__o21ai_4 _33134_ (.A1(_20641_),
    .A2(_03155_),
    .B1(_03161_),
    .Y(_01264_));
 sky130_fd_sc_hd__buf_1 _33135_ (.A(_23640_),
    .X(_03162_));
 sky130_fd_sc_hd__a41o_4 _33136_ (.A1(_02687_),
    .A2(_03162_),
    .A3(_02688_),
    .A4(_02689_),
    .B1(_03157_),
    .X(_03163_));
 sky130_fd_sc_hd__o21ai_4 _33137_ (.A1(_20687_),
    .A2(_03155_),
    .B1(_03163_),
    .Y(_01265_));
 sky130_fd_sc_hd__buf_1 _33138_ (.A(_03107_),
    .X(_03164_));
 sky130_fd_sc_hd__buf_1 _33139_ (.A(_23647_),
    .X(_03165_));
 sky130_fd_sc_hd__a41o_4 _33140_ (.A1(_02692_),
    .A2(_03165_),
    .A3(_02693_),
    .A4(_02694_),
    .B1(_03157_),
    .X(_03166_));
 sky130_fd_sc_hd__o21ai_4 _33141_ (.A1(_20734_),
    .A2(_03164_),
    .B1(_03166_),
    .Y(_01266_));
 sky130_fd_sc_hd__buf_1 _33142_ (.A(_23655_),
    .X(_03167_));
 sky130_fd_sc_hd__a41o_4 _33143_ (.A1(_02696_),
    .A2(_03167_),
    .A3(_02697_),
    .A4(_02698_),
    .B1(_03102_),
    .X(_03168_));
 sky130_fd_sc_hd__o21ai_4 _33144_ (.A1(_20777_),
    .A2(_03164_),
    .B1(_03168_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_4 _33145_ (.A(_03032_),
    .B(_03149_),
    .Y(_03169_));
 sky130_fd_sc_hd__o21ai_4 _33146_ (.A1(_20809_),
    .A2(_03164_),
    .B1(_03169_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand2_4 _33147_ (.A(_03035_),
    .B(_03149_),
    .Y(_03170_));
 sky130_fd_sc_hd__o21ai_4 _33148_ (.A1(_20866_),
    .A2(_03164_),
    .B1(_03170_),
    .Y(_01269_));
 sky130_fd_sc_hd__nand2_4 _33149_ (.A(_03037_),
    .B(_03105_),
    .Y(_03171_));
 sky130_fd_sc_hd__o21ai_4 _33150_ (.A1(_20915_),
    .A2(_03108_),
    .B1(_03171_),
    .Y(_01270_));
 sky130_fd_sc_hd__nand2_4 _33151_ (.A(_03039_),
    .B(_03105_),
    .Y(_03172_));
 sky130_fd_sc_hd__o21ai_4 _33152_ (.A1(_20955_),
    .A2(_03108_),
    .B1(_03172_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_4 _33153_ (.A(_03041_),
    .B(_03105_),
    .Y(_03173_));
 sky130_fd_sc_hd__o21ai_4 _33154_ (.A1(_20998_),
    .A2(_03108_),
    .B1(_03173_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor4_4 _33155_ (.A(_02705_),
    .B(_01787_),
    .C(_03044_),
    .D(_02818_),
    .Y(_03174_));
 sky130_vsdinv _33156_ (.A(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__buf_1 _33157_ (.A(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__buf_1 _33158_ (.A(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__nor3_4 _33159_ (.A(_03049_),
    .B(_02248_),
    .C(_02393_),
    .Y(_03178_));
 sky130_fd_sc_hd__a21o_4 _33160_ (.A1(\cpuregs[5][0] ),
    .A2(_03177_),
    .B1(_03178_),
    .X(_01217_));
 sky130_fd_sc_hd__and2_4 _33161_ (.A(_03174_),
    .B(_02253_),
    .X(_03179_));
 sky130_fd_sc_hd__a21o_4 _33162_ (.A1(\cpuregs[5][1] ),
    .A2(_03177_),
    .B1(_03179_),
    .X(_01228_));
 sky130_fd_sc_hd__buf_1 _33163_ (.A(_03175_),
    .X(_03180_));
 sky130_fd_sc_hd__buf_1 _33164_ (.A(_03180_),
    .X(_03181_));
 sky130_fd_sc_hd__nor2_4 _33165_ (.A(_03181_),
    .B(_02827_),
    .Y(_03182_));
 sky130_fd_sc_hd__a21o_4 _33166_ (.A1(\cpuregs[5][2] ),
    .A2(_03177_),
    .B1(_03182_),
    .X(_01239_));
 sky130_fd_sc_hd__buf_1 _33167_ (.A(_01828_),
    .X(_03183_));
 sky130_fd_sc_hd__nor2_4 _33168_ (.A(_03181_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__a21o_4 _33169_ (.A1(\cpuregs[5][3] ),
    .A2(_03177_),
    .B1(_03184_),
    .X(_01242_));
 sky130_fd_sc_hd__buf_1 _33170_ (.A(_03176_),
    .X(_03185_));
 sky130_fd_sc_hd__a41oi_4 _33171_ (.A1(_02831_),
    .A2(_02832_),
    .A3(_02833_),
    .A4(_02834_),
    .B1(_03181_),
    .Y(_03186_));
 sky130_fd_sc_hd__a21o_4 _33172_ (.A1(\cpuregs[5][4] ),
    .A2(_03185_),
    .B1(_03186_),
    .X(_01243_));
 sky130_fd_sc_hd__a41oi_4 _33173_ (.A1(_02836_),
    .A2(_02837_),
    .A3(_02838_),
    .A4(_02839_),
    .B1(_03181_),
    .Y(_03187_));
 sky130_fd_sc_hd__a21o_4 _33174_ (.A1(\cpuregs[5][5] ),
    .A2(_03185_),
    .B1(_03187_),
    .X(_01244_));
 sky130_fd_sc_hd__buf_1 _33175_ (.A(_03175_),
    .X(_03188_));
 sky130_fd_sc_hd__buf_1 _33176_ (.A(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__a41oi_4 _33177_ (.A1(_02841_),
    .A2(_02842_),
    .A3(_02843_),
    .A4(_02844_),
    .B1(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__a21o_4 _33178_ (.A1(\cpuregs[5][6] ),
    .A2(_03185_),
    .B1(_03190_),
    .X(_01245_));
 sky130_fd_sc_hd__a41oi_4 _33179_ (.A1(_02848_),
    .A2(_02849_),
    .A3(_02850_),
    .A4(_02851_),
    .B1(_03189_),
    .Y(_03191_));
 sky130_fd_sc_hd__a21o_4 _33180_ (.A1(\cpuregs[5][7] ),
    .A2(_03185_),
    .B1(_03191_),
    .X(_01246_));
 sky130_fd_sc_hd__buf_1 _33181_ (.A(_03176_),
    .X(_03192_));
 sky130_fd_sc_hd__a41oi_4 _33182_ (.A1(_02854_),
    .A2(_02855_),
    .A3(_02856_),
    .A4(_02857_),
    .B1(_03189_),
    .Y(_03193_));
 sky130_fd_sc_hd__a21o_4 _33183_ (.A1(\cpuregs[5][8] ),
    .A2(_03192_),
    .B1(_03193_),
    .X(_01247_));
 sky130_fd_sc_hd__a41oi_4 _33184_ (.A1(_02859_),
    .A2(_02860_),
    .A3(_02861_),
    .A4(_02862_),
    .B1(_03189_),
    .Y(_03194_));
 sky130_fd_sc_hd__a21o_4 _33185_ (.A1(\cpuregs[5][9] ),
    .A2(_03192_),
    .B1(_03194_),
    .X(_01248_));
 sky130_fd_sc_hd__buf_1 _33186_ (.A(_03188_),
    .X(_03195_));
 sky130_fd_sc_hd__a41oi_4 _33187_ (.A1(_02864_),
    .A2(_02865_),
    .A3(_02866_),
    .A4(_02867_),
    .B1(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__a21o_4 _33188_ (.A1(\cpuregs[5][10] ),
    .A2(_03192_),
    .B1(_03196_),
    .X(_01218_));
 sky130_fd_sc_hd__a41oi_4 _33189_ (.A1(_02870_),
    .A2(_02871_),
    .A3(_02872_),
    .A4(_02873_),
    .B1(_03195_),
    .Y(_03197_));
 sky130_fd_sc_hd__a21o_4 _33190_ (.A1(\cpuregs[5][11] ),
    .A2(_03192_),
    .B1(_03197_),
    .X(_01219_));
 sky130_fd_sc_hd__buf_1 _33191_ (.A(_03175_),
    .X(_03198_));
 sky130_fd_sc_hd__buf_1 _33192_ (.A(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__a41oi_4 _33193_ (.A1(_02877_),
    .A2(_02878_),
    .A3(_02879_),
    .A4(_02880_),
    .B1(_03195_),
    .Y(_03200_));
 sky130_fd_sc_hd__a21o_4 _33194_ (.A1(\cpuregs[5][12] ),
    .A2(_03199_),
    .B1(_03200_),
    .X(_01220_));
 sky130_fd_sc_hd__a41oi_4 _33195_ (.A1(_02882_),
    .A2(_02883_),
    .A3(_02884_),
    .A4(_02885_),
    .B1(_03195_),
    .Y(_03201_));
 sky130_fd_sc_hd__a21o_4 _33196_ (.A1(\cpuregs[5][13] ),
    .A2(_03199_),
    .B1(_03201_),
    .X(_01221_));
 sky130_fd_sc_hd__buf_1 _33197_ (.A(_03188_),
    .X(_03202_));
 sky130_fd_sc_hd__a41oi_4 _33198_ (.A1(_02887_),
    .A2(_02888_),
    .A3(_02889_),
    .A4(_02890_),
    .B1(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__a21o_4 _33199_ (.A1(\cpuregs[5][14] ),
    .A2(_03199_),
    .B1(_03203_),
    .X(_01222_));
 sky130_fd_sc_hd__a41oi_4 _33200_ (.A1(_02893_),
    .A2(_02894_),
    .A3(_02895_),
    .A4(_02896_),
    .B1(_03202_),
    .Y(_03204_));
 sky130_fd_sc_hd__a21o_4 _33201_ (.A1(\cpuregs[5][15] ),
    .A2(_03199_),
    .B1(_03204_),
    .X(_01223_));
 sky130_fd_sc_hd__buf_1 _33202_ (.A(_03198_),
    .X(_03205_));
 sky130_fd_sc_hd__a41oi_4 _33203_ (.A1(_02899_),
    .A2(_02900_),
    .A3(_02901_),
    .A4(_02902_),
    .B1(_03202_),
    .Y(_03206_));
 sky130_fd_sc_hd__a21o_4 _33204_ (.A1(\cpuregs[5][16] ),
    .A2(_03205_),
    .B1(_03206_),
    .X(_01224_));
 sky130_fd_sc_hd__a41oi_4 _33205_ (.A1(_02904_),
    .A2(_02905_),
    .A3(_02906_),
    .A4(_02907_),
    .B1(_03202_),
    .Y(_03207_));
 sky130_fd_sc_hd__a21o_4 _33206_ (.A1(\cpuregs[5][17] ),
    .A2(_03205_),
    .B1(_03207_),
    .X(_01225_));
 sky130_fd_sc_hd__buf_1 _33207_ (.A(_03180_),
    .X(_03208_));
 sky130_fd_sc_hd__a41oi_4 _33208_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_02911_),
    .A4(_02912_),
    .B1(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__a21o_4 _33209_ (.A1(\cpuregs[5][18] ),
    .A2(_03205_),
    .B1(_03209_),
    .X(_01226_));
 sky130_fd_sc_hd__a41oi_4 _33210_ (.A1(_02915_),
    .A2(_02916_),
    .A3(_02917_),
    .A4(_02918_),
    .B1(_03208_),
    .Y(_03210_));
 sky130_fd_sc_hd__a21o_4 _33211_ (.A1(\cpuregs[5][19] ),
    .A2(_03205_),
    .B1(_03210_),
    .X(_01227_));
 sky130_fd_sc_hd__buf_1 _33212_ (.A(_03198_),
    .X(_03211_));
 sky130_fd_sc_hd__a41oi_4 _33213_ (.A1(_02921_),
    .A2(_02922_),
    .A3(_02923_),
    .A4(_02924_),
    .B1(_03208_),
    .Y(_03212_));
 sky130_fd_sc_hd__a21o_4 _33214_ (.A1(\cpuregs[5][20] ),
    .A2(_03211_),
    .B1(_03212_),
    .X(_01229_));
 sky130_fd_sc_hd__a41oi_4 _33215_ (.A1(_02926_),
    .A2(_02927_),
    .A3(_02928_),
    .A4(_02929_),
    .B1(_03208_),
    .Y(_03213_));
 sky130_fd_sc_hd__a21o_4 _33216_ (.A1(\cpuregs[5][21] ),
    .A2(_03211_),
    .B1(_03213_),
    .X(_01230_));
 sky130_fd_sc_hd__buf_1 _33217_ (.A(_03180_),
    .X(_03214_));
 sky130_fd_sc_hd__a41oi_4 _33218_ (.A1(_02931_),
    .A2(_02932_),
    .A3(_02933_),
    .A4(_02934_),
    .B1(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__a21o_4 _33219_ (.A1(\cpuregs[5][22] ),
    .A2(_03211_),
    .B1(_03215_),
    .X(_01231_));
 sky130_fd_sc_hd__a41oi_4 _33220_ (.A1(_02937_),
    .A2(_02938_),
    .A3(_02939_),
    .A4(_02940_),
    .B1(_03214_),
    .Y(_03216_));
 sky130_fd_sc_hd__a21o_4 _33221_ (.A1(\cpuregs[5][23] ),
    .A2(_03211_),
    .B1(_03216_),
    .X(_01232_));
 sky130_fd_sc_hd__buf_1 _33222_ (.A(_03198_),
    .X(_03217_));
 sky130_fd_sc_hd__a41oi_4 _33223_ (.A1(_02943_),
    .A2(_02944_),
    .A3(_02945_),
    .A4(_02946_),
    .B1(_03214_),
    .Y(_03218_));
 sky130_fd_sc_hd__a21o_4 _33224_ (.A1(\cpuregs[5][24] ),
    .A2(_03217_),
    .B1(_03218_),
    .X(_01233_));
 sky130_fd_sc_hd__a41oi_4 _33225_ (.A1(_02948_),
    .A2(_02949_),
    .A3(_02950_),
    .A4(_02951_),
    .B1(_03214_),
    .Y(_03219_));
 sky130_fd_sc_hd__a21o_4 _33226_ (.A1(\cpuregs[5][25] ),
    .A2(_03217_),
    .B1(_03219_),
    .X(_01234_));
 sky130_fd_sc_hd__buf_1 _33227_ (.A(_03180_),
    .X(_03220_));
 sky130_fd_sc_hd__a41oi_4 _33228_ (.A1(_02953_),
    .A2(_02954_),
    .A3(_02955_),
    .A4(_02956_),
    .B1(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__a21o_4 _33229_ (.A1(\cpuregs[5][26] ),
    .A2(_03217_),
    .B1(_03221_),
    .X(_01235_));
 sky130_fd_sc_hd__a41oi_4 _33230_ (.A1(_02959_),
    .A2(_02960_),
    .A3(_02961_),
    .A4(_02962_),
    .B1(_03220_),
    .Y(_03222_));
 sky130_fd_sc_hd__a21o_4 _33231_ (.A1(\cpuregs[5][27] ),
    .A2(_03217_),
    .B1(_03222_),
    .X(_01236_));
 sky130_fd_sc_hd__buf_1 _33232_ (.A(_03188_),
    .X(_03223_));
 sky130_fd_sc_hd__and2_4 _33233_ (.A(_02759_),
    .B(_03174_),
    .X(_03224_));
 sky130_fd_sc_hd__a21o_4 _33234_ (.A1(\cpuregs[5][28] ),
    .A2(_03223_),
    .B1(_03224_),
    .X(_01237_));
 sky130_fd_sc_hd__a41oi_4 _33235_ (.A1(_02966_),
    .A2(_02967_),
    .A3(_02968_),
    .A4(_02969_),
    .B1(_03220_),
    .Y(_03225_));
 sky130_fd_sc_hd__a21o_4 _33236_ (.A1(\cpuregs[5][29] ),
    .A2(_03223_),
    .B1(_03225_),
    .X(_01238_));
 sky130_fd_sc_hd__a41oi_4 _33237_ (.A1(_02971_),
    .A2(_02972_),
    .A3(_02973_),
    .A4(_02974_),
    .B1(_03220_),
    .Y(_03226_));
 sky130_fd_sc_hd__a21o_4 _33238_ (.A1(\cpuregs[5][30] ),
    .A2(_03223_),
    .B1(_03226_),
    .X(_01240_));
 sky130_fd_sc_hd__a41oi_4 _33239_ (.A1(_02976_),
    .A2(_02977_),
    .A3(_02978_),
    .A4(_02979_),
    .B1(_03176_),
    .Y(_03227_));
 sky130_fd_sc_hd__a21o_4 _33240_ (.A1(\cpuregs[5][31] ),
    .A2(_03223_),
    .B1(_03227_),
    .X(_01241_));
 sky130_fd_sc_hd__buf_1 _33241_ (.A(\pcpi_mul.rs1[0] ),
    .X(_03228_));
 sky130_vsdinv _33242_ (.A(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__and4_4 _33243_ (.A(_18822_),
    .B(_18814_),
    .C(_18823_),
    .D(_18824_),
    .X(_03230_));
 sky130_fd_sc_hd__nor2_4 _33244_ (.A(_18810_),
    .B(_18813_),
    .Y(_03231_));
 sky130_fd_sc_hd__nor2_4 _33245_ (.A(\pcpi_mul.active[1] ),
    .B(\pcpi_mul.active[0] ),
    .Y(_03232_));
 sky130_fd_sc_hd__and3_4 _33246_ (.A(_03230_),
    .B(_03231_),
    .C(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__buf_1 _33247_ (.A(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__buf_1 _33248_ (.A(_03234_),
    .X(_00669_));
 sky130_fd_sc_hd__buf_1 _33249_ (.A(_03230_),
    .X(_03235_));
 sky130_fd_sc_hd__buf_1 _33250_ (.A(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_1 _33251_ (.A(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__buf_1 _33252_ (.A(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__buf_1 _33253_ (.A(_03231_),
    .X(_03239_));
 sky130_fd_sc_hd__buf_1 _33254_ (.A(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__buf_1 _33255_ (.A(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__buf_1 _33256_ (.A(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__buf_1 _33257_ (.A(_03232_),
    .X(_03243_));
 sky130_fd_sc_hd__buf_1 _33258_ (.A(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__buf_1 _33259_ (.A(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__buf_1 _33260_ (.A(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__nand4_4 _33261_ (.A(_21351_),
    .B(_03238_),
    .C(_03242_),
    .D(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__o21ai_4 _33262_ (.A1(_03229_),
    .A2(_00669_),
    .B1(_03247_),
    .Y(_00671_));
 sky130_fd_sc_hd__buf_1 _33263_ (.A(\pcpi_mul.rs1[1] ),
    .X(_03248_));
 sky130_vsdinv _33264_ (.A(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__buf_1 _33265_ (.A(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__nand4_4 _33266_ (.A(_21380_),
    .B(_03238_),
    .C(_03242_),
    .D(_03246_),
    .Y(_03251_));
 sky130_fd_sc_hd__o21ai_4 _33267_ (.A1(_03250_),
    .A2(_00669_),
    .B1(_03251_),
    .Y(_00682_));
 sky130_fd_sc_hd__buf_1 _33268_ (.A(\pcpi_mul.rs1[2] ),
    .X(_03252_));
 sky130_fd_sc_hd__buf_1 _33269_ (.A(_03252_),
    .X(_03253_));
 sky130_vsdinv _33270_ (.A(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand4_4 _33271_ (.A(_21397_),
    .B(_03238_),
    .C(_03242_),
    .D(_03246_),
    .Y(_03255_));
 sky130_fd_sc_hd__o21ai_4 _33272_ (.A1(_03254_),
    .A2(_00669_),
    .B1(_03255_),
    .Y(_00693_));
 sky130_fd_sc_hd__buf_1 _33273_ (.A(\pcpi_mul.rs1[3] ),
    .X(_03256_));
 sky130_vsdinv _33274_ (.A(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__buf_1 _33275_ (.A(_03233_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_1 _33276_ (.A(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__nand4_4 _33277_ (.A(_21421_),
    .B(_03238_),
    .C(_03242_),
    .D(_03246_),
    .Y(_03260_));
 sky130_fd_sc_hd__o21ai_4 _33278_ (.A1(_03257_),
    .A2(_03259_),
    .B1(_03260_),
    .Y(_00697_));
 sky130_fd_sc_hd__buf_1 _33279_ (.A(\pcpi_mul.rs1[4] ),
    .X(_03261_));
 sky130_vsdinv _33280_ (.A(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__buf_1 _33281_ (.A(_03237_),
    .X(_03263_));
 sky130_fd_sc_hd__buf_1 _33282_ (.A(_03241_),
    .X(_03264_));
 sky130_fd_sc_hd__buf_1 _33283_ (.A(_03245_),
    .X(_03265_));
 sky130_fd_sc_hd__nand4_4 _33284_ (.A(_21434_),
    .B(_03263_),
    .C(_03264_),
    .D(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__o21ai_4 _33285_ (.A1(_03262_),
    .A2(_03259_),
    .B1(_03266_),
    .Y(_00698_));
 sky130_fd_sc_hd__buf_1 _33286_ (.A(\pcpi_mul.rs1[5] ),
    .X(_03267_));
 sky130_fd_sc_hd__buf_1 _33287_ (.A(_03267_),
    .X(_03268_));
 sky130_vsdinv _33288_ (.A(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand4_4 _33289_ (.A(_21462_),
    .B(_03263_),
    .C(_03264_),
    .D(_03265_),
    .Y(_03270_));
 sky130_fd_sc_hd__o21ai_4 _33290_ (.A1(_03269_),
    .A2(_03259_),
    .B1(_03270_),
    .Y(_00699_));
 sky130_fd_sc_hd__buf_1 _33291_ (.A(\pcpi_mul.rs1[6] ),
    .X(_03271_));
 sky130_vsdinv _33292_ (.A(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__nand4_4 _33293_ (.A(_21479_),
    .B(_03263_),
    .C(_03264_),
    .D(_03265_),
    .Y(_03273_));
 sky130_fd_sc_hd__o21ai_4 _33294_ (.A1(_03272_),
    .A2(_03259_),
    .B1(_03273_),
    .Y(_00700_));
 sky130_fd_sc_hd__buf_1 _33295_ (.A(\pcpi_mul.rs1[7] ),
    .X(_03274_));
 sky130_fd_sc_hd__buf_1 _33296_ (.A(_03274_),
    .X(_03275_));
 sky130_vsdinv _33297_ (.A(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__buf_1 _33298_ (.A(_03258_),
    .X(_03277_));
 sky130_fd_sc_hd__nand4_4 _33299_ (.A(_21493_),
    .B(_03263_),
    .C(_03264_),
    .D(_03265_),
    .Y(_03278_));
 sky130_fd_sc_hd__o21ai_4 _33300_ (.A1(_03276_),
    .A2(_03277_),
    .B1(_03278_),
    .Y(_00701_));
 sky130_fd_sc_hd__buf_1 _33301_ (.A(\pcpi_mul.rs1[8] ),
    .X(_03279_));
 sky130_fd_sc_hd__buf_1 _33302_ (.A(_03279_),
    .X(_03280_));
 sky130_vsdinv _33303_ (.A(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__buf_1 _33304_ (.A(_03236_),
    .X(_03282_));
 sky130_fd_sc_hd__buf_1 _33305_ (.A(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__buf_1 _33306_ (.A(_03240_),
    .X(_03284_));
 sky130_fd_sc_hd__buf_1 _33307_ (.A(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__buf_1 _33308_ (.A(_03244_),
    .X(_03286_));
 sky130_fd_sc_hd__buf_1 _33309_ (.A(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__nand4_4 _33310_ (.A(_21507_),
    .B(_03283_),
    .C(_03285_),
    .D(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__o21ai_4 _33311_ (.A1(_03281_),
    .A2(_03277_),
    .B1(_03288_),
    .Y(_00702_));
 sky130_fd_sc_hd__buf_1 _33312_ (.A(\pcpi_mul.rs1[9] ),
    .X(_03289_));
 sky130_fd_sc_hd__buf_1 _33313_ (.A(_03289_),
    .X(_03290_));
 sky130_vsdinv _33314_ (.A(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__nand4_4 _33315_ (.A(_21530_),
    .B(_03283_),
    .C(_03285_),
    .D(_03287_),
    .Y(_03292_));
 sky130_fd_sc_hd__o21ai_4 _33316_ (.A1(_03291_),
    .A2(_03277_),
    .B1(_03292_),
    .Y(_00703_));
 sky130_fd_sc_hd__buf_1 _33317_ (.A(\pcpi_mul.rs1[10] ),
    .X(_03293_));
 sky130_fd_sc_hd__buf_1 _33318_ (.A(_03293_),
    .X(_03294_));
 sky130_vsdinv _33319_ (.A(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand4_4 _33320_ (.A(_01611_),
    .B(_03283_),
    .C(_03285_),
    .D(_03287_),
    .Y(_03296_));
 sky130_fd_sc_hd__o21ai_4 _33321_ (.A1(_03295_),
    .A2(_03277_),
    .B1(_03296_),
    .Y(_00672_));
 sky130_fd_sc_hd__buf_1 _33322_ (.A(\pcpi_mul.rs1[11] ),
    .X(_03297_));
 sky130_fd_sc_hd__buf_1 _33323_ (.A(_03297_),
    .X(_03298_));
 sky130_vsdinv _33324_ (.A(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__buf_1 _33325_ (.A(_03258_),
    .X(_03300_));
 sky130_fd_sc_hd__nand4_4 _33326_ (.A(_21565_),
    .B(_03283_),
    .C(_03285_),
    .D(_03287_),
    .Y(_03301_));
 sky130_fd_sc_hd__o21ai_4 _33327_ (.A1(_03299_),
    .A2(_03300_),
    .B1(_03301_),
    .Y(_00673_));
 sky130_fd_sc_hd__buf_1 _33328_ (.A(\pcpi_mul.rs1[12] ),
    .X(_03302_));
 sky130_fd_sc_hd__buf_1 _33329_ (.A(_03302_),
    .X(_03303_));
 sky130_vsdinv _33330_ (.A(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__buf_1 _33331_ (.A(_03282_),
    .X(_03305_));
 sky130_fd_sc_hd__buf_1 _33332_ (.A(_03284_),
    .X(_03306_));
 sky130_fd_sc_hd__buf_1 _33333_ (.A(_03286_),
    .X(_03307_));
 sky130_fd_sc_hd__nand4_4 _33334_ (.A(_21590_),
    .B(_03305_),
    .C(_03306_),
    .D(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__o21ai_4 _33335_ (.A1(_03304_),
    .A2(_03300_),
    .B1(_03308_),
    .Y(_00674_));
 sky130_fd_sc_hd__buf_1 _33336_ (.A(\pcpi_mul.rs1[13] ),
    .X(_03309_));
 sky130_fd_sc_hd__buf_1 _33337_ (.A(_03309_),
    .X(_03310_));
 sky130_vsdinv _33338_ (.A(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand4_4 _33339_ (.A(_21605_),
    .B(_03305_),
    .C(_03306_),
    .D(_03307_),
    .Y(_03312_));
 sky130_fd_sc_hd__o21ai_4 _33340_ (.A1(_03311_),
    .A2(_03300_),
    .B1(_03312_),
    .Y(_00675_));
 sky130_fd_sc_hd__buf_1 _33341_ (.A(\pcpi_mul.rs1[14] ),
    .X(_03313_));
 sky130_fd_sc_hd__buf_1 _33342_ (.A(_03313_),
    .X(_03314_));
 sky130_vsdinv _33343_ (.A(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand4_4 _33344_ (.A(_01630_),
    .B(_03305_),
    .C(_03306_),
    .D(_03307_),
    .Y(_03316_));
 sky130_fd_sc_hd__o21ai_4 _33345_ (.A1(_03315_),
    .A2(_03300_),
    .B1(_03316_),
    .Y(_00676_));
 sky130_fd_sc_hd__buf_1 _33346_ (.A(\pcpi_mul.rs1[15] ),
    .X(_03317_));
 sky130_fd_sc_hd__buf_1 _33347_ (.A(_03317_),
    .X(_03318_));
 sky130_vsdinv _33348_ (.A(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__buf_1 _33349_ (.A(_03234_),
    .X(_03320_));
 sky130_fd_sc_hd__buf_1 _33350_ (.A(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__nand4_4 _33351_ (.A(_01636_),
    .B(_03305_),
    .C(_03306_),
    .D(_03307_),
    .Y(_03322_));
 sky130_fd_sc_hd__o21ai_4 _33352_ (.A1(_03319_),
    .A2(_03321_),
    .B1(_03322_),
    .Y(_00677_));
 sky130_fd_sc_hd__buf_1 _33353_ (.A(\pcpi_mul.rs1[16] ),
    .X(_03323_));
 sky130_fd_sc_hd__buf_1 _33354_ (.A(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__buf_1 _33355_ (.A(_03324_),
    .X(_03325_));
 sky130_vsdinv _33356_ (.A(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__buf_1 _33357_ (.A(_03282_),
    .X(_03327_));
 sky130_fd_sc_hd__buf_1 _33358_ (.A(_03284_),
    .X(_03328_));
 sky130_fd_sc_hd__buf_1 _33359_ (.A(_03286_),
    .X(_03329_));
 sky130_fd_sc_hd__nand4_4 _33360_ (.A(_21678_),
    .B(_03327_),
    .C(_03328_),
    .D(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__o21ai_4 _33361_ (.A1(_03326_),
    .A2(_03321_),
    .B1(_03330_),
    .Y(_00678_));
 sky130_fd_sc_hd__buf_1 _33362_ (.A(\pcpi_mul.rs1[17] ),
    .X(_03331_));
 sky130_fd_sc_hd__buf_1 _33363_ (.A(_03331_),
    .X(_03332_));
 sky130_vsdinv _33364_ (.A(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__nand4_4 _33365_ (.A(_18715_),
    .B(_03327_),
    .C(_03328_),
    .D(_03329_),
    .Y(_03334_));
 sky130_fd_sc_hd__o21ai_4 _33366_ (.A1(_03333_),
    .A2(_03321_),
    .B1(_03334_),
    .Y(_00679_));
 sky130_fd_sc_hd__buf_1 _33367_ (.A(\pcpi_mul.rs1[18] ),
    .X(_03335_));
 sky130_fd_sc_hd__buf_1 _33368_ (.A(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__buf_1 _33369_ (.A(_03336_),
    .X(_03337_));
 sky130_vsdinv _33370_ (.A(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand4_4 _33371_ (.A(_18705_),
    .B(_03327_),
    .C(_03328_),
    .D(_03329_),
    .Y(_03339_));
 sky130_fd_sc_hd__o21ai_4 _33372_ (.A1(_03338_),
    .A2(_03321_),
    .B1(_03339_),
    .Y(_00680_));
 sky130_fd_sc_hd__buf_1 _33373_ (.A(\pcpi_mul.rs1[19] ),
    .X(_03340_));
 sky130_fd_sc_hd__buf_1 _33374_ (.A(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__buf_1 _33375_ (.A(_03341_),
    .X(_03342_));
 sky130_vsdinv _33376_ (.A(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__buf_1 _33377_ (.A(_03320_),
    .X(_03344_));
 sky130_fd_sc_hd__nand4_4 _33378_ (.A(_18694_),
    .B(_03327_),
    .C(_03328_),
    .D(_03329_),
    .Y(_03345_));
 sky130_fd_sc_hd__o21ai_4 _33379_ (.A1(_03343_),
    .A2(_03344_),
    .B1(_03345_),
    .Y(_00681_));
 sky130_fd_sc_hd__buf_1 _33380_ (.A(\pcpi_mul.rs1[20] ),
    .X(_03346_));
 sky130_vsdinv _33381_ (.A(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__buf_1 _33382_ (.A(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__buf_1 _33383_ (.A(_03282_),
    .X(_03349_));
 sky130_fd_sc_hd__buf_1 _33384_ (.A(_03284_),
    .X(_03350_));
 sky130_fd_sc_hd__buf_1 _33385_ (.A(_03286_),
    .X(_03351_));
 sky130_fd_sc_hd__nand4_4 _33386_ (.A(_21721_),
    .B(_03349_),
    .C(_03350_),
    .D(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__o21ai_4 _33387_ (.A1(_03348_),
    .A2(_03344_),
    .B1(_03352_),
    .Y(_00683_));
 sky130_fd_sc_hd__buf_1 _33388_ (.A(\pcpi_mul.rs1[21] ),
    .X(_03353_));
 sky130_vsdinv _33389_ (.A(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__buf_1 _33390_ (.A(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__nand4_4 _33391_ (.A(_21739_),
    .B(_03349_),
    .C(_03350_),
    .D(_03351_),
    .Y(_03356_));
 sky130_fd_sc_hd__o21ai_4 _33392_ (.A1(_03355_),
    .A2(_03344_),
    .B1(_03356_),
    .Y(_00684_));
 sky130_fd_sc_hd__buf_1 _33393_ (.A(\pcpi_mul.rs1[22] ),
    .X(_03357_));
 sky130_fd_sc_hd__buf_1 _33394_ (.A(_03357_),
    .X(_03358_));
 sky130_vsdinv _33395_ (.A(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand4_4 _33396_ (.A(_18676_),
    .B(_03349_),
    .C(_03350_),
    .D(_03351_),
    .Y(_03360_));
 sky130_fd_sc_hd__o21ai_4 _33397_ (.A1(_03359_),
    .A2(_03344_),
    .B1(_03360_),
    .Y(_00685_));
 sky130_fd_sc_hd__buf_1 _33398_ (.A(\pcpi_mul.rs1[23] ),
    .X(_03361_));
 sky130_vsdinv _33399_ (.A(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__buf_1 _33400_ (.A(_03320_),
    .X(_03363_));
 sky130_fd_sc_hd__nand4_4 _33401_ (.A(_01671_),
    .B(_03349_),
    .C(_03350_),
    .D(_03351_),
    .Y(_03364_));
 sky130_fd_sc_hd__o21ai_4 _33402_ (.A1(_03362_),
    .A2(_03363_),
    .B1(_03364_),
    .Y(_00686_));
 sky130_fd_sc_hd__buf_1 _33403_ (.A(\pcpi_mul.rs1[24] ),
    .X(_03365_));
 sky130_vsdinv _33404_ (.A(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__buf_1 _33405_ (.A(_03235_),
    .X(_03367_));
 sky130_fd_sc_hd__buf_1 _33406_ (.A(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__buf_1 _33407_ (.A(_03239_),
    .X(_03369_));
 sky130_fd_sc_hd__buf_1 _33408_ (.A(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__buf_1 _33409_ (.A(_03243_),
    .X(_03371_));
 sky130_fd_sc_hd__buf_1 _33410_ (.A(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__nand4_4 _33411_ (.A(_18732_),
    .B(_03368_),
    .C(_03370_),
    .D(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__o21ai_4 _33412_ (.A1(_03366_),
    .A2(_03363_),
    .B1(_03373_),
    .Y(_00687_));
 sky130_fd_sc_hd__buf_1 _33413_ (.A(\pcpi_mul.rs1[25] ),
    .X(_03374_));
 sky130_fd_sc_hd__buf_1 _33414_ (.A(_03374_),
    .X(_03375_));
 sky130_vsdinv _33415_ (.A(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__buf_1 _33416_ (.A(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__nand4_4 _33417_ (.A(_18766_),
    .B(_03368_),
    .C(_03370_),
    .D(_03372_),
    .Y(_03378_));
 sky130_fd_sc_hd__o21ai_4 _33418_ (.A1(_03377_),
    .A2(_03363_),
    .B1(_03378_),
    .Y(_00688_));
 sky130_fd_sc_hd__buf_1 _33419_ (.A(\pcpi_mul.rs1[26] ),
    .X(_03379_));
 sky130_vsdinv _33420_ (.A(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand4_4 _33421_ (.A(_18721_),
    .B(_03368_),
    .C(_03370_),
    .D(_03372_),
    .Y(_03381_));
 sky130_fd_sc_hd__o21ai_4 _33422_ (.A1(_03380_),
    .A2(_03363_),
    .B1(_03381_),
    .Y(_00689_));
 sky130_fd_sc_hd__buf_1 _33423_ (.A(\pcpi_mul.rs1[27] ),
    .X(_03382_));
 sky130_fd_sc_hd__buf_1 _33424_ (.A(_03382_),
    .X(_03383_));
 sky130_vsdinv _33425_ (.A(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__buf_1 _33426_ (.A(_03320_),
    .X(_03385_));
 sky130_fd_sc_hd__nand4_4 _33427_ (.A(_01689_),
    .B(_03368_),
    .C(_03370_),
    .D(_03372_),
    .Y(_03386_));
 sky130_fd_sc_hd__o21ai_4 _33428_ (.A1(_03384_),
    .A2(_03385_),
    .B1(_03386_),
    .Y(_00690_));
 sky130_fd_sc_hd__buf_1 _33429_ (.A(\pcpi_mul.rs1[28] ),
    .X(_03387_));
 sky130_vsdinv _33430_ (.A(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__buf_1 _33431_ (.A(_03367_),
    .X(_03389_));
 sky130_fd_sc_hd__buf_1 _33432_ (.A(_03369_),
    .X(_03390_));
 sky130_fd_sc_hd__buf_1 _33433_ (.A(_03371_),
    .X(_03391_));
 sky130_fd_sc_hd__nand4_4 _33434_ (.A(_01694_),
    .B(_03389_),
    .C(_03390_),
    .D(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__o21ai_4 _33435_ (.A1(_03388_),
    .A2(_03385_),
    .B1(_03392_),
    .Y(_00691_));
 sky130_fd_sc_hd__buf_1 _33436_ (.A(\pcpi_mul.rs1[29] ),
    .X(_03393_));
 sky130_vsdinv _33437_ (.A(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand4_4 _33438_ (.A(_21879_),
    .B(_03389_),
    .C(_03390_),
    .D(_03391_),
    .Y(_03395_));
 sky130_fd_sc_hd__o21ai_4 _33439_ (.A1(_03394_),
    .A2(_03385_),
    .B1(_03395_),
    .Y(_00692_));
 sky130_fd_sc_hd__buf_1 _33440_ (.A(\pcpi_mul.rs1[30] ),
    .X(_03396_));
 sky130_fd_sc_hd__buf_1 _33441_ (.A(_03396_),
    .X(_03397_));
 sky130_vsdinv _33442_ (.A(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand4_4 _33443_ (.A(_21871_),
    .B(_03389_),
    .C(_03390_),
    .D(_03391_),
    .Y(_03399_));
 sky130_fd_sc_hd__o21ai_4 _33444_ (.A1(_03398_),
    .A2(_03385_),
    .B1(_03399_),
    .Y(_00694_));
 sky130_vsdinv _33445_ (.A(\pcpi_mul.rs1[31] ),
    .Y(_03400_));
 sky130_fd_sc_hd__buf_1 _33446_ (.A(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__buf_1 _33447_ (.A(_03234_),
    .X(_03402_));
 sky130_fd_sc_hd__and4_4 _33448_ (.A(_03235_),
    .B(_21905_),
    .C(_03239_),
    .D(_03243_),
    .X(_03403_));
 sky130_vsdinv _33449_ (.A(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__o21ai_4 _33450_ (.A1(_03401_),
    .A2(_03402_),
    .B1(_03404_),
    .Y(_00695_));
 sky130_fd_sc_hd__buf_1 _33451_ (.A(\pcpi_mul.rs1[32] ),
    .X(_03405_));
 sky130_fd_sc_hd__buf_8 _33452_ (.A(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__buf_8 _33453_ (.A(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__buf_1 _33454_ (.A(_03407_),
    .X(_03408_));
 sky130_fd_sc_hd__buf_1 _33455_ (.A(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__buf_1 _33456_ (.A(_03409_),
    .X(_03410_));
 sky130_vsdinv _33457_ (.A(_03233_),
    .Y(_03411_));
 sky130_fd_sc_hd__buf_1 _33458_ (.A(_03411_),
    .X(_03412_));
 sky130_vsdinv _33459_ (.A(_18826_),
    .Y(_03413_));
 sky130_fd_sc_hd__nor3_4 _33460_ (.A(pcpi_insn[13]),
    .B(_24155_),
    .C(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__o21ai_4 _33461_ (.A1(pcpi_insn[13]),
    .A2(pcpi_insn[12]),
    .B1(_18826_),
    .Y(_03415_));
 sky130_fd_sc_hd__nor2_4 _33462_ (.A(_03415_),
    .B(_03404_),
    .Y(_03416_));
 sky130_fd_sc_hd__o21a_4 _33463_ (.A1(_24155_),
    .A2(_03414_),
    .B1(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__a21o_4 _33464_ (.A1(_03410_),
    .A2(_03412_),
    .B1(_03417_),
    .X(_00696_));
 sky130_fd_sc_hd__buf_1 _33465_ (.A(_03412_),
    .X(_03418_));
 sky130_fd_sc_hd__buf_1 _33466_ (.A(\pcpi_mul.rs2[0] ),
    .X(_03419_));
 sky130_fd_sc_hd__buf_1 _33467_ (.A(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__buf_1 _33468_ (.A(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__buf_1 _33469_ (.A(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__buf_1 _33470_ (.A(_03236_),
    .X(_03423_));
 sky130_fd_sc_hd__buf_1 _33471_ (.A(_18628_),
    .X(_03424_));
 sky130_fd_sc_hd__buf_1 _33472_ (.A(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__buf_1 _33473_ (.A(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__buf_1 _33474_ (.A(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__buf_1 _33475_ (.A(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__buf_1 _33476_ (.A(_03239_),
    .X(_03429_));
 sky130_fd_sc_hd__buf_1 _33477_ (.A(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__buf_1 _33478_ (.A(_03243_),
    .X(_03431_));
 sky130_fd_sc_hd__buf_1 _33479_ (.A(_03431_),
    .X(_03432_));
 sky130_fd_sc_hd__and4_4 _33480_ (.A(_03423_),
    .B(_03428_),
    .C(_03430_),
    .D(_03432_),
    .X(_03433_));
 sky130_fd_sc_hd__a21o_4 _33481_ (.A1(_03418_),
    .A2(_03422_),
    .B1(_03433_),
    .X(_00704_));
 sky130_fd_sc_hd__buf_1 _33482_ (.A(\pcpi_mul.rs2[1] ),
    .X(_03434_));
 sky130_fd_sc_hd__buf_1 _33483_ (.A(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__buf_1 _33484_ (.A(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__buf_1 _33485_ (.A(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__buf_1 _33486_ (.A(_18623_),
    .X(_03438_));
 sky130_fd_sc_hd__buf_1 _33487_ (.A(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__buf_1 _33488_ (.A(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__and4_4 _33489_ (.A(_03423_),
    .B(_03440_),
    .C(_03430_),
    .D(_03432_),
    .X(_03441_));
 sky130_fd_sc_hd__a21o_4 _33490_ (.A1(_03418_),
    .A2(_03437_),
    .B1(_03441_),
    .X(_00715_));
 sky130_fd_sc_hd__buf_1 _33491_ (.A(\pcpi_mul.rs2[2] ),
    .X(_03442_));
 sky130_fd_sc_hd__buf_1 _33492_ (.A(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__buf_1 _33493_ (.A(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__buf_1 _33494_ (.A(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__buf_1 _33495_ (.A(_18614_),
    .X(_03446_));
 sky130_fd_sc_hd__buf_1 _33496_ (.A(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_1 _33497_ (.A(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__buf_1 _33498_ (.A(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__buf_1 _33499_ (.A(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__and4_4 _33500_ (.A(_03423_),
    .B(_03450_),
    .C(_03430_),
    .D(_03432_),
    .X(_03451_));
 sky130_fd_sc_hd__a21o_4 _33501_ (.A1(_03418_),
    .A2(_03445_),
    .B1(_03451_),
    .X(_00726_));
 sky130_fd_sc_hd__buf_1 _33502_ (.A(\pcpi_mul.rs2[3] ),
    .X(_03452_));
 sky130_fd_sc_hd__buf_1 _33503_ (.A(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__buf_1 _33504_ (.A(_03453_),
    .X(_03454_));
 sky130_fd_sc_hd__buf_1 _33505_ (.A(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__buf_1 _33506_ (.A(_03235_),
    .X(_03456_));
 sky130_fd_sc_hd__buf_1 _33507_ (.A(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__buf_1 _33508_ (.A(_18608_),
    .X(_03458_));
 sky130_fd_sc_hd__buf_1 _33509_ (.A(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_1 _33510_ (.A(_03429_),
    .X(_03460_));
 sky130_fd_sc_hd__buf_1 _33511_ (.A(_03431_),
    .X(_03461_));
 sky130_fd_sc_hd__and4_4 _33512_ (.A(_03457_),
    .B(_03459_),
    .C(_03460_),
    .D(_03461_),
    .X(_03462_));
 sky130_fd_sc_hd__a21o_4 _33513_ (.A1(_03418_),
    .A2(_03455_),
    .B1(_03462_),
    .X(_00730_));
 sky130_fd_sc_hd__buf_1 _33514_ (.A(_03412_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_1 _33515_ (.A(\pcpi_mul.rs2[4] ),
    .X(_03464_));
 sky130_fd_sc_hd__buf_1 _33516_ (.A(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__buf_1 _33517_ (.A(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__buf_1 _33518_ (.A(_18602_),
    .X(_03467_));
 sky130_fd_sc_hd__buf_1 _33519_ (.A(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__and4_4 _33520_ (.A(_03457_),
    .B(_03468_),
    .C(_03460_),
    .D(_03461_),
    .X(_03469_));
 sky130_fd_sc_hd__a21o_4 _33521_ (.A1(_03463_),
    .A2(_03466_),
    .B1(_03469_),
    .X(_00731_));
 sky130_fd_sc_hd__buf_1 _33522_ (.A(\pcpi_mul.rs2[5] ),
    .X(_03470_));
 sky130_fd_sc_hd__buf_1 _33523_ (.A(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__buf_1 _33524_ (.A(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__buf_1 _33525_ (.A(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__and4_4 _33526_ (.A(_03457_),
    .B(_18583_),
    .C(_03460_),
    .D(_03461_),
    .X(_03474_));
 sky130_fd_sc_hd__a21o_4 _33527_ (.A1(_03463_),
    .A2(_03473_),
    .B1(_03474_),
    .X(_00732_));
 sky130_fd_sc_hd__buf_1 _33528_ (.A(\pcpi_mul.rs2[6] ),
    .X(_03475_));
 sky130_fd_sc_hd__buf_1 _33529_ (.A(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__buf_1 _33530_ (.A(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__buf_1 _33531_ (.A(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__and4_4 _33532_ (.A(_03457_),
    .B(_18595_),
    .C(_03460_),
    .D(_03461_),
    .X(_03479_));
 sky130_fd_sc_hd__a21o_4 _33533_ (.A1(_03463_),
    .A2(_03478_),
    .B1(_03479_),
    .X(_00733_));
 sky130_fd_sc_hd__buf_1 _33534_ (.A(\pcpi_mul.rs2[7] ),
    .X(_03480_));
 sky130_fd_sc_hd__buf_1 _33535_ (.A(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__buf_1 _33536_ (.A(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__buf_1 _33537_ (.A(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__buf_1 _33538_ (.A(_03456_),
    .X(_03484_));
 sky130_fd_sc_hd__buf_1 _33539_ (.A(_03429_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_1 _33540_ (.A(_03431_),
    .X(_03486_));
 sky130_fd_sc_hd__and4_4 _33541_ (.A(_03484_),
    .B(_18589_),
    .C(_03485_),
    .D(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__a21o_4 _33542_ (.A1(_03463_),
    .A2(_03483_),
    .B1(_03487_),
    .X(_00734_));
 sky130_fd_sc_hd__buf_1 _33543_ (.A(_03411_),
    .X(_03488_));
 sky130_fd_sc_hd__buf_1 _33544_ (.A(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__buf_1 _33545_ (.A(\pcpi_mul.rs2[8] ),
    .X(_03490_));
 sky130_fd_sc_hd__buf_1 _33546_ (.A(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_1 _33547_ (.A(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__buf_1 _33548_ (.A(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__and4_4 _33549_ (.A(_03484_),
    .B(_24236_),
    .C(_03485_),
    .D(_03486_),
    .X(_03494_));
 sky130_fd_sc_hd__a21o_4 _33550_ (.A1(_03489_),
    .A2(_03493_),
    .B1(_03494_),
    .X(_00735_));
 sky130_fd_sc_hd__buf_1 _33551_ (.A(\pcpi_mul.rs2[9] ),
    .X(_03495_));
 sky130_fd_sc_hd__buf_1 _33552_ (.A(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__buf_1 _33553_ (.A(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__and4_4 _33554_ (.A(_03484_),
    .B(_24243_),
    .C(_03485_),
    .D(_03486_),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_4 _33555_ (.A1(_03489_),
    .A2(_03497_),
    .B1(_03498_),
    .X(_00736_));
 sky130_fd_sc_hd__buf_1 _33556_ (.A(\pcpi_mul.rs2[10] ),
    .X(_03499_));
 sky130_fd_sc_hd__buf_1 _33557_ (.A(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__buf_1 _33558_ (.A(_03500_),
    .X(_03501_));
 sky130_vsdinv _33559_ (.A(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__nand4_4 _33560_ (.A(_21228_),
    .B(_03389_),
    .C(_03390_),
    .D(_03391_),
    .Y(_03503_));
 sky130_fd_sc_hd__o21ai_4 _33561_ (.A1(_03502_),
    .A2(_03402_),
    .B1(_03503_),
    .Y(_00705_));
 sky130_fd_sc_hd__buf_1 _33562_ (.A(\pcpi_mul.rs2[11] ),
    .X(_03504_));
 sky130_vsdinv _33563_ (.A(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__buf_1 _33564_ (.A(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__buf_1 _33565_ (.A(_03367_),
    .X(_03507_));
 sky130_fd_sc_hd__buf_1 _33566_ (.A(_03369_),
    .X(_03508_));
 sky130_fd_sc_hd__buf_1 _33567_ (.A(_03371_),
    .X(_03509_));
 sky130_fd_sc_hd__nand4_4 _33568_ (.A(_24248_),
    .B(_03507_),
    .C(_03508_),
    .D(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__o21ai_4 _33569_ (.A1(_03506_),
    .A2(_03402_),
    .B1(_03510_),
    .Y(_00706_));
 sky130_fd_sc_hd__buf_8 _33570_ (.A(\pcpi_mul.rs2[12] ),
    .X(_03511_));
 sky130_fd_sc_hd__buf_1 _33571_ (.A(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__buf_1 _33572_ (.A(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__buf_1 _33573_ (.A(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__and4_4 _33574_ (.A(_03484_),
    .B(_24252_),
    .C(_03485_),
    .D(_03486_),
    .X(_03515_));
 sky130_fd_sc_hd__a21o_4 _33575_ (.A1(_03489_),
    .A2(_03514_),
    .B1(_03515_),
    .X(_00707_));
 sky130_fd_sc_hd__buf_1 _33576_ (.A(\pcpi_mul.rs2[13] ),
    .X(_03516_));
 sky130_fd_sc_hd__buf_1 _33577_ (.A(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__buf_1 _33578_ (.A(_03517_),
    .X(_03518_));
 sky130_fd_sc_hd__buf_1 _33579_ (.A(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__buf_1 _33580_ (.A(_03456_),
    .X(_03520_));
 sky130_fd_sc_hd__buf_1 _33581_ (.A(_03429_),
    .X(_03521_));
 sky130_fd_sc_hd__buf_1 _33582_ (.A(_03431_),
    .X(_03522_));
 sky130_fd_sc_hd__and4_4 _33583_ (.A(_03520_),
    .B(_01476_),
    .C(_03521_),
    .D(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__a21o_4 _33584_ (.A1(_03489_),
    .A2(_03519_),
    .B1(_03523_),
    .X(_00708_));
 sky130_fd_sc_hd__buf_1 _33585_ (.A(\pcpi_mul.rs2[14] ),
    .X(_03524_));
 sky130_fd_sc_hd__buf_1 _33586_ (.A(_03524_),
    .X(_03525_));
 sky130_vsdinv _33587_ (.A(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand4_4 _33588_ (.A(_01478_),
    .B(_03507_),
    .C(_03508_),
    .D(_03509_),
    .Y(_03527_));
 sky130_fd_sc_hd__o21ai_4 _33589_ (.A1(_03526_),
    .A2(_03402_),
    .B1(_03527_),
    .Y(_00709_));
 sky130_fd_sc_hd__buf_1 _33590_ (.A(_03488_),
    .X(_03528_));
 sky130_fd_sc_hd__buf_1 _33591_ (.A(\pcpi_mul.rs2[15] ),
    .X(_03529_));
 sky130_fd_sc_hd__buf_1 _33592_ (.A(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__buf_1 _33593_ (.A(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__buf_1 _33594_ (.A(_03531_),
    .X(_03532_));
 sky130_fd_sc_hd__and4_4 _33595_ (.A(_03520_),
    .B(_01480_),
    .C(_03521_),
    .D(_03522_),
    .X(_03533_));
 sky130_fd_sc_hd__a21o_4 _33596_ (.A1(_03528_),
    .A2(_03532_),
    .B1(_03533_),
    .X(_00710_));
 sky130_fd_sc_hd__buf_1 _33597_ (.A(\pcpi_mul.rs2[16] ),
    .X(_03534_));
 sky130_fd_sc_hd__buf_1 _33598_ (.A(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__buf_1 _33599_ (.A(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__buf_1 _33600_ (.A(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__and4_4 _33601_ (.A(_03520_),
    .B(_18712_),
    .C(_03521_),
    .D(_03522_),
    .X(_03538_));
 sky130_fd_sc_hd__a21o_4 _33602_ (.A1(_03528_),
    .A2(_03537_),
    .B1(_03538_),
    .X(_00711_));
 sky130_fd_sc_hd__buf_1 _33603_ (.A(\pcpi_mul.rs2[17] ),
    .X(_03539_));
 sky130_fd_sc_hd__buf_1 _33604_ (.A(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__buf_1 _33605_ (.A(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__buf_1 _33606_ (.A(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__and4_4 _33607_ (.A(_03520_),
    .B(_18717_),
    .C(_03521_),
    .D(_03522_),
    .X(_03543_));
 sky130_fd_sc_hd__a21o_4 _33608_ (.A1(_03528_),
    .A2(_03542_),
    .B1(_03543_),
    .X(_00712_));
 sky130_fd_sc_hd__buf_1 _33609_ (.A(\pcpi_mul.rs2[18] ),
    .X(_03544_));
 sky130_fd_sc_hd__buf_1 _33610_ (.A(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__buf_1 _33611_ (.A(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__buf_1 _33612_ (.A(_03456_),
    .X(_03547_));
 sky130_fd_sc_hd__buf_1 _33613_ (.A(_03240_),
    .X(_03548_));
 sky130_fd_sc_hd__buf_1 _33614_ (.A(_03244_),
    .X(_03549_));
 sky130_fd_sc_hd__and4_4 _33615_ (.A(_03547_),
    .B(_18706_),
    .C(_03548_),
    .D(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__a21o_4 _33616_ (.A1(_03528_),
    .A2(_03546_),
    .B1(_03550_),
    .X(_00713_));
 sky130_fd_sc_hd__buf_1 _33617_ (.A(\pcpi_mul.rs2[19] ),
    .X(_03551_));
 sky130_fd_sc_hd__buf_1 _33618_ (.A(_03551_),
    .X(_03552_));
 sky130_vsdinv _33619_ (.A(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hd__buf_1 _33620_ (.A(_03234_),
    .X(_03554_));
 sky130_fd_sc_hd__nand4_4 _33621_ (.A(_18696_),
    .B(_03507_),
    .C(_03508_),
    .D(_03509_),
    .Y(_03555_));
 sky130_fd_sc_hd__o21ai_4 _33622_ (.A1(_03553_),
    .A2(_03554_),
    .B1(_03555_),
    .Y(_00714_));
 sky130_fd_sc_hd__buf_1 _33623_ (.A(\pcpi_mul.rs2[20] ),
    .X(_03556_));
 sky130_fd_sc_hd__buf_1 _33624_ (.A(_03556_),
    .X(_03557_));
 sky130_vsdinv _33625_ (.A(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__buf_1 _33626_ (.A(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__nand4_4 _33627_ (.A(_18668_),
    .B(_03507_),
    .C(_03508_),
    .D(_03509_),
    .Y(_03560_));
 sky130_fd_sc_hd__o21ai_4 _33628_ (.A1(_03559_),
    .A2(_03554_),
    .B1(_03560_),
    .Y(_00716_));
 sky130_fd_sc_hd__buf_1 _33629_ (.A(_03488_),
    .X(_03561_));
 sky130_fd_sc_hd__buf_1 _33630_ (.A(\pcpi_mul.rs2[21] ),
    .X(_03562_));
 sky130_fd_sc_hd__buf_1 _33631_ (.A(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__buf_1 _33632_ (.A(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__buf_1 _33633_ (.A(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__buf_1 _33634_ (.A(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__and4_4 _33635_ (.A(_03547_),
    .B(_18682_),
    .C(_03548_),
    .D(_03549_),
    .X(_03567_));
 sky130_fd_sc_hd__a21o_4 _33636_ (.A1(_03561_),
    .A2(_03566_),
    .B1(_03567_),
    .X(_00717_));
 sky130_fd_sc_hd__buf_1 _33637_ (.A(\pcpi_mul.rs2[22] ),
    .X(_03568_));
 sky130_fd_sc_hd__buf_1 _33638_ (.A(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__buf_1 _33639_ (.A(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__buf_1 _33640_ (.A(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__buf_1 _33641_ (.A(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__and4_4 _33642_ (.A(_03547_),
    .B(_18677_),
    .C(_03548_),
    .D(_03549_),
    .X(_03573_));
 sky130_fd_sc_hd__a21o_4 _33643_ (.A1(_03561_),
    .A2(_03572_),
    .B1(_03573_),
    .X(_00718_));
 sky130_fd_sc_hd__buf_1 _33644_ (.A(\pcpi_mul.rs2[23] ),
    .X(_03574_));
 sky130_fd_sc_hd__buf_1 _33645_ (.A(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__buf_1 _33646_ (.A(_03575_),
    .X(_03576_));
 sky130_vsdinv _33647_ (.A(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__buf_1 _33648_ (.A(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nand4_4 _33649_ (.A(_18689_),
    .B(_03423_),
    .C(_03430_),
    .D(_03432_),
    .Y(_03579_));
 sky130_fd_sc_hd__o21ai_4 _33650_ (.A1(_03578_),
    .A2(_03554_),
    .B1(_03579_),
    .Y(_00719_));
 sky130_fd_sc_hd__buf_1 _33651_ (.A(\pcpi_mul.rs2[24] ),
    .X(_03580_));
 sky130_fd_sc_hd__buf_1 _33652_ (.A(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__buf_1 _33653_ (.A(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__buf_1 _33654_ (.A(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__buf_1 _33655_ (.A(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__and4_4 _33656_ (.A(_03547_),
    .B(_18734_),
    .C(_03548_),
    .D(_03549_),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_4 _33657_ (.A1(_03561_),
    .A2(_03584_),
    .B1(_03585_),
    .X(_00720_));
 sky130_fd_sc_hd__buf_1 _33658_ (.A(\pcpi_mul.rs2[25] ),
    .X(_03586_));
 sky130_fd_sc_hd__buf_1 _33659_ (.A(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__buf_1 _33660_ (.A(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__buf_1 _33661_ (.A(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__buf_1 _33662_ (.A(_03236_),
    .X(_03590_));
 sky130_fd_sc_hd__buf_1 _33663_ (.A(_03240_),
    .X(_03591_));
 sky130_fd_sc_hd__buf_1 _33664_ (.A(_03244_),
    .X(_03592_));
 sky130_fd_sc_hd__and4_4 _33665_ (.A(_03590_),
    .B(_18767_),
    .C(_03591_),
    .D(_03592_),
    .X(_03593_));
 sky130_fd_sc_hd__a21o_4 _33666_ (.A1(_03561_),
    .A2(_03589_),
    .B1(_03593_),
    .X(_00721_));
 sky130_fd_sc_hd__buf_1 _33667_ (.A(_03488_),
    .X(_03594_));
 sky130_fd_sc_hd__buf_1 _33668_ (.A(\pcpi_mul.rs2[26] ),
    .X(_03595_));
 sky130_fd_sc_hd__buf_1 _33669_ (.A(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__buf_1 _33670_ (.A(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__buf_1 _33671_ (.A(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__and4_4 _33672_ (.A(_03590_),
    .B(_18722_),
    .C(_03591_),
    .D(_03592_),
    .X(_03599_));
 sky130_fd_sc_hd__a21o_4 _33673_ (.A1(_03594_),
    .A2(_03598_),
    .B1(_03599_),
    .X(_00722_));
 sky130_fd_sc_hd__buf_1 _33674_ (.A(\pcpi_mul.rs2[27] ),
    .X(_03600_));
 sky130_fd_sc_hd__buf_1 _33675_ (.A(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__buf_1 _33676_ (.A(_03601_),
    .X(_03602_));
 sky130_fd_sc_hd__buf_1 _33677_ (.A(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__and4_4 _33678_ (.A(_03590_),
    .B(_18762_),
    .C(_03591_),
    .D(_03592_),
    .X(_03604_));
 sky130_fd_sc_hd__a21o_4 _33679_ (.A1(_03594_),
    .A2(_03603_),
    .B1(_03604_),
    .X(_00723_));
 sky130_fd_sc_hd__buf_8 _33680_ (.A(\pcpi_mul.rs2[28] ),
    .X(_03605_));
 sky130_fd_sc_hd__buf_1 _33681_ (.A(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__buf_4 _33682_ (.A(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__buf_4 _33683_ (.A(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__buf_1 _33684_ (.A(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__buf_1 _33685_ (.A(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__and4_4 _33686_ (.A(_03590_),
    .B(_18747_),
    .C(_03591_),
    .D(_03592_),
    .X(_03611_));
 sky130_fd_sc_hd__a21o_4 _33687_ (.A1(_03594_),
    .A2(_03610_),
    .B1(_03611_),
    .X(_00724_));
 sky130_fd_sc_hd__buf_4 _33688_ (.A(\pcpi_mul.rs2[29] ),
    .X(_03612_));
 sky130_fd_sc_hd__buf_4 _33689_ (.A(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__buf_4 _33690_ (.A(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__buf_4 _33691_ (.A(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__buf_4 _33692_ (.A(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__buf_1 _33693_ (.A(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__and4_4 _33694_ (.A(_03237_),
    .B(_01506_),
    .C(_03241_),
    .D(_03245_),
    .X(_03618_));
 sky130_fd_sc_hd__a21o_4 _33695_ (.A1(_03594_),
    .A2(_03617_),
    .B1(_03618_),
    .X(_00725_));
 sky130_fd_sc_hd__buf_8 _33696_ (.A(\pcpi_mul.rs2[30] ),
    .X(_03619_));
 sky130_fd_sc_hd__buf_8 _33697_ (.A(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_8 _33698_ (.A(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__buf_8 _33699_ (.A(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__buf_1 _33700_ (.A(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__buf_1 _33701_ (.A(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__buf_1 _33702_ (.A(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__and4_4 _33703_ (.A(_03237_),
    .B(_18737_),
    .C(_03241_),
    .D(_03245_),
    .X(_03626_));
 sky130_fd_sc_hd__a21o_4 _33704_ (.A1(_03412_),
    .A2(_03625_),
    .B1(_03626_),
    .X(_00727_));
 sky130_fd_sc_hd__buf_1 _33705_ (.A(\pcpi_mul.rs2[31] ),
    .X(_03627_));
 sky130_fd_sc_hd__buf_1 _33706_ (.A(_03627_),
    .X(_03628_));
 sky130_vsdinv _33707_ (.A(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__and4_4 _33708_ (.A(_03367_),
    .B(_21339_),
    .C(_03369_),
    .D(_03371_),
    .X(_03630_));
 sky130_vsdinv _33709_ (.A(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__o21ai_4 _33710_ (.A1(_03629_),
    .A2(_03554_),
    .B1(_03631_),
    .Y(_00728_));
 sky130_vsdinv _33711_ (.A(\pcpi_mul.rs2[32] ),
    .Y(_03632_));
 sky130_fd_sc_hd__buf_1 _33712_ (.A(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__buf_1 _33713_ (.A(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__buf_1 _33714_ (.A(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_1 _33715_ (.A(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_1 _33716_ (.A(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__nand2_4 _33717_ (.A(_03414_),
    .B(_03630_),
    .Y(_03638_));
 sky130_fd_sc_hd__o21ai_4 _33718_ (.A1(_03637_),
    .A2(_03258_),
    .B1(_03638_),
    .Y(_00729_));
 sky130_fd_sc_hd__nor2_4 _33719_ (.A(_18239_),
    .B(\cpu_state[4] ),
    .Y(_03639_));
 sky130_fd_sc_hd__and2_4 _33720_ (.A(_21225_),
    .B(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_1 _33721_ (.A(_03640_),
    .X(_03641_));
 sky130_vsdinv _33722_ (.A(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__buf_1 _33723_ (.A(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__nand2_4 _33724_ (.A(_21369_),
    .B(mem_rdata[8]),
    .Y(_03644_));
 sky130_fd_sc_hd__buf_1 _33725_ (.A(_21378_),
    .X(_03645_));
 sky130_fd_sc_hd__nand2_4 _33726_ (.A(_03645_),
    .B(mem_rdata[24]),
    .Y(_03646_));
 sky130_fd_sc_hd__nand2_4 _33727_ (.A(_18297_),
    .B(\mem_wordsize[1] ),
    .Y(_03647_));
 sky130_fd_sc_hd__buf_1 _33728_ (.A(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_1 _33729_ (.A(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__a21o_4 _33730_ (.A1(_03644_),
    .A2(_03646_),
    .B1(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__buf_1 _33731_ (.A(_24206_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_1 _33732_ (.A(_21378_),
    .X(_03652_));
 sky130_fd_sc_hd__nand3_4 _33733_ (.A(_03651_),
    .B(_03652_),
    .C(mem_rdata[16]),
    .Y(_03653_));
 sky130_fd_sc_hd__buf_1 _33734_ (.A(_24228_),
    .X(_03654_));
 sky130_fd_sc_hd__a21oi_4 _33735_ (.A1(_03650_),
    .A2(_03653_),
    .B1(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__a21o_4 _33736_ (.A1(mem_rdata[0]),
    .A2(mem_la_wstrb[0]),
    .B1(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__buf_1 _33737_ (.A(_03640_),
    .X(_03657_));
 sky130_fd_sc_hd__buf_1 _33738_ (.A(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_1 _33739_ (.A(_19036_),
    .X(_03659_));
 sky130_fd_sc_hd__nor2_4 _33740_ (.A(_21361_),
    .B(_21345_),
    .Y(_03660_));
 sky130_fd_sc_hd__nand2_4 _33741_ (.A(\reg_pc[0] ),
    .B(\decoded_imm[0] ),
    .Y(_03661_));
 sky130_vsdinv _33742_ (.A(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__nor3_4 _33743_ (.A(_03659_),
    .B(_03660_),
    .C(_03662_),
    .Y(_03663_));
 sky130_vsdinv _33744_ (.A(\pcpi_mul.shift_out ),
    .Y(_03664_));
 sky130_fd_sc_hd__buf_1 _33745_ (.A(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__buf_1 _33746_ (.A(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__buf_1 _33747_ (.A(\pcpi_mul.shift_out ),
    .X(_03667_));
 sky130_fd_sc_hd__buf_1 _33748_ (.A(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__buf_1 _33749_ (.A(_18533_),
    .X(_03669_));
 sky130_fd_sc_hd__buf_1 _33750_ (.A(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__o21a_4 _33751_ (.A1(\pcpi_mul.rd[0] ),
    .A2(_03668_),
    .B1(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__o21a_4 _33752_ (.A1(\pcpi_mul.rd[32] ),
    .A2(_03666_),
    .B1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__a2111oi_4 _33753_ (.A1(_03656_),
    .A2(_18365_),
    .B1(_03658_),
    .C1(_03663_),
    .D1(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__o21ai_4 _33754_ (.A1(_19096_),
    .A2(instr_getq),
    .B1(_19282_),
    .Y(_03674_));
 sky130_fd_sc_hd__buf_1 _33755_ (.A(_18800_),
    .X(_03675_));
 sky130_fd_sc_hd__buf_1 _33756_ (.A(_21058_),
    .X(_03676_));
 sky130_fd_sc_hd__a22oi_4 _33757_ (.A1(_24044_),
    .A2(_19145_),
    .B1(_03676_),
    .B2(\irq_mask[0] ),
    .Y(_03677_));
 sky130_fd_sc_hd__nand3_4 _33758_ (.A(_03674_),
    .B(_03675_),
    .C(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__buf_1 _33759_ (.A(_21061_),
    .X(_03679_));
 sky130_fd_sc_hd__buf_1 _33760_ (.A(_18513_),
    .X(_03680_));
 sky130_fd_sc_hd__buf_1 _33761_ (.A(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__buf_1 _33762_ (.A(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__nand4_4 _33763_ (.A(_24087_),
    .B(_24074_),
    .C(_24095_),
    .D(\count_cycle[0] ),
    .Y(_03683_));
 sky130_fd_sc_hd__buf_1 _33764_ (.A(instr_rdinstrh),
    .X(_03684_));
 sky130_fd_sc_hd__buf_1 _33765_ (.A(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__buf_1 _33766_ (.A(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__nand2_4 _33767_ (.A(_03686_),
    .B(_23251_),
    .Y(_03687_));
 sky130_fd_sc_hd__buf_1 _33768_ (.A(instr_rdinstr),
    .X(_03688_));
 sky130_fd_sc_hd__buf_1 _33769_ (.A(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__buf_1 _33770_ (.A(_03689_),
    .X(_03690_));
 sky130_fd_sc_hd__buf_1 _33771_ (.A(instr_rdcycleh),
    .X(_03691_));
 sky130_fd_sc_hd__buf_1 _33772_ (.A(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__buf_1 _33773_ (.A(\count_cycle[32] ),
    .X(_03693_));
 sky130_fd_sc_hd__a22oi_4 _33774_ (.A1(_03690_),
    .A2(_22999_),
    .B1(_03692_),
    .B2(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__nand4_4 _33775_ (.A(_03682_),
    .B(_03683_),
    .C(_03687_),
    .D(_03694_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand3_4 _33776_ (.A(_03678_),
    .B(_03679_),
    .C(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__a2bb2oi_4 _33777_ (.A1_N(_18907_),
    .A2_N(_03643_),
    .B1(_03673_),
    .B2(_03696_),
    .Y(_24253_));
 sky130_fd_sc_hd__buf_1 _33778_ (.A(_21368_),
    .X(_03697_));
 sky130_fd_sc_hd__nand2_4 _33779_ (.A(_03697_),
    .B(mem_rdata[9]),
    .Y(_03698_));
 sky130_fd_sc_hd__nand2_4 _33780_ (.A(_03645_),
    .B(mem_rdata[25]),
    .Y(_03699_));
 sky130_fd_sc_hd__a21o_4 _33781_ (.A1(_03698_),
    .A2(_03699_),
    .B1(_03649_),
    .X(_03700_));
 sky130_fd_sc_hd__nand3_4 _33782_ (.A(_03651_),
    .B(_03652_),
    .C(mem_rdata[17]),
    .Y(_03701_));
 sky130_fd_sc_hd__a21oi_4 _33783_ (.A1(_03700_),
    .A2(_03701_),
    .B1(_03654_),
    .Y(_03702_));
 sky130_fd_sc_hd__a21o_4 _33784_ (.A1(mem_rdata[1]),
    .A2(mem_la_wstrb[0]),
    .B1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__nor2_4 _33785_ (.A(\reg_pc[1] ),
    .B(_21135_),
    .Y(_03704_));
 sky130_vsdinv _33786_ (.A(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__nand2_4 _33787_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_03706_));
 sky130_fd_sc_hd__a21oi_4 _33788_ (.A1(_03705_),
    .A2(_03706_),
    .B1(_03662_),
    .Y(_03707_));
 sky130_fd_sc_hd__and3_4 _33789_ (.A(_03705_),
    .B(_03662_),
    .C(_03706_),
    .X(_03708_));
 sky130_fd_sc_hd__nor3_4 _33790_ (.A(_03659_),
    .B(_03707_),
    .C(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__buf_1 _33791_ (.A(_03665_),
    .X(_03710_));
 sky130_fd_sc_hd__buf_1 _33792_ (.A(_03667_),
    .X(_03711_));
 sky130_fd_sc_hd__o21a_4 _33793_ (.A1(_03711_),
    .A2(\pcpi_mul.rd[1] ),
    .B1(_03670_),
    .X(_03712_));
 sky130_fd_sc_hd__o21a_4 _33794_ (.A1(_03710_),
    .A2(\pcpi_mul.rd[33] ),
    .B1(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__a2111oi_4 _33795_ (.A1(_03703_),
    .A2(_18838_),
    .B1(_03658_),
    .C1(_03709_),
    .D1(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__nor3_4 _33796_ (.A(_19141_),
    .B(_19096_),
    .C(instr_getq),
    .Y(_03715_));
 sky130_fd_sc_hd__buf_1 _33797_ (.A(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__buf_1 _33798_ (.A(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__a2111o_4 _33799_ (.A1(_19332_),
    .A2(_19379_),
    .B1(_20267_),
    .C1(_19412_),
    .D1(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__a22oi_4 _33800_ (.A1(_24044_),
    .A2(_19422_),
    .B1(_03676_),
    .B2(\irq_mask[1] ),
    .Y(_03719_));
 sky130_fd_sc_hd__nand3_4 _33801_ (.A(_03718_),
    .B(_03675_),
    .C(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__buf_1 _33802_ (.A(_03685_),
    .X(_03721_));
 sky130_fd_sc_hd__buf_1 _33803_ (.A(_18320_),
    .X(_03722_));
 sky130_fd_sc_hd__buf_1 _33804_ (.A(\count_cycle[1] ),
    .X(_03723_));
 sky130_fd_sc_hd__nand4_4 _33805_ (.A(_24086_),
    .B(_24073_),
    .C(_03722_),
    .D(_03723_),
    .Y(_03724_));
 sky130_vsdinv _33806_ (.A(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__buf_1 _33807_ (.A(_03722_),
    .X(_03726_));
 sky130_vsdinv _33808_ (.A(\count_cycle[33] ),
    .Y(_03727_));
 sky130_fd_sc_hd__buf_1 _33809_ (.A(_03689_),
    .X(_03728_));
 sky130_fd_sc_hd__a2bb2o_4 _33810_ (.A1_N(_03726_),
    .A2_N(_03727_),
    .B1(_03728_),
    .B2(\count_instr[1] ),
    .X(_03729_));
 sky130_fd_sc_hd__a2111o_4 _33811_ (.A1(_03721_),
    .A2(_23260_),
    .B1(_03725_),
    .C1(_03729_),
    .D1(_18800_),
    .X(_03730_));
 sky130_fd_sc_hd__nand3_4 _33812_ (.A(_03720_),
    .B(_03679_),
    .C(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__a2bb2oi_4 _33813_ (.A1_N(_18935_),
    .A2_N(_03643_),
    .B1(_03714_),
    .B2(_03731_),
    .Y(_24264_));
 sky130_fd_sc_hd__buf_1 _33814_ (.A(_24209_),
    .X(_03732_));
 sky130_fd_sc_hd__nand2_4 _33815_ (.A(_03697_),
    .B(mem_rdata[10]),
    .Y(_03733_));
 sky130_fd_sc_hd__nand2_4 _33816_ (.A(mem_rdata[26]),
    .B(_24217_),
    .Y(_03734_));
 sky130_fd_sc_hd__a21o_4 _33817_ (.A1(_03733_),
    .A2(_03734_),
    .B1(_03648_),
    .X(_03735_));
 sky130_fd_sc_hd__nand3_4 _33818_ (.A(_03651_),
    .B(_03652_),
    .C(mem_rdata[18]),
    .Y(_03736_));
 sky130_fd_sc_hd__a21oi_4 _33819_ (.A1(_03735_),
    .A2(_03736_),
    .B1(_24229_),
    .Y(_03737_));
 sky130_fd_sc_hd__a21o_4 _33820_ (.A1(mem_rdata[2]),
    .A2(_03732_),
    .B1(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__buf_1 _33821_ (.A(_03657_),
    .X(_03739_));
 sky130_fd_sc_hd__buf_1 _33822_ (.A(_03664_),
    .X(_03740_));
 sky130_fd_sc_hd__buf_1 _33823_ (.A(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__buf_1 _33824_ (.A(\pcpi_mul.shift_out ),
    .X(_03742_));
 sky130_fd_sc_hd__buf_1 _33825_ (.A(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__o21a_4 _33826_ (.A1(_03743_),
    .A2(\pcpi_mul.rd[2] ),
    .B1(_18502_),
    .X(_03744_));
 sky130_fd_sc_hd__o21a_4 _33827_ (.A1(_03741_),
    .A2(\pcpi_mul.rd[34] ),
    .B1(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__nand2_4 _33828_ (.A(\decoded_imm[2] ),
    .B(\reg_pc[2] ),
    .Y(_03746_));
 sky130_vsdinv _33829_ (.A(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__nor2_4 _33830_ (.A(\decoded_imm[2] ),
    .B(\reg_pc[2] ),
    .Y(_03748_));
 sky130_fd_sc_hd__o21a_4 _33831_ (.A1(_03661_),
    .A2(_03704_),
    .B1(_03706_),
    .X(_03749_));
 sky130_fd_sc_hd__o21a_4 _33832_ (.A1(_03747_),
    .A2(_03748_),
    .B1(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__nor3_4 _33833_ (.A(_03747_),
    .B(_03748_),
    .C(_03749_),
    .Y(_03751_));
 sky130_fd_sc_hd__or3_4 _33834_ (.A(_19036_),
    .B(_03750_),
    .C(_03751_),
    .X(_03752_));
 sky130_vsdinv _33835_ (.A(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__a2111oi_4 _33836_ (.A1(_18365_),
    .A2(_03738_),
    .B1(_03739_),
    .C1(_03745_),
    .D1(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__a2111o_4 _33837_ (.A1(_19450_),
    .A2(_19478_),
    .B1(_20267_),
    .C1(_19489_),
    .D1(_03717_),
    .X(_03755_));
 sky130_fd_sc_hd__a22oi_4 _33838_ (.A1(_18311_),
    .A2(_21059_),
    .B1(_24044_),
    .B2(\timer[2] ),
    .Y(_03756_));
 sky130_fd_sc_hd__nand3_4 _33839_ (.A(_03755_),
    .B(_03675_),
    .C(_03756_),
    .Y(_03757_));
 sky130_vsdinv _33840_ (.A(\count_cycle[2] ),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_4 _33841_ (.A(_03685_),
    .B(_23270_),
    .Y(_03759_));
 sky130_fd_sc_hd__buf_1 _33842_ (.A(instr_rdcycleh),
    .X(_03760_));
 sky130_fd_sc_hd__a22oi_4 _33843_ (.A1(_03689_),
    .A2(_23023_),
    .B1(_03760_),
    .B2(\count_cycle[34] ),
    .Y(_03761_));
 sky130_fd_sc_hd__and3_4 _33844_ (.A(_03681_),
    .B(_03759_),
    .C(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__o41ai_4 _33845_ (.A1(_03690_),
    .A2(_03686_),
    .A3(_03692_),
    .A4(_03758_),
    .B1(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand3_4 _33846_ (.A(_03757_),
    .B(_03679_),
    .C(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__a2bb2oi_4 _33847_ (.A1_N(_21991_),
    .A2_N(_03643_),
    .B1(_03754_),
    .B2(_03764_),
    .Y(_24275_));
 sky130_fd_sc_hd__xor2_4 _33848_ (.A(_21159_),
    .B(_21418_),
    .X(_03765_));
 sky130_fd_sc_hd__o21a_4 _33849_ (.A1(_03748_),
    .A2(_03749_),
    .B1(_03746_),
    .X(_03766_));
 sky130_vsdinv _33850_ (.A(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__a21oi_4 _33851_ (.A1(_03767_),
    .A2(_03765_),
    .B1(_19037_),
    .Y(_03768_));
 sky130_fd_sc_hd__o21ai_4 _33852_ (.A1(_03765_),
    .A2(_03767_),
    .B1(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__nand2_4 _33853_ (.A(_21369_),
    .B(mem_rdata[11]),
    .Y(_03770_));
 sky130_fd_sc_hd__nand2_4 _33854_ (.A(mem_rdata[27]),
    .B(_03645_),
    .Y(_03771_));
 sky130_fd_sc_hd__a21o_4 _33855_ (.A1(_03770_),
    .A2(_03771_),
    .B1(_03649_),
    .X(_03772_));
 sky130_fd_sc_hd__nand3_4 _33856_ (.A(_24226_),
    .B(_24218_),
    .C(mem_rdata[19]),
    .Y(_03773_));
 sky130_fd_sc_hd__a21oi_4 _33857_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03654_),
    .Y(_03774_));
 sky130_fd_sc_hd__and2_4 _33858_ (.A(_24209_),
    .B(mem_rdata[3]),
    .X(_03775_));
 sky130_fd_sc_hd__o21ai_4 _33859_ (.A1(_03774_),
    .A2(_03775_),
    .B1(_18838_),
    .Y(_03776_));
 sky130_fd_sc_hd__o21a_4 _33860_ (.A1(_03668_),
    .A2(\pcpi_mul.rd[3] ),
    .B1(_18855_),
    .X(_03777_));
 sky130_fd_sc_hd__o21ai_4 _33861_ (.A1(_03666_),
    .A2(\pcpi_mul.rd[35] ),
    .B1(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__nand4_4 _33862_ (.A(_03642_),
    .B(_03769_),
    .C(_03776_),
    .D(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__buf_1 _33863_ (.A(_03715_),
    .X(_03780_));
 sky130_fd_sc_hd__a2111o_4 _33864_ (.A1(_19523_),
    .A2(_19551_),
    .B1(_21519_),
    .C1(_19562_),
    .D1(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__buf_1 _33865_ (.A(_18515_),
    .X(_03782_));
 sky130_fd_sc_hd__a22oi_4 _33866_ (.A1(_24043_),
    .A2(\timer[3] ),
    .B1(_21058_),
    .B2(\irq_mask[3] ),
    .Y(_03783_));
 sky130_fd_sc_hd__nand3_4 _33867_ (.A(_03781_),
    .B(_03782_),
    .C(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__buf_1 _33868_ (.A(_03760_),
    .X(_03785_));
 sky130_vsdinv _33869_ (.A(\count_cycle[3] ),
    .Y(_03786_));
 sky130_fd_sc_hd__buf_1 _33870_ (.A(_03684_),
    .X(_03787_));
 sky130_fd_sc_hd__nand2_4 _33871_ (.A(_03787_),
    .B(\count_instr[35] ),
    .Y(_03788_));
 sky130_fd_sc_hd__a22oi_4 _33872_ (.A1(_03688_),
    .A2(\count_instr[3] ),
    .B1(_03760_),
    .B2(\count_cycle[35] ),
    .Y(_03789_));
 sky130_fd_sc_hd__and3_4 _33873_ (.A(_03680_),
    .B(_03788_),
    .C(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__o41ai_4 _33874_ (.A1(_03728_),
    .A2(_03721_),
    .A3(_03785_),
    .A4(_03786_),
    .B1(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__and3_4 _33875_ (.A(_03784_),
    .B(_20232_),
    .C(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__o22a_4 _33876_ (.A1(_18946_),
    .A2(_03642_),
    .B1(_03779_),
    .B2(_03792_),
    .X(_24278_));
 sky130_fd_sc_hd__buf_1 _33877_ (.A(_03739_),
    .X(_03793_));
 sky130_fd_sc_hd__a2111o_4 _33878_ (.A1(_19604_),
    .A2(_19629_),
    .B1(_20267_),
    .C1(_19648_),
    .D1(_03717_),
    .X(_03794_));
 sky130_fd_sc_hd__buf_1 _33879_ (.A(_24043_),
    .X(_03795_));
 sky130_fd_sc_hd__a22oi_4 _33880_ (.A1(_03795_),
    .A2(\timer[4] ),
    .B1(_03676_),
    .B2(\irq_mask[4] ),
    .Y(_03796_));
 sky130_fd_sc_hd__nand3_4 _33881_ (.A(_03794_),
    .B(_03675_),
    .C(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__nand4_4 _33882_ (.A(_24087_),
    .B(_24074_),
    .C(_24095_),
    .D(\count_cycle[4] ),
    .Y(_03798_));
 sky130_fd_sc_hd__nand2_4 _33883_ (.A(_03686_),
    .B(_23289_),
    .Y(_03799_));
 sky130_fd_sc_hd__a22oi_4 _33884_ (.A1(_03690_),
    .A2(_23037_),
    .B1(_03692_),
    .B2(\count_cycle[36] ),
    .Y(_03800_));
 sky130_fd_sc_hd__nand4_4 _33885_ (.A(_03682_),
    .B(_03798_),
    .C(_03799_),
    .D(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__nand3_4 _33886_ (.A(_03797_),
    .B(_03679_),
    .C(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_4 _33887_ (.A(\decoded_imm[4] ),
    .B(\reg_pc[4] ),
    .Y(_03803_));
 sky130_fd_sc_hd__nor2_4 _33888_ (.A(\decoded_imm[4] ),
    .B(\reg_pc[4] ),
    .Y(_03804_));
 sky130_vsdinv _33889_ (.A(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__nor2_4 _33890_ (.A(\decoded_imm[3] ),
    .B(\reg_pc[3] ),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_4 _33891_ (.A(\decoded_imm[3] ),
    .B(\reg_pc[3] ),
    .Y(_03807_));
 sky130_fd_sc_hd__o21ai_4 _33892_ (.A1(_03806_),
    .A2(_03766_),
    .B1(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__a21o_4 _33893_ (.A1(_03803_),
    .A2(_03805_),
    .B1(_03808_),
    .X(_03809_));
 sky130_vsdinv _33894_ (.A(_03803_),
    .Y(_03810_));
 sky130_fd_sc_hd__nor2_4 _33895_ (.A(_03804_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__a21oi_4 _33896_ (.A1(_03808_),
    .A2(_03811_),
    .B1(_03659_),
    .Y(_03812_));
 sky130_fd_sc_hd__buf_1 _33897_ (.A(_03657_),
    .X(_03813_));
 sky130_fd_sc_hd__nand2_4 _33898_ (.A(_21368_),
    .B(mem_rdata[12]),
    .Y(_03814_));
 sky130_fd_sc_hd__nand2_4 _33899_ (.A(_24217_),
    .B(mem_rdata[28]),
    .Y(_03815_));
 sky130_fd_sc_hd__a21o_4 _33900_ (.A1(_03814_),
    .A2(_03815_),
    .B1(_03648_),
    .X(_03816_));
 sky130_fd_sc_hd__nand3_4 _33901_ (.A(_24226_),
    .B(_24218_),
    .C(mem_rdata[20]),
    .Y(_03817_));
 sky130_fd_sc_hd__a21o_4 _33902_ (.A1(_03816_),
    .A2(_03817_),
    .B1(_24229_),
    .X(_03818_));
 sky130_fd_sc_hd__nand2_4 _33903_ (.A(_03732_),
    .B(mem_rdata[4]),
    .Y(_03819_));
 sky130_fd_sc_hd__buf_1 _33904_ (.A(_18270_),
    .X(_03820_));
 sky130_fd_sc_hd__a21oi_4 _33905_ (.A1(_03818_),
    .A2(_03819_),
    .B1(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__buf_1 _33906_ (.A(_03669_),
    .X(_03822_));
 sky130_fd_sc_hd__o21a_4 _33907_ (.A1(_03711_),
    .A2(\pcpi_mul.rd[4] ),
    .B1(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__o21a_4 _33908_ (.A1(_03710_),
    .A2(\pcpi_mul.rd[36] ),
    .B1(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__a2111oi_4 _33909_ (.A1(_03809_),
    .A2(_03812_),
    .B1(_03813_),
    .C1(_03821_),
    .D1(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__a22oi_4 _33910_ (.A1(_21993_),
    .A2(_03793_),
    .B1(_03802_),
    .B2(_03825_),
    .Y(_24279_));
 sky130_fd_sc_hd__a2111o_4 _33911_ (.A1(_19671_),
    .A2(_19686_),
    .B1(_19194_),
    .C1(_19693_),
    .D1(_03717_),
    .X(_03826_));
 sky130_fd_sc_hd__buf_1 _33912_ (.A(_18800_),
    .X(_03827_));
 sky130_fd_sc_hd__a22oi_4 _33913_ (.A1(_03795_),
    .A2(\timer[5] ),
    .B1(_03676_),
    .B2(\irq_mask[5] ),
    .Y(_03828_));
 sky130_fd_sc_hd__nand3_4 _33914_ (.A(_03826_),
    .B(_03827_),
    .C(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__buf_1 _33915_ (.A(\count_cycle[5] ),
    .X(_03830_));
 sky130_fd_sc_hd__nand4_4 _33916_ (.A(_24087_),
    .B(_24074_),
    .C(_24095_),
    .D(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_4 _33917_ (.A(_03686_),
    .B(_23292_),
    .Y(_03832_));
 sky130_fd_sc_hd__a22oi_4 _33918_ (.A1(_03690_),
    .A2(\count_instr[5] ),
    .B1(_03692_),
    .B2(\count_cycle[37] ),
    .Y(_03833_));
 sky130_fd_sc_hd__nand4_4 _33919_ (.A(_03682_),
    .B(_03831_),
    .C(_03832_),
    .D(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand3_4 _33920_ (.A(_03829_),
    .B(_21583_),
    .C(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__a21oi_4 _33921_ (.A1(_03808_),
    .A2(_03805_),
    .B1(_03810_),
    .Y(_03836_));
 sky130_vsdinv _33922_ (.A(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__xor2_4 _33923_ (.A(_21186_),
    .B(_21458_),
    .X(_03838_));
 sky130_fd_sc_hd__a21oi_4 _33924_ (.A1(_03837_),
    .A2(_03838_),
    .B1(_03659_),
    .Y(_03839_));
 sky130_fd_sc_hd__a211o_4 _33925_ (.A1(_03808_),
    .A2(_03805_),
    .B1(_03810_),
    .C1(_03838_),
    .X(_03840_));
 sky130_fd_sc_hd__nand2_4 _33926_ (.A(_21368_),
    .B(mem_rdata[13]),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2_4 _33927_ (.A(_24217_),
    .B(mem_rdata[29]),
    .Y(_03842_));
 sky130_fd_sc_hd__a21o_4 _33928_ (.A1(_03841_),
    .A2(_03842_),
    .B1(_03648_),
    .X(_03843_));
 sky130_fd_sc_hd__buf_1 _33929_ (.A(_21378_),
    .X(_03844_));
 sky130_fd_sc_hd__nand3_4 _33930_ (.A(_03651_),
    .B(_03844_),
    .C(mem_rdata[21]),
    .Y(_03845_));
 sky130_fd_sc_hd__a21o_4 _33931_ (.A1(_03843_),
    .A2(_03845_),
    .B1(_24229_),
    .X(_03846_));
 sky130_fd_sc_hd__nand2_4 _33932_ (.A(_03732_),
    .B(mem_rdata[5]),
    .Y(_03847_));
 sky130_fd_sc_hd__a21oi_4 _33933_ (.A1(_03846_),
    .A2(_03847_),
    .B1(_03820_),
    .Y(_03848_));
 sky130_fd_sc_hd__o21a_4 _33934_ (.A1(_03711_),
    .A2(\pcpi_mul.rd[5] ),
    .B1(_03822_),
    .X(_03849_));
 sky130_fd_sc_hd__o21a_4 _33935_ (.A1(_03710_),
    .A2(\pcpi_mul.rd[37] ),
    .B1(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__a2111oi_4 _33936_ (.A1(_03839_),
    .A2(_03840_),
    .B1(_03813_),
    .C1(_03848_),
    .D1(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__a22oi_4 _33937_ (.A1(_21994_),
    .A2(_03793_),
    .B1(_03835_),
    .B2(_03851_),
    .Y(_24280_));
 sky130_fd_sc_hd__buf_1 _33938_ (.A(_03716_),
    .X(_03852_));
 sky130_fd_sc_hd__a2111o_4 _33939_ (.A1(_19719_),
    .A2(_19738_),
    .B1(_20874_),
    .C1(_19749_),
    .D1(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__a22oi_4 _33940_ (.A1(_03795_),
    .A2(\timer[6] ),
    .B1(_21059_),
    .B2(\irq_mask[6] ),
    .Y(_03854_));
 sky130_fd_sc_hd__nand3_4 _33941_ (.A(_03853_),
    .B(_03827_),
    .C(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__buf_1 _33942_ (.A(_24085_),
    .X(_03856_));
 sky130_fd_sc_hd__buf_1 _33943_ (.A(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__buf_1 _33944_ (.A(_24072_),
    .X(_03858_));
 sky130_fd_sc_hd__buf_1 _33945_ (.A(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_1 _33946_ (.A(_03722_),
    .X(_03860_));
 sky130_fd_sc_hd__nand4_4 _33947_ (.A(_03857_),
    .B(_03859_),
    .C(_03860_),
    .D(\count_cycle[6] ),
    .Y(_03861_));
 sky130_fd_sc_hd__nand2_4 _33948_ (.A(_03721_),
    .B(\count_instr[38] ),
    .Y(_03862_));
 sky130_fd_sc_hd__buf_1 _33949_ (.A(\count_cycle[38] ),
    .X(_03863_));
 sky130_fd_sc_hd__a22oi_4 _33950_ (.A1(_03728_),
    .A2(\count_instr[6] ),
    .B1(_03785_),
    .B2(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__a41oi_4 _33951_ (.A1(_03682_),
    .A2(_03861_),
    .A3(_03862_),
    .A4(_03864_),
    .B1(_21116_),
    .Y(_03865_));
 sky130_fd_sc_hd__buf_1 _33952_ (.A(_03640_),
    .X(_03866_));
 sky130_fd_sc_hd__buf_1 _33953_ (.A(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__nand2_4 _33954_ (.A(_03697_),
    .B(mem_rdata[14]),
    .Y(_03868_));
 sky130_fd_sc_hd__nand2_4 _33955_ (.A(_03645_),
    .B(mem_rdata[30]),
    .Y(_03869_));
 sky130_fd_sc_hd__a21o_4 _33956_ (.A1(_03868_),
    .A2(_03869_),
    .B1(_03649_),
    .X(_03870_));
 sky130_fd_sc_hd__nand3_4 _33957_ (.A(_24226_),
    .B(_24218_),
    .C(mem_rdata[22]),
    .Y(_03871_));
 sky130_fd_sc_hd__a21o_4 _33958_ (.A1(_03870_),
    .A2(_03871_),
    .B1(_03654_),
    .X(_03872_));
 sky130_fd_sc_hd__nand2_4 _33959_ (.A(_03732_),
    .B(mem_rdata[6]),
    .Y(_03873_));
 sky130_fd_sc_hd__buf_1 _33960_ (.A(_18270_),
    .X(_03874_));
 sky130_fd_sc_hd__a21oi_4 _33961_ (.A1(_03872_),
    .A2(_03873_),
    .B1(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__buf_1 _33962_ (.A(_18534_),
    .X(_03876_));
 sky130_fd_sc_hd__o21a_4 _33963_ (.A1(_03668_),
    .A2(\pcpi_mul.rd[6] ),
    .B1(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__o21a_4 _33964_ (.A1(_03666_),
    .A2(\pcpi_mul.rd[38] ),
    .B1(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__a2111oi_4 _33965_ (.A1(_03855_),
    .A2(_03865_),
    .B1(_03867_),
    .C1(_03875_),
    .D1(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__xor2_4 _33966_ (.A(\decoded_imm[6] ),
    .B(\reg_pc[6] ),
    .X(_03880_));
 sky130_fd_sc_hd__nor2_4 _33967_ (.A(\decoded_imm[5] ),
    .B(\reg_pc[5] ),
    .Y(_03881_));
 sky130_fd_sc_hd__nand2_4 _33968_ (.A(\decoded_imm[5] ),
    .B(_21457_),
    .Y(_03882_));
 sky130_fd_sc_hd__o21ai_4 _33969_ (.A1(_03881_),
    .A2(_03836_),
    .B1(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__or2_4 _33970_ (.A(_03880_),
    .B(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__buf_1 _33971_ (.A(_18400_),
    .X(_03885_));
 sky130_fd_sc_hd__nand2_4 _33972_ (.A(_03883_),
    .B(_03880_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand3_4 _33973_ (.A(_03884_),
    .B(_03885_),
    .C(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__a22oi_4 _33974_ (.A1(_21995_),
    .A2(_03793_),
    .B1(_03879_),
    .B2(_03887_),
    .Y(_24281_));
 sky130_fd_sc_hd__a2111o_4 _33975_ (.A1(_19770_),
    .A2(_19785_),
    .B1(_20874_),
    .C1(_19797_),
    .D1(_03852_),
    .X(_03888_));
 sky130_fd_sc_hd__a22oi_4 _33976_ (.A1(_03795_),
    .A2(\timer[7] ),
    .B1(_21059_),
    .B2(\irq_mask[7] ),
    .Y(_03889_));
 sky130_fd_sc_hd__nand3_4 _33977_ (.A(_03888_),
    .B(_03827_),
    .C(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__buf_1 _33978_ (.A(_03681_),
    .X(_03891_));
 sky130_fd_sc_hd__nand4_4 _33979_ (.A(_03857_),
    .B(_03859_),
    .C(_03860_),
    .D(\count_cycle[7] ),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_4 _33980_ (.A(_03721_),
    .B(\count_instr[39] ),
    .Y(_03893_));
 sky130_fd_sc_hd__a22oi_4 _33981_ (.A1(_03728_),
    .A2(\count_instr[7] ),
    .B1(_03785_),
    .B2(\count_cycle[39] ),
    .Y(_03894_));
 sky130_fd_sc_hd__a41oi_4 _33982_ (.A1(_03891_),
    .A2(_03892_),
    .A3(_03893_),
    .A4(_03894_),
    .B1(_21116_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_4 _33983_ (.A(_21367_),
    .B(mem_rdata[15]),
    .Y(_03896_));
 sky130_fd_sc_hd__nand2_4 _33984_ (.A(pcpi_rs1[1]),
    .B(mem_rdata[31]),
    .Y(_03897_));
 sky130_fd_sc_hd__a21o_4 _33985_ (.A1(_03896_),
    .A2(_03897_),
    .B1(_03647_),
    .X(_03898_));
 sky130_fd_sc_hd__nand3_4 _33986_ (.A(_24206_),
    .B(_18301_),
    .C(mem_rdata[23]),
    .Y(_03899_));
 sky130_fd_sc_hd__a21oi_4 _33987_ (.A1(_03898_),
    .A2(_03899_),
    .B1(_24207_),
    .Y(_03900_));
 sky130_fd_sc_hd__a21oi_4 _33988_ (.A1(mem_rdata[7]),
    .A2(_24209_),
    .B1(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__nor2_4 _33989_ (.A(_03874_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__o21a_4 _33990_ (.A1(_03668_),
    .A2(\pcpi_mul.rd[7] ),
    .B1(_03876_),
    .X(_03903_));
 sky130_fd_sc_hd__o21a_4 _33991_ (.A1(_03666_),
    .A2(\pcpi_mul.rd[39] ),
    .B1(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__a2111oi_4 _33992_ (.A1(_03890_),
    .A2(_03895_),
    .B1(_03867_),
    .C1(_03902_),
    .D1(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__xor2_4 _33993_ (.A(_21201_),
    .B(_21490_),
    .X(_03906_));
 sky130_vsdinv _33994_ (.A(_03886_),
    .Y(_03907_));
 sky130_fd_sc_hd__a211o_4 _33995_ (.A1(_21193_),
    .A2(_21476_),
    .B1(_03906_),
    .C1(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__nand2_4 _33996_ (.A(_21193_),
    .B(_21476_),
    .Y(_03909_));
 sky130_fd_sc_hd__a21bo_4 _33997_ (.A1(_03886_),
    .A2(_03909_),
    .B1_N(_03906_),
    .X(_03910_));
 sky130_fd_sc_hd__nand3_4 _33998_ (.A(_03908_),
    .B(_03885_),
    .C(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__a22oi_4 _33999_ (.A1(_21996_),
    .A2(_03793_),
    .B1(_03905_),
    .B2(_03911_),
    .Y(_24282_));
 sky130_fd_sc_hd__buf_1 _34000_ (.A(_03739_),
    .X(_03912_));
 sky130_fd_sc_hd__a2111o_4 _34001_ (.A1(_19829_),
    .A2(_19853_),
    .B1(_20874_),
    .C1(_19862_),
    .D1(_03852_),
    .X(_03913_));
 sky130_fd_sc_hd__buf_1 _34002_ (.A(_24043_),
    .X(_03914_));
 sky130_fd_sc_hd__buf_1 _34003_ (.A(_21058_),
    .X(_03915_));
 sky130_fd_sc_hd__a22oi_4 _34004_ (.A1(_03914_),
    .A2(\timer[8] ),
    .B1(_03915_),
    .B2(\irq_mask[8] ),
    .Y(_03916_));
 sky130_fd_sc_hd__nand3_4 _34005_ (.A(_03913_),
    .B(_03827_),
    .C(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__buf_1 _34006_ (.A(\count_cycle[8] ),
    .X(_03918_));
 sky130_fd_sc_hd__nand4_4 _34007_ (.A(_03857_),
    .B(_03859_),
    .C(_03860_),
    .D(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__buf_1 _34008_ (.A(_03685_),
    .X(_03920_));
 sky130_fd_sc_hd__nand2_4 _34009_ (.A(_03920_),
    .B(\count_instr[40] ),
    .Y(_03921_));
 sky130_fd_sc_hd__buf_1 _34010_ (.A(_03689_),
    .X(_03922_));
 sky130_fd_sc_hd__a22oi_4 _34011_ (.A1(_03922_),
    .A2(_23073_),
    .B1(_03785_),
    .B2(\count_cycle[40] ),
    .Y(_03923_));
 sky130_fd_sc_hd__a41oi_4 _34012_ (.A1(_03891_),
    .A2(_03919_),
    .A3(_03921_),
    .A4(_03923_),
    .B1(_21116_),
    .Y(_03924_));
 sky130_vsdinv _34013_ (.A(latched_is_lb),
    .Y(_03925_));
 sky130_fd_sc_hd__or2_4 _34014_ (.A(_03925_),
    .B(_03901_),
    .X(_03926_));
 sky130_fd_sc_hd__buf_1 _34015_ (.A(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__buf_1 _34016_ (.A(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__nor2_4 _34017_ (.A(_18619_),
    .B(_01484_),
    .Y(_03929_));
 sky130_fd_sc_hd__buf_1 _34018_ (.A(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__buf_1 _34019_ (.A(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__o21ai_4 _34020_ (.A1(_01503_),
    .A2(_03931_),
    .B1(mem_rdata[8]),
    .Y(_03932_));
 sky130_fd_sc_hd__nand3_4 _34021_ (.A(_01481_),
    .B(_03844_),
    .C(mem_rdata[24]),
    .Y(_03933_));
 sky130_fd_sc_hd__nor2_4 _34022_ (.A(latched_is_lh),
    .B(_03925_),
    .Y(_03934_));
 sky130_fd_sc_hd__buf_1 _34023_ (.A(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__a21o_4 _34024_ (.A1(_03932_),
    .A2(_03933_),
    .B1(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__buf_1 _34025_ (.A(_18362_),
    .X(_03937_));
 sky130_fd_sc_hd__a21oi_4 _34026_ (.A1(_03928_),
    .A2(_03936_),
    .B1(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__buf_1 _34027_ (.A(_03665_),
    .X(_03939_));
 sky130_fd_sc_hd__buf_1 _34028_ (.A(_03667_),
    .X(_03940_));
 sky130_fd_sc_hd__o21a_4 _34029_ (.A1(_03940_),
    .A2(\pcpi_mul.rd[8] ),
    .B1(_03876_),
    .X(_03941_));
 sky130_fd_sc_hd__o21a_4 _34030_ (.A1(_03939_),
    .A2(\pcpi_mul.rd[40] ),
    .B1(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__a2111oi_4 _34031_ (.A1(_03917_),
    .A2(_03924_),
    .B1(_03867_),
    .C1(_03938_),
    .D1(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__a22oi_4 _34032_ (.A1(\decoded_imm[6] ),
    .A2(\reg_pc[6] ),
    .B1(\decoded_imm[7] ),
    .B2(\reg_pc[7] ),
    .Y(_03944_));
 sky130_fd_sc_hd__nand2_4 _34033_ (.A(_03886_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__nor2_4 _34034_ (.A(_21200_),
    .B(\reg_pc[7] ),
    .Y(_03946_));
 sky130_vsdinv _34035_ (.A(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__xor2_4 _34036_ (.A(\decoded_imm[8] ),
    .B(\reg_pc[8] ),
    .X(_03948_));
 sky130_fd_sc_hd__a21o_4 _34037_ (.A1(_03945_),
    .A2(_03947_),
    .B1(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__nand3_4 _34038_ (.A(_03945_),
    .B(_03947_),
    .C(_03948_),
    .Y(_03950_));
 sky130_fd_sc_hd__nand3_4 _34039_ (.A(_03949_),
    .B(_18866_),
    .C(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__a22oi_4 _34040_ (.A1(_22026_),
    .A2(_03912_),
    .B1(_03943_),
    .B2(_03951_),
    .Y(_24283_));
 sky130_fd_sc_hd__a2111o_4 _34041_ (.A1(_19888_),
    .A2(_19907_),
    .B1(_20156_),
    .C1(_19919_),
    .D1(_03852_),
    .X(_03952_));
 sky130_fd_sc_hd__buf_1 _34042_ (.A(_18514_),
    .X(_03953_));
 sky130_fd_sc_hd__buf_1 _34043_ (.A(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__a22oi_4 _34044_ (.A1(_03914_),
    .A2(\timer[9] ),
    .B1(_03915_),
    .B2(\irq_mask[9] ),
    .Y(_03955_));
 sky130_fd_sc_hd__nand3_4 _34045_ (.A(_03952_),
    .B(_03954_),
    .C(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__buf_1 _34046_ (.A(\count_cycle[9] ),
    .X(_03957_));
 sky130_fd_sc_hd__nand4_4 _34047_ (.A(_03857_),
    .B(_03859_),
    .C(_03860_),
    .D(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__nand2_4 _34048_ (.A(_03920_),
    .B(_23317_),
    .Y(_03959_));
 sky130_fd_sc_hd__buf_1 _34049_ (.A(_03760_),
    .X(_03960_));
 sky130_fd_sc_hd__a22oi_4 _34050_ (.A1(_03922_),
    .A2(\count_instr[9] ),
    .B1(_03960_),
    .B2(\count_cycle[41] ),
    .Y(_03961_));
 sky130_fd_sc_hd__buf_1 _34051_ (.A(_21133_),
    .X(_03962_));
 sky130_fd_sc_hd__a41oi_4 _34052_ (.A1(_03891_),
    .A2(_03958_),
    .A3(_03959_),
    .A4(_03961_),
    .B1(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__o21ai_4 _34053_ (.A1(_01503_),
    .A2(_03931_),
    .B1(mem_rdata[9]),
    .Y(_03964_));
 sky130_fd_sc_hd__nand3_4 _34054_ (.A(_01481_),
    .B(_03844_),
    .C(mem_rdata[25]),
    .Y(_03965_));
 sky130_fd_sc_hd__a21o_4 _34055_ (.A1(_03964_),
    .A2(_03965_),
    .B1(_03935_),
    .X(_03966_));
 sky130_fd_sc_hd__a21oi_4 _34056_ (.A1(_03928_),
    .A2(_03966_),
    .B1(_03937_),
    .Y(_03967_));
 sky130_fd_sc_hd__o21a_4 _34057_ (.A1(_03940_),
    .A2(\pcpi_mul.rd[9] ),
    .B1(_03876_),
    .X(_03968_));
 sky130_fd_sc_hd__o21a_4 _34058_ (.A1(_03939_),
    .A2(\pcpi_mul.rd[41] ),
    .B1(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__a2111oi_4 _34059_ (.A1(_03956_),
    .A2(_03963_),
    .B1(_03867_),
    .C1(_03967_),
    .D1(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__xor2_4 _34060_ (.A(\decoded_imm[9] ),
    .B(\reg_pc[9] ),
    .X(_03971_));
 sky130_vsdinv _34061_ (.A(_03971_),
    .Y(_03972_));
 sky130_fd_sc_hd__nand2_4 _34062_ (.A(_21206_),
    .B(\reg_pc[8] ),
    .Y(_03973_));
 sky130_fd_sc_hd__a21bo_4 _34063_ (.A1(_03945_),
    .A2(_03947_),
    .B1_N(_03973_),
    .X(_03974_));
 sky130_fd_sc_hd__o21ai_4 _34064_ (.A1(_21207_),
    .A2(_21523_),
    .B1(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__a21oi_4 _34065_ (.A1(_03975_),
    .A2(_03972_),
    .B1(_19038_),
    .Y(_03976_));
 sky130_fd_sc_hd__o21ai_4 _34066_ (.A1(_03972_),
    .A2(_03975_),
    .B1(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__a22oi_4 _34067_ (.A1(_22027_),
    .A2(_03912_),
    .B1(_03970_),
    .B2(_03977_),
    .Y(_24284_));
 sky130_fd_sc_hd__a21o_4 _34068_ (.A1(_24050_),
    .A2(_18511_),
    .B1(_19975_),
    .X(_03978_));
 sky130_fd_sc_hd__a22oi_4 _34069_ (.A1(_03914_),
    .A2(\timer[10] ),
    .B1(_03915_),
    .B2(\irq_mask[10] ),
    .Y(_03979_));
 sky130_fd_sc_hd__nand3_4 _34070_ (.A(_03978_),
    .B(_03954_),
    .C(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__buf_1 _34071_ (.A(_03856_),
    .X(_03981_));
 sky130_fd_sc_hd__buf_1 _34072_ (.A(_03858_),
    .X(_03982_));
 sky130_fd_sc_hd__buf_1 _34073_ (.A(\count_cycle[10] ),
    .X(_03983_));
 sky130_fd_sc_hd__nand4_4 _34074_ (.A(_03981_),
    .B(_03982_),
    .C(_03726_),
    .D(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_4 _34075_ (.A(_03920_),
    .B(_23324_),
    .Y(_03985_));
 sky130_fd_sc_hd__buf_1 _34076_ (.A(\count_cycle[42] ),
    .X(_03986_));
 sky130_fd_sc_hd__a22oi_4 _34077_ (.A1(_03922_),
    .A2(\count_instr[10] ),
    .B1(_03960_),
    .B2(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__a41oi_4 _34078_ (.A1(_03891_),
    .A2(_03984_),
    .A3(_03985_),
    .A4(_03987_),
    .B1(_03962_),
    .Y(_03988_));
 sky130_fd_sc_hd__buf_1 _34079_ (.A(_24227_),
    .X(_03989_));
 sky130_fd_sc_hd__o21ai_4 _34080_ (.A1(_03989_),
    .A2(_03931_),
    .B1(mem_rdata[10]),
    .Y(_03990_));
 sky130_fd_sc_hd__nand3_4 _34081_ (.A(mem_rdata[26]),
    .B(_24219_),
    .C(_03652_),
    .Y(_03991_));
 sky130_fd_sc_hd__a21o_4 _34082_ (.A1(_03990_),
    .A2(_03991_),
    .B1(_03935_),
    .X(_03992_));
 sky130_fd_sc_hd__a21oi_4 _34083_ (.A1(_03928_),
    .A2(_03992_),
    .B1(_03937_),
    .Y(_03993_));
 sky130_fd_sc_hd__o21a_4 _34084_ (.A1(_03940_),
    .A2(\pcpi_mul.rd[10] ),
    .B1(_03670_),
    .X(_03994_));
 sky130_fd_sc_hd__o21a_4 _34085_ (.A1(_03939_),
    .A2(\pcpi_mul.rd[42] ),
    .B1(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__a2111oi_4 _34086_ (.A1(_03980_),
    .A2(_03988_),
    .B1(_03658_),
    .C1(_03993_),
    .D1(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__xor2_4 _34087_ (.A(\decoded_imm[10] ),
    .B(\reg_pc[10] ),
    .X(_03997_));
 sky130_fd_sc_hd__nand4_4 _34088_ (.A(_03947_),
    .B(_03945_),
    .C(_03948_),
    .D(_03971_),
    .Y(_03998_));
 sky130_vsdinv _34089_ (.A(\reg_pc[9] ),
    .Y(_03999_));
 sky130_fd_sc_hd__maj3_4 _34090_ (.A(_21218_),
    .B(_03973_),
    .C(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__nand2_4 _34091_ (.A(_03998_),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__buf_1 _34092_ (.A(_19037_),
    .X(_04002_));
 sky130_fd_sc_hd__a21oi_4 _34093_ (.A1(_04001_),
    .A2(_03997_),
    .B1(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__o21ai_4 _34094_ (.A1(_03997_),
    .A2(_04001_),
    .B1(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__a22oi_4 _34095_ (.A1(_22028_),
    .A2(_03912_),
    .B1(_03996_),
    .B2(_04004_),
    .Y(_24254_));
 sky130_fd_sc_hd__xor2_4 _34096_ (.A(\decoded_imm[11] ),
    .B(\reg_pc[11] ),
    .X(_04005_));
 sky130_fd_sc_hd__maj3_4 _34097_ (.A(_21222_),
    .B(_04001_),
    .C(_21559_),
    .X(_04006_));
 sky130_fd_sc_hd__o21ai_4 _34098_ (.A1(_04005_),
    .A2(_04006_),
    .B1(_18866_),
    .Y(_04007_));
 sky130_fd_sc_hd__a21o_4 _34099_ (.A1(_04005_),
    .A2(_04006_),
    .B1(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__buf_1 _34100_ (.A(_03716_),
    .X(_04009_));
 sky130_fd_sc_hd__a2111o_4 _34101_ (.A1(_20004_),
    .A2(_20028_),
    .B1(_20649_),
    .C1(_20049_),
    .D1(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__buf_1 _34102_ (.A(_19163_),
    .X(_04011_));
 sky130_fd_sc_hd__buf_1 _34103_ (.A(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__buf_1 _34104_ (.A(_21016_),
    .X(_04013_));
 sky130_fd_sc_hd__buf_1 _34105_ (.A(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__a22oi_4 _34106_ (.A1(_04012_),
    .A2(\timer[11] ),
    .B1(_04014_),
    .B2(\irq_mask[11] ),
    .Y(_04015_));
 sky130_fd_sc_hd__nand3_4 _34107_ (.A(_04010_),
    .B(_03954_),
    .C(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__buf_1 _34108_ (.A(_03680_),
    .X(_04017_));
 sky130_fd_sc_hd__buf_1 _34109_ (.A(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__nand4_4 _34110_ (.A(_03981_),
    .B(_03982_),
    .C(_03726_),
    .D(\count_cycle[11] ),
    .Y(_04019_));
 sky130_fd_sc_hd__buf_1 _34111_ (.A(_03787_),
    .X(_04020_));
 sky130_fd_sc_hd__nand2_4 _34112_ (.A(_04020_),
    .B(\count_instr[43] ),
    .Y(_04021_));
 sky130_fd_sc_hd__buf_1 _34113_ (.A(_03688_),
    .X(_04022_));
 sky130_fd_sc_hd__buf_1 _34114_ (.A(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__buf_1 _34115_ (.A(\count_cycle[43] ),
    .X(_04024_));
 sky130_fd_sc_hd__a22oi_4 _34116_ (.A1(_04023_),
    .A2(_23094_),
    .B1(_03960_),
    .B2(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__a41oi_4 _34117_ (.A1(_04018_),
    .A2(_04019_),
    .A3(_04021_),
    .A4(_04025_),
    .B1(_03962_),
    .Y(_04026_));
 sky130_fd_sc_hd__o21ai_4 _34118_ (.A1(_03989_),
    .A2(_03930_),
    .B1(mem_rdata[11]),
    .Y(_04027_));
 sky130_fd_sc_hd__nand3_4 _34119_ (.A(mem_rdata[27]),
    .B(_24219_),
    .C(_21379_),
    .Y(_04028_));
 sky130_fd_sc_hd__a21o_4 _34120_ (.A1(_04027_),
    .A2(_04028_),
    .B1(_03934_),
    .X(_04029_));
 sky130_fd_sc_hd__a21oi_4 _34121_ (.A1(_03927_),
    .A2(_04029_),
    .B1(_03820_),
    .Y(_04030_));
 sky130_fd_sc_hd__o21a_4 _34122_ (.A1(_03711_),
    .A2(\pcpi_mul.rd[11] ),
    .B1(_03822_),
    .X(_04031_));
 sky130_fd_sc_hd__o21a_4 _34123_ (.A1(_03710_),
    .A2(\pcpi_mul.rd[43] ),
    .B1(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__a2111oi_4 _34124_ (.A1(_04016_),
    .A2(_04026_),
    .B1(_03813_),
    .C1(_04030_),
    .D1(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__a22oi_4 _34125_ (.A1(_22029_),
    .A2(_03912_),
    .B1(_04008_),
    .B2(_04033_),
    .Y(_24255_));
 sky130_fd_sc_hd__buf_1 _34126_ (.A(_03739_),
    .X(_04034_));
 sky130_fd_sc_hd__a2111o_4 _34127_ (.A1(_20079_),
    .A2(_20101_),
    .B1(_20156_),
    .C1(_20110_),
    .D1(_04009_),
    .X(_04035_));
 sky130_fd_sc_hd__a22oi_4 _34128_ (.A1(_03914_),
    .A2(\timer[12] ),
    .B1(_03915_),
    .B2(\irq_mask[12] ),
    .Y(_04036_));
 sky130_fd_sc_hd__nand3_4 _34129_ (.A(_04035_),
    .B(_03954_),
    .C(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__nand4_4 _34130_ (.A(_03981_),
    .B(_03982_),
    .C(_03726_),
    .D(\count_cycle[12] ),
    .Y(_04038_));
 sky130_fd_sc_hd__nand2_4 _34131_ (.A(_03920_),
    .B(_23337_),
    .Y(_04039_));
 sky130_fd_sc_hd__a22oi_4 _34132_ (.A1(_03922_),
    .A2(_23101_),
    .B1(_03960_),
    .B2(\count_cycle[44] ),
    .Y(_04040_));
 sky130_fd_sc_hd__a41oi_4 _34133_ (.A1(_04018_),
    .A2(_04038_),
    .A3(_04039_),
    .A4(_04040_),
    .B1(_03962_),
    .Y(_04041_));
 sky130_fd_sc_hd__o21ai_4 _34134_ (.A1(_03989_),
    .A2(_03931_),
    .B1(mem_rdata[12]),
    .Y(_04042_));
 sky130_fd_sc_hd__nand3_4 _34135_ (.A(_01481_),
    .B(_03844_),
    .C(mem_rdata[28]),
    .Y(_04043_));
 sky130_fd_sc_hd__a21o_4 _34136_ (.A1(_04042_),
    .A2(_04043_),
    .B1(_03935_),
    .X(_04044_));
 sky130_fd_sc_hd__a21oi_4 _34137_ (.A1(_03928_),
    .A2(_04044_),
    .B1(_03937_),
    .Y(_04045_));
 sky130_fd_sc_hd__o21a_4 _34138_ (.A1(_03940_),
    .A2(\pcpi_mul.rd[12] ),
    .B1(_03670_),
    .X(_04046_));
 sky130_fd_sc_hd__o21a_4 _34139_ (.A1(_03939_),
    .A2(\pcpi_mul.rd[44] ),
    .B1(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__a2111oi_4 _34140_ (.A1(_04037_),
    .A2(_04041_),
    .B1(_03658_),
    .C1(_04045_),
    .D1(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__xnor2_4 _34141_ (.A(\decoded_imm[12] ),
    .B(\reg_pc[12] ),
    .Y(_04049_));
 sky130_fd_sc_hd__and2_4 _34142_ (.A(_03997_),
    .B(_04005_),
    .X(_04050_));
 sky130_fd_sc_hd__nand2_4 _34143_ (.A(_21221_),
    .B(\reg_pc[10] ),
    .Y(_04051_));
 sky130_vsdinv _34144_ (.A(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__maj3_4 _34145_ (.A(\decoded_imm[11] ),
    .B(_04052_),
    .C(\reg_pc[11] ),
    .X(_04053_));
 sky130_fd_sc_hd__a21oi_4 _34146_ (.A1(_04001_),
    .A2(_04050_),
    .B1(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__buf_1 _34147_ (.A(_18399_),
    .X(_04055_));
 sky130_fd_sc_hd__o21ai_4 _34148_ (.A1(_04049_),
    .A2(_04054_),
    .B1(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__a21o_4 _34149_ (.A1(_04049_),
    .A2(_04054_),
    .B1(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__a22oi_4 _34150_ (.A1(_22021_),
    .A2(_04034_),
    .B1(_04048_),
    .B2(_04057_),
    .Y(_24256_));
 sky130_fd_sc_hd__xor2_4 _34151_ (.A(\decoded_imm[13] ),
    .B(\reg_pc[13] ),
    .X(_04058_));
 sky130_vsdinv _34152_ (.A(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__nor2_4 _34153_ (.A(_21239_),
    .B(_21587_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_4 _34154_ (.A(_21238_),
    .B(\reg_pc[12] ),
    .Y(_04061_));
 sky130_fd_sc_hd__o21a_4 _34155_ (.A1(_04060_),
    .A2(_04054_),
    .B1(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__a21oi_4 _34156_ (.A1(_04062_),
    .A2(_04059_),
    .B1(_19038_),
    .Y(_04063_));
 sky130_fd_sc_hd__o21ai_4 _34157_ (.A1(_04059_),
    .A2(_04062_),
    .B1(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__buf_1 _34158_ (.A(_19193_),
    .X(_04065_));
 sky130_fd_sc_hd__a2111o_4 _34159_ (.A1(_20134_),
    .A2(_20154_),
    .B1(_04065_),
    .C1(_20169_),
    .D1(_04009_),
    .X(_04066_));
 sky130_fd_sc_hd__buf_1 _34160_ (.A(_03953_),
    .X(_04067_));
 sky130_fd_sc_hd__a22oi_4 _34161_ (.A1(_04012_),
    .A2(_18908_),
    .B1(_04014_),
    .B2(\irq_mask[13] ),
    .Y(_04068_));
 sky130_fd_sc_hd__nand3_4 _34162_ (.A(_04066_),
    .B(_04067_),
    .C(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__buf_1 _34163_ (.A(_03722_),
    .X(_04070_));
 sky130_fd_sc_hd__nand4_4 _34164_ (.A(_03981_),
    .B(_03982_),
    .C(_04070_),
    .D(\count_cycle[13] ),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_4 _34165_ (.A(_04020_),
    .B(\count_instr[45] ),
    .Y(_04072_));
 sky130_fd_sc_hd__buf_1 _34166_ (.A(instr_rdcycleh),
    .X(_04073_));
 sky130_fd_sc_hd__buf_1 _34167_ (.A(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__a22oi_4 _34168_ (.A1(_04023_),
    .A2(_23110_),
    .B1(_04074_),
    .B2(\count_cycle[45] ),
    .Y(_04075_));
 sky130_fd_sc_hd__buf_1 _34169_ (.A(_21133_),
    .X(_04076_));
 sky130_fd_sc_hd__a41oi_4 _34170_ (.A1(_04018_),
    .A2(_04071_),
    .A3(_04072_),
    .A4(_04075_),
    .B1(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__o21ai_4 _34171_ (.A1(_03989_),
    .A2(_03930_),
    .B1(mem_rdata[13]),
    .Y(_04078_));
 sky130_fd_sc_hd__nand3_4 _34172_ (.A(_24216_),
    .B(_21379_),
    .C(mem_rdata[29]),
    .Y(_04079_));
 sky130_fd_sc_hd__a21o_4 _34173_ (.A1(_04078_),
    .A2(_04079_),
    .B1(_03934_),
    .X(_04080_));
 sky130_fd_sc_hd__a21oi_4 _34174_ (.A1(_03927_),
    .A2(_04080_),
    .B1(_03820_),
    .Y(_04081_));
 sky130_fd_sc_hd__buf_1 _34175_ (.A(_03665_),
    .X(_04082_));
 sky130_fd_sc_hd__buf_1 _34176_ (.A(_03667_),
    .X(_04083_));
 sky130_fd_sc_hd__o21a_4 _34177_ (.A1(_04083_),
    .A2(\pcpi_mul.rd[13] ),
    .B1(_03822_),
    .X(_04084_));
 sky130_fd_sc_hd__o21a_4 _34178_ (.A1(_04082_),
    .A2(\pcpi_mul.rd[45] ),
    .B1(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__a2111oi_4 _34179_ (.A1(_04069_),
    .A2(_04077_),
    .B1(_03813_),
    .C1(_04081_),
    .D1(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__a22oi_4 _34180_ (.A1(_22022_),
    .A2(_04034_),
    .B1(_04064_),
    .B2(_04086_),
    .Y(_24257_));
 sky130_fd_sc_hd__xor2_4 _34181_ (.A(\decoded_imm[14] ),
    .B(\reg_pc[14] ),
    .X(_04087_));
 sky130_fd_sc_hd__or2_4 _34182_ (.A(_04049_),
    .B(_04059_),
    .X(_04088_));
 sky130_vsdinv _34183_ (.A(\reg_pc[13] ),
    .Y(_04089_));
 sky130_fd_sc_hd__maj3_4 _34184_ (.A(_21246_),
    .B(_04061_),
    .C(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__o21ai_4 _34185_ (.A1(_04088_),
    .A2(_04054_),
    .B1(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__or2_4 _34186_ (.A(_04087_),
    .B(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__buf_1 _34187_ (.A(_04055_),
    .X(_04093_));
 sky130_fd_sc_hd__nand2_4 _34188_ (.A(_04091_),
    .B(_04087_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand3_4 _34189_ (.A(_04092_),
    .B(_04093_),
    .C(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__a2111o_4 _34190_ (.A1(_20201_),
    .A2(_20218_),
    .B1(_04065_),
    .C1(_20225_),
    .D1(_04009_),
    .X(_04096_));
 sky130_fd_sc_hd__a22oi_4 _34191_ (.A1(_04012_),
    .A2(\timer[14] ),
    .B1(_04014_),
    .B2(\irq_mask[14] ),
    .Y(_04097_));
 sky130_fd_sc_hd__nand3_4 _34192_ (.A(_04096_),
    .B(_04067_),
    .C(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__buf_1 _34193_ (.A(_03856_),
    .X(_04099_));
 sky130_fd_sc_hd__buf_1 _34194_ (.A(_03858_),
    .X(_04100_));
 sky130_fd_sc_hd__buf_1 _34195_ (.A(\count_cycle[14] ),
    .X(_04101_));
 sky130_fd_sc_hd__nand4_4 _34196_ (.A(_04099_),
    .B(_04100_),
    .C(_04070_),
    .D(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand2_4 _34197_ (.A(_04020_),
    .B(\count_instr[46] ),
    .Y(_04103_));
 sky130_fd_sc_hd__a22oi_4 _34198_ (.A1(_04023_),
    .A2(_23116_),
    .B1(_04074_),
    .B2(\count_cycle[46] ),
    .Y(_04104_));
 sky130_fd_sc_hd__a41oi_4 _34199_ (.A1(_04018_),
    .A2(_04102_),
    .A3(_04103_),
    .A4(_04104_),
    .B1(_04076_),
    .Y(_04105_));
 sky130_fd_sc_hd__buf_1 _34200_ (.A(_03657_),
    .X(_04106_));
 sky130_fd_sc_hd__o21ai_4 _34201_ (.A1(_24228_),
    .A2(_03930_),
    .B1(mem_rdata[14]),
    .Y(_04107_));
 sky130_fd_sc_hd__nand3_4 _34202_ (.A(_24216_),
    .B(_21379_),
    .C(mem_rdata[30]),
    .Y(_04108_));
 sky130_fd_sc_hd__a21o_4 _34203_ (.A1(_04107_),
    .A2(_04108_),
    .B1(_03934_),
    .X(_04109_));
 sky130_fd_sc_hd__a21oi_4 _34204_ (.A1(_03927_),
    .A2(_04109_),
    .B1(_18362_),
    .Y(_04110_));
 sky130_fd_sc_hd__buf_1 _34205_ (.A(_03669_),
    .X(_04111_));
 sky130_fd_sc_hd__o21a_4 _34206_ (.A1(_04083_),
    .A2(\pcpi_mul.rd[14] ),
    .B1(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__o21a_4 _34207_ (.A1(_04082_),
    .A2(\pcpi_mul.rd[46] ),
    .B1(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__a2111oi_4 _34208_ (.A1(_04098_),
    .A2(_04105_),
    .B1(_04106_),
    .C1(_04110_),
    .D1(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__a22oi_4 _34209_ (.A1(_22023_),
    .A2(_04034_),
    .B1(_04095_),
    .B2(_04114_),
    .Y(_24258_));
 sky130_fd_sc_hd__xor2_4 _34210_ (.A(\decoded_imm[15] ),
    .B(\reg_pc[15] ),
    .X(_04115_));
 sky130_fd_sc_hd__nand2_4 _34211_ (.A(\decoded_imm[14] ),
    .B(\reg_pc[14] ),
    .Y(_04116_));
 sky130_fd_sc_hd__nand2_4 _34212_ (.A(_04094_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__or2_4 _34213_ (.A(_04115_),
    .B(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__nand2_4 _34214_ (.A(_04117_),
    .B(_04115_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand3_4 _34215_ (.A(_04118_),
    .B(_04093_),
    .C(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__buf_1 _34216_ (.A(_03716_),
    .X(_04121_));
 sky130_fd_sc_hd__a2111o_4 _34217_ (.A1(_20251_),
    .A2(_20266_),
    .B1(_04065_),
    .C1(_20274_),
    .D1(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__a22oi_4 _34218_ (.A1(_04012_),
    .A2(_20174_),
    .B1(_04014_),
    .B2(\irq_mask[15] ),
    .Y(_04123_));
 sky130_fd_sc_hd__nand3_4 _34219_ (.A(_04122_),
    .B(_04067_),
    .C(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__buf_1 _34220_ (.A(_04017_),
    .X(_04125_));
 sky130_fd_sc_hd__nand4_4 _34221_ (.A(_04099_),
    .B(_04100_),
    .C(_04070_),
    .D(\count_cycle[15] ),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_4 _34222_ (.A(_04020_),
    .B(\count_instr[47] ),
    .Y(_04127_));
 sky130_fd_sc_hd__buf_1 _34223_ (.A(\count_cycle[47] ),
    .X(_04128_));
 sky130_fd_sc_hd__a22oi_4 _34224_ (.A1(_04023_),
    .A2(\count_instr[15] ),
    .B1(_04074_),
    .B2(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__a41oi_4 _34225_ (.A1(_04125_),
    .A2(_04126_),
    .A3(_04127_),
    .A4(_04129_),
    .B1(_04076_),
    .Y(_04130_));
 sky130_vsdinv _34226_ (.A(latched_is_lh),
    .Y(_04131_));
 sky130_fd_sc_hd__o21ai_4 _34227_ (.A1(_24227_),
    .A2(_03929_),
    .B1(mem_rdata[15]),
    .Y(_04132_));
 sky130_fd_sc_hd__nand3_4 _34228_ (.A(_18295_),
    .B(_18619_),
    .C(mem_rdata[31]),
    .Y(_04133_));
 sky130_fd_sc_hd__nor2_4 _34229_ (.A(latched_is_lh),
    .B(latched_is_lb),
    .Y(_04134_));
 sky130_fd_sc_hd__a21oi_4 _34230_ (.A1(_04132_),
    .A2(_04133_),
    .B1(_04131_),
    .Y(_04135_));
 sky130_fd_sc_hd__nor2_4 _34231_ (.A(_04134_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__a21o_4 _34232_ (.A1(_03926_),
    .A2(_04136_),
    .B1(_18269_),
    .X(_04137_));
 sky130_fd_sc_hd__buf_1 _34233_ (.A(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__a41oi_4 _34234_ (.A1(_04131_),
    .A2(_03925_),
    .A3(_04132_),
    .A4(_04133_),
    .B1(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__o21a_4 _34235_ (.A1(_04083_),
    .A2(\pcpi_mul.rd[15] ),
    .B1(_04111_),
    .X(_04140_));
 sky130_fd_sc_hd__o21a_4 _34236_ (.A1(_04082_),
    .A2(\pcpi_mul.rd[47] ),
    .B1(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__a2111oi_4 _34237_ (.A1(_04124_),
    .A2(_04130_),
    .B1(_04106_),
    .C1(_04139_),
    .D1(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__a22oi_4 _34238_ (.A1(_22024_),
    .A2(_04034_),
    .B1(_04120_),
    .B2(_04142_),
    .Y(_24259_));
 sky130_fd_sc_hd__buf_1 _34239_ (.A(_03866_),
    .X(_04143_));
 sky130_fd_sc_hd__buf_1 _34240_ (.A(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__nand2_4 _34241_ (.A(_21258_),
    .B(_21649_),
    .Y(_04145_));
 sky130_fd_sc_hd__nor2_4 _34242_ (.A(_21263_),
    .B(_21664_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_4 _34243_ (.A(\decoded_imm[16] ),
    .B(\reg_pc[16] ),
    .Y(_04147_));
 sky130_vsdinv _34244_ (.A(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__nor2_4 _34245_ (.A(_04146_),
    .B(_04148_),
    .Y(_04149_));
 sky130_vsdinv _34246_ (.A(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__a21oi_4 _34247_ (.A1(_04119_),
    .A2(_04145_),
    .B1(_04150_),
    .Y(_04151_));
 sky130_vsdinv _34248_ (.A(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__nand3_4 _34249_ (.A(_04119_),
    .B(_04145_),
    .C(_04150_),
    .Y(_04153_));
 sky130_fd_sc_hd__nand3_4 _34250_ (.A(_04152_),
    .B(_04093_),
    .C(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__a2111o_4 _34251_ (.A1(_20297_),
    .A2(_20317_),
    .B1(_04065_),
    .C1(_20325_),
    .D1(_04121_),
    .X(_04155_));
 sky130_fd_sc_hd__buf_1 _34252_ (.A(_04011_),
    .X(_04156_));
 sky130_fd_sc_hd__buf_1 _34253_ (.A(_04013_),
    .X(_04157_));
 sky130_fd_sc_hd__a22oi_4 _34254_ (.A1(_04156_),
    .A2(_20328_),
    .B1(_04157_),
    .B2(\irq_mask[16] ),
    .Y(_04158_));
 sky130_fd_sc_hd__nand3_4 _34255_ (.A(_04155_),
    .B(_04067_),
    .C(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__nand4_4 _34256_ (.A(_04099_),
    .B(_04100_),
    .C(_04070_),
    .D(\count_cycle[16] ),
    .Y(_04160_));
 sky130_fd_sc_hd__buf_1 _34257_ (.A(_03787_),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_4 _34258_ (.A(_04161_),
    .B(_23361_),
    .Y(_04162_));
 sky130_fd_sc_hd__buf_1 _34259_ (.A(_04022_),
    .X(_04163_));
 sky130_fd_sc_hd__a22oi_4 _34260_ (.A1(_04163_),
    .A2(_23131_),
    .B1(_04074_),
    .B2(\count_cycle[48] ),
    .Y(_04164_));
 sky130_fd_sc_hd__a41oi_4 _34261_ (.A1(_04125_),
    .A2(_04160_),
    .A3(_04162_),
    .A4(_04164_),
    .B1(_04076_),
    .Y(_04165_));
 sky130_fd_sc_hd__buf_1 _34262_ (.A(_04134_),
    .X(_04166_));
 sky130_fd_sc_hd__buf_1 _34263_ (.A(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__buf_1 _34264_ (.A(_01485_),
    .X(_04168_));
 sky130_fd_sc_hd__buf_1 _34265_ (.A(_01487_),
    .X(_04169_));
 sky130_fd_sc_hd__nand3_4 _34266_ (.A(_04168_),
    .B(_04169_),
    .C(mem_rdata[16]),
    .Y(_04170_));
 sky130_fd_sc_hd__buf_1 _34267_ (.A(_04138_),
    .X(_04171_));
 sky130_fd_sc_hd__a21oi_4 _34268_ (.A1(_04167_),
    .A2(_04170_),
    .B1(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__o21a_4 _34269_ (.A1(_04083_),
    .A2(\pcpi_mul.rd[16] ),
    .B1(_04111_),
    .X(_04173_));
 sky130_fd_sc_hd__o21a_4 _34270_ (.A1(_04082_),
    .A2(\pcpi_mul.rd[48] ),
    .B1(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__a2111oi_4 _34271_ (.A1(_04159_),
    .A2(_04165_),
    .B1(_04106_),
    .C1(_04172_),
    .D1(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__a22oi_4 _34272_ (.A1(_22004_),
    .A2(_04144_),
    .B1(_04154_),
    .B2(_04175_),
    .Y(_24260_));
 sky130_fd_sc_hd__xor2_4 _34273_ (.A(\decoded_imm[17] ),
    .B(\reg_pc[17] ),
    .X(_04176_));
 sky130_fd_sc_hd__a211o_4 _34274_ (.A1(_21264_),
    .A2(_21665_),
    .B1(_04176_),
    .C1(_04151_),
    .X(_04177_));
 sky130_fd_sc_hd__o21ai_4 _34275_ (.A1(_04148_),
    .A2(_04151_),
    .B1(_04176_),
    .Y(_04178_));
 sky130_fd_sc_hd__nand3_4 _34276_ (.A(_04177_),
    .B(_04178_),
    .C(_03885_),
    .Y(_04179_));
 sky130_fd_sc_hd__buf_1 _34277_ (.A(_20029_),
    .X(_04180_));
 sky130_fd_sc_hd__a2111o_4 _34278_ (.A1(_20351_),
    .A2(_20365_),
    .B1(_04180_),
    .C1(_20373_),
    .D1(_04121_),
    .X(_04181_));
 sky130_fd_sc_hd__buf_1 _34279_ (.A(_03953_),
    .X(_04182_));
 sky130_fd_sc_hd__a22oi_4 _34280_ (.A1(_04156_),
    .A2(\timer[17] ),
    .B1(_04157_),
    .B2(\irq_mask[17] ),
    .Y(_04183_));
 sky130_fd_sc_hd__nand3_4 _34281_ (.A(_04181_),
    .B(_04182_),
    .C(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__buf_1 _34282_ (.A(_24093_),
    .X(_04185_));
 sky130_fd_sc_hd__nand4_4 _34283_ (.A(_04099_),
    .B(_04100_),
    .C(_04185_),
    .D(\count_cycle[17] ),
    .Y(_04186_));
 sky130_fd_sc_hd__nand2_4 _34284_ (.A(_04161_),
    .B(\count_instr[49] ),
    .Y(_04187_));
 sky130_fd_sc_hd__buf_1 _34285_ (.A(_04073_),
    .X(_04188_));
 sky130_fd_sc_hd__a22oi_4 _34286_ (.A1(_04163_),
    .A2(_23146_),
    .B1(_04188_),
    .B2(\count_cycle[49] ),
    .Y(_04189_));
 sky130_fd_sc_hd__buf_1 _34287_ (.A(_21133_),
    .X(_04190_));
 sky130_fd_sc_hd__a41oi_4 _34288_ (.A1(_04125_),
    .A2(_04186_),
    .A3(_04187_),
    .A4(_04189_),
    .B1(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand3_4 _34289_ (.A(_04168_),
    .B(_04169_),
    .C(mem_rdata[17]),
    .Y(_04192_));
 sky130_fd_sc_hd__a21oi_4 _34290_ (.A1(_04167_),
    .A2(_04192_),
    .B1(_04171_),
    .Y(_04193_));
 sky130_fd_sc_hd__buf_1 _34291_ (.A(_03740_),
    .X(_04194_));
 sky130_fd_sc_hd__buf_1 _34292_ (.A(_03742_),
    .X(_04195_));
 sky130_fd_sc_hd__o21a_4 _34293_ (.A1(_04195_),
    .A2(\pcpi_mul.rd[17] ),
    .B1(_04111_),
    .X(_04196_));
 sky130_fd_sc_hd__o21a_4 _34294_ (.A1(_04194_),
    .A2(\pcpi_mul.rd[49] ),
    .B1(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__a2111oi_4 _34295_ (.A1(_04184_),
    .A2(_04191_),
    .B1(_04106_),
    .C1(_04193_),
    .D1(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__a22oi_4 _34296_ (.A1(_22005_),
    .A2(_04144_),
    .B1(_04179_),
    .B2(_04198_),
    .Y(_24261_));
 sky130_fd_sc_hd__xor2_4 _34297_ (.A(\decoded_imm[18] ),
    .B(\reg_pc[18] ),
    .X(_04199_));
 sky130_fd_sc_hd__maj3_4 _34298_ (.A(\decoded_imm[17] ),
    .B(_04148_),
    .C(\reg_pc[17] ),
    .X(_04200_));
 sky130_fd_sc_hd__and2_4 _34299_ (.A(_04176_),
    .B(_04149_),
    .X(_04201_));
 sky130_fd_sc_hd__a21boi_4 _34300_ (.A1(_04119_),
    .A2(_04145_),
    .B1_N(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__or3_4 _34301_ (.A(_04199_),
    .B(_04200_),
    .C(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__o21ai_4 _34302_ (.A1(_04200_),
    .A2(_04202_),
    .B1(_04199_),
    .Y(_04204_));
 sky130_fd_sc_hd__nand3_4 _34303_ (.A(_04203_),
    .B(_04093_),
    .C(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__a2111o_4 _34304_ (.A1(_20406_),
    .A2(_20420_),
    .B1(_04180_),
    .C1(_20427_),
    .D1(_04121_),
    .X(_04206_));
 sky130_fd_sc_hd__a22oi_4 _34305_ (.A1(_04156_),
    .A2(_20387_),
    .B1(_04157_),
    .B2(\irq_mask[18] ),
    .Y(_04207_));
 sky130_fd_sc_hd__nand3_4 _34306_ (.A(_04206_),
    .B(_04182_),
    .C(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__buf_1 _34307_ (.A(_03856_),
    .X(_04209_));
 sky130_fd_sc_hd__buf_1 _34308_ (.A(_03858_),
    .X(_04210_));
 sky130_fd_sc_hd__nand4_4 _34309_ (.A(_04209_),
    .B(_04210_),
    .C(_04185_),
    .D(\count_cycle[18] ),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2_4 _34310_ (.A(_04161_),
    .B(_23374_),
    .Y(_04212_));
 sky130_fd_sc_hd__a22oi_4 _34311_ (.A1(_04163_),
    .A2(\count_instr[18] ),
    .B1(_04188_),
    .B2(\count_cycle[50] ),
    .Y(_04213_));
 sky130_fd_sc_hd__a41oi_4 _34312_ (.A1(_04125_),
    .A2(_04211_),
    .A3(_04212_),
    .A4(_04213_),
    .B1(_04190_),
    .Y(_04214_));
 sky130_fd_sc_hd__buf_1 _34313_ (.A(_03641_),
    .X(_04215_));
 sky130_fd_sc_hd__nand3_4 _34314_ (.A(_04168_),
    .B(_04169_),
    .C(mem_rdata[18]),
    .Y(_04216_));
 sky130_fd_sc_hd__a21oi_4 _34315_ (.A1(_04167_),
    .A2(_04216_),
    .B1(_04171_),
    .Y(_04217_));
 sky130_fd_sc_hd__buf_1 _34316_ (.A(_03669_),
    .X(_04218_));
 sky130_fd_sc_hd__o21a_4 _34317_ (.A1(_04195_),
    .A2(\pcpi_mul.rd[18] ),
    .B1(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__o21a_4 _34318_ (.A1(_04194_),
    .A2(\pcpi_mul.rd[50] ),
    .B1(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__a2111oi_4 _34319_ (.A1(_04208_),
    .A2(_04214_),
    .B1(_04215_),
    .C1(_04217_),
    .D1(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a22oi_4 _34320_ (.A1(_22006_),
    .A2(_04144_),
    .B1(_04205_),
    .B2(_04221_),
    .Y(_24262_));
 sky130_fd_sc_hd__nand2_4 _34321_ (.A(\decoded_imm[18] ),
    .B(\reg_pc[18] ),
    .Y(_04222_));
 sky130_fd_sc_hd__xor2_4 _34322_ (.A(\decoded_imm[19] ),
    .B(\reg_pc[19] ),
    .X(_04223_));
 sky130_vsdinv _34323_ (.A(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__a21oi_4 _34324_ (.A1(_04204_),
    .A2(_04222_),
    .B1(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__and3_4 _34325_ (.A(_04204_),
    .B(_04222_),
    .C(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__or3_4 _34326_ (.A(_04002_),
    .B(_04225_),
    .C(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__buf_1 _34327_ (.A(_03715_),
    .X(_04228_));
 sky130_fd_sc_hd__a2111o_4 _34328_ (.A1(_20456_),
    .A2(_20470_),
    .B1(_04180_),
    .C1(_20477_),
    .D1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__a22oi_4 _34329_ (.A1(_04156_),
    .A2(\timer[19] ),
    .B1(_04157_),
    .B2(\irq_mask[19] ),
    .Y(_04230_));
 sky130_fd_sc_hd__nand3_4 _34330_ (.A(_04229_),
    .B(_04182_),
    .C(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__buf_1 _34331_ (.A(_04017_),
    .X(_04232_));
 sky130_fd_sc_hd__nand4_4 _34332_ (.A(_04209_),
    .B(_04210_),
    .C(_04185_),
    .D(\count_cycle[19] ),
    .Y(_04233_));
 sky130_fd_sc_hd__nand2_4 _34333_ (.A(_04161_),
    .B(\count_instr[51] ),
    .Y(_04234_));
 sky130_fd_sc_hd__buf_1 _34334_ (.A(\count_cycle[51] ),
    .X(_04235_));
 sky130_fd_sc_hd__a22oi_4 _34335_ (.A1(_04163_),
    .A2(\count_instr[19] ),
    .B1(_04188_),
    .B2(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__a41oi_4 _34336_ (.A1(_04232_),
    .A2(_04233_),
    .A3(_04234_),
    .A4(_04236_),
    .B1(_04190_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand3_4 _34337_ (.A(_04168_),
    .B(_04169_),
    .C(mem_rdata[19]),
    .Y(_04238_));
 sky130_fd_sc_hd__a21oi_4 _34338_ (.A1(_04167_),
    .A2(_04238_),
    .B1(_04171_),
    .Y(_04239_));
 sky130_fd_sc_hd__o21a_4 _34339_ (.A1(_04195_),
    .A2(\pcpi_mul.rd[19] ),
    .B1(_04218_),
    .X(_04240_));
 sky130_fd_sc_hd__o21a_4 _34340_ (.A1(_04194_),
    .A2(\pcpi_mul.rd[51] ),
    .B1(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__a2111oi_4 _34341_ (.A1(_04231_),
    .A2(_04237_),
    .B1(_04215_),
    .C1(_04239_),
    .D1(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__a22oi_4 _34342_ (.A1(_22007_),
    .A2(_04144_),
    .B1(_04227_),
    .B2(_04242_),
    .Y(_24263_));
 sky130_fd_sc_hd__buf_1 _34343_ (.A(_04143_),
    .X(_04243_));
 sky130_fd_sc_hd__xor2_4 _34344_ (.A(\decoded_imm[20] ),
    .B(\reg_pc[20] ),
    .X(_04244_));
 sky130_fd_sc_hd__a211o_4 _34345_ (.A1(_21281_),
    .A2(_21717_),
    .B1(_04244_),
    .C1(_04225_),
    .X(_04245_));
 sky130_fd_sc_hd__buf_1 _34346_ (.A(_04055_),
    .X(_04246_));
 sky130_fd_sc_hd__nand2_4 _34347_ (.A(\decoded_imm[19] ),
    .B(_21716_),
    .Y(_04247_));
 sky130_vsdinv _34348_ (.A(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__o21ai_4 _34349_ (.A1(_04248_),
    .A2(_04225_),
    .B1(_04244_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand3_4 _34350_ (.A(_04245_),
    .B(_04246_),
    .C(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__a2111o_4 _34351_ (.A1(_20500_),
    .A2(_20514_),
    .B1(_04180_),
    .C1(_20524_),
    .D1(_04228_),
    .X(_04251_));
 sky130_fd_sc_hd__buf_1 _34352_ (.A(_04011_),
    .X(_04252_));
 sky130_fd_sc_hd__buf_1 _34353_ (.A(_04013_),
    .X(_04253_));
 sky130_fd_sc_hd__a22oi_4 _34354_ (.A1(_04252_),
    .A2(\timer[20] ),
    .B1(_04253_),
    .B2(\irq_mask[20] ),
    .Y(_04254_));
 sky130_fd_sc_hd__nand3_4 _34355_ (.A(_04251_),
    .B(_04182_),
    .C(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand4_4 _34356_ (.A(_04209_),
    .B(_04210_),
    .C(_04185_),
    .D(\count_cycle[20] ),
    .Y(_04256_));
 sky130_fd_sc_hd__buf_1 _34357_ (.A(_03787_),
    .X(_04257_));
 sky130_fd_sc_hd__nand2_4 _34358_ (.A(_04257_),
    .B(_23384_),
    .Y(_04258_));
 sky130_fd_sc_hd__buf_1 _34359_ (.A(_04022_),
    .X(_04259_));
 sky130_fd_sc_hd__buf_1 _34360_ (.A(\count_cycle[52] ),
    .X(_04260_));
 sky130_fd_sc_hd__a22oi_4 _34361_ (.A1(_04259_),
    .A2(_23170_),
    .B1(_04188_),
    .B2(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__a41oi_4 _34362_ (.A1(_04232_),
    .A2(_04256_),
    .A3(_04258_),
    .A4(_04261_),
    .B1(_04190_),
    .Y(_04262_));
 sky130_fd_sc_hd__buf_1 _34363_ (.A(_04166_),
    .X(_04263_));
 sky130_fd_sc_hd__buf_1 _34364_ (.A(_01485_),
    .X(_04264_));
 sky130_fd_sc_hd__buf_1 _34365_ (.A(_01487_),
    .X(_04265_));
 sky130_fd_sc_hd__nand3_4 _34366_ (.A(_04264_),
    .B(_04265_),
    .C(mem_rdata[20]),
    .Y(_04266_));
 sky130_fd_sc_hd__buf_1 _34367_ (.A(_04138_),
    .X(_04267_));
 sky130_fd_sc_hd__a21oi_4 _34368_ (.A1(_04263_),
    .A2(_04266_),
    .B1(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__o21a_4 _34369_ (.A1(_04195_),
    .A2(\pcpi_mul.rd[20] ),
    .B1(_04218_),
    .X(_04269_));
 sky130_fd_sc_hd__o21a_4 _34370_ (.A1(_04194_),
    .A2(\pcpi_mul.rd[52] ),
    .B1(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__a2111oi_4 _34371_ (.A1(_04255_),
    .A2(_04262_),
    .B1(_04215_),
    .C1(_04268_),
    .D1(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__a22oi_4 _34372_ (.A1(_21999_),
    .A2(_04243_),
    .B1(_04250_),
    .B2(_04271_),
    .Y(_24265_));
 sky130_fd_sc_hd__nand2_4 _34373_ (.A(\decoded_imm[20] ),
    .B(\reg_pc[20] ),
    .Y(_04272_));
 sky130_fd_sc_hd__xor2_4 _34374_ (.A(\decoded_imm[21] ),
    .B(\reg_pc[21] ),
    .X(_04273_));
 sky130_vsdinv _34375_ (.A(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__a21oi_4 _34376_ (.A1(_04249_),
    .A2(_04272_),
    .B1(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__and3_4 _34377_ (.A(_04249_),
    .B(_04272_),
    .C(_04274_),
    .X(_04276_));
 sky130_fd_sc_hd__or3_4 _34378_ (.A(_04002_),
    .B(_04275_),
    .C(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__buf_1 _34379_ (.A(_20029_),
    .X(_04278_));
 sky130_fd_sc_hd__a2111o_4 _34380_ (.A1(_20551_),
    .A2(_20565_),
    .B1(_04278_),
    .C1(_20572_),
    .D1(_04228_),
    .X(_04279_));
 sky130_fd_sc_hd__buf_1 _34381_ (.A(_03953_),
    .X(_04280_));
 sky130_fd_sc_hd__a22oi_4 _34382_ (.A1(_04252_),
    .A2(\timer[21] ),
    .B1(_04253_),
    .B2(\irq_mask[21] ),
    .Y(_04281_));
 sky130_fd_sc_hd__nand3_4 _34383_ (.A(_04279_),
    .B(_04280_),
    .C(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__buf_1 _34384_ (.A(_24093_),
    .X(_04283_));
 sky130_fd_sc_hd__nand4_4 _34385_ (.A(_04209_),
    .B(_04210_),
    .C(_04283_),
    .D(\count_cycle[21] ),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_4 _34386_ (.A(_04257_),
    .B(\count_instr[53] ),
    .Y(_04285_));
 sky130_fd_sc_hd__buf_1 _34387_ (.A(_04073_),
    .X(_04286_));
 sky130_fd_sc_hd__buf_1 _34388_ (.A(\count_cycle[53] ),
    .X(_04287_));
 sky130_fd_sc_hd__a22oi_4 _34389_ (.A1(_04259_),
    .A2(\count_instr[21] ),
    .B1(_04286_),
    .B2(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__buf_1 _34390_ (.A(_21214_),
    .X(_04289_));
 sky130_fd_sc_hd__a41oi_4 _34391_ (.A1(_04232_),
    .A2(_04284_),
    .A3(_04285_),
    .A4(_04288_),
    .B1(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand3_4 _34392_ (.A(_04264_),
    .B(_04265_),
    .C(mem_rdata[21]),
    .Y(_04291_));
 sky130_fd_sc_hd__a21oi_4 _34393_ (.A1(_04263_),
    .A2(_04291_),
    .B1(_04267_),
    .Y(_04292_));
 sky130_fd_sc_hd__buf_1 _34394_ (.A(_03740_),
    .X(_04293_));
 sky130_fd_sc_hd__buf_1 _34395_ (.A(_03742_),
    .X(_04294_));
 sky130_fd_sc_hd__o21a_4 _34396_ (.A1(_04294_),
    .A2(\pcpi_mul.rd[21] ),
    .B1(_04218_),
    .X(_04295_));
 sky130_fd_sc_hd__o21a_4 _34397_ (.A1(_04293_),
    .A2(\pcpi_mul.rd[53] ),
    .B1(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__a2111oi_4 _34398_ (.A1(_04282_),
    .A2(_04290_),
    .B1(_04215_),
    .C1(_04292_),
    .D1(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__a22oi_4 _34399_ (.A1(_22000_),
    .A2(_04243_),
    .B1(_04277_),
    .B2(_04297_),
    .Y(_24266_));
 sky130_fd_sc_hd__a21o_4 _34400_ (.A1(\decoded_imm[21] ),
    .A2(\reg_pc[21] ),
    .B1(_04275_),
    .X(_04298_));
 sky130_fd_sc_hd__xor2_4 _34401_ (.A(\decoded_imm[22] ),
    .B(\reg_pc[22] ),
    .X(_04299_));
 sky130_fd_sc_hd__nand2_4 _34402_ (.A(_04298_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__a211o_4 _34403_ (.A1(_21292_),
    .A2(_21743_),
    .B1(_04299_),
    .C1(_04275_),
    .X(_04301_));
 sky130_fd_sc_hd__nand3_4 _34404_ (.A(_04300_),
    .B(_04301_),
    .C(_03885_),
    .Y(_04302_));
 sky130_fd_sc_hd__a21o_4 _34405_ (.A1(_24050_),
    .A2(_18511_),
    .B1(_20617_),
    .X(_04303_));
 sky130_fd_sc_hd__a22oi_4 _34406_ (.A1(_04252_),
    .A2(_20575_),
    .B1(_04253_),
    .B2(\irq_mask[22] ),
    .Y(_04304_));
 sky130_fd_sc_hd__nand3_4 _34407_ (.A(_04303_),
    .B(_04280_),
    .C(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__buf_1 _34408_ (.A(_24085_),
    .X(_04306_));
 sky130_fd_sc_hd__buf_1 _34409_ (.A(_24072_),
    .X(_04307_));
 sky130_fd_sc_hd__buf_1 _34410_ (.A(\count_cycle[22] ),
    .X(_04308_));
 sky130_fd_sc_hd__nand4_4 _34411_ (.A(_04306_),
    .B(_04307_),
    .C(_04283_),
    .D(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__nand2_4 _34412_ (.A(_04257_),
    .B(\count_instr[54] ),
    .Y(_04310_));
 sky130_fd_sc_hd__buf_1 _34413_ (.A(\count_cycle[54] ),
    .X(_04311_));
 sky130_fd_sc_hd__a22oi_4 _34414_ (.A1(_04259_),
    .A2(_23185_),
    .B1(_04286_),
    .B2(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__a41oi_4 _34415_ (.A1(_04232_),
    .A2(_04309_),
    .A3(_04310_),
    .A4(_04312_),
    .B1(_04289_),
    .Y(_04313_));
 sky130_fd_sc_hd__buf_1 _34416_ (.A(_03641_),
    .X(_04314_));
 sky130_fd_sc_hd__nand3_4 _34417_ (.A(_04264_),
    .B(_04265_),
    .C(mem_rdata[22]),
    .Y(_04315_));
 sky130_fd_sc_hd__a21oi_4 _34418_ (.A1(_04263_),
    .A2(_04315_),
    .B1(_04267_),
    .Y(_04316_));
 sky130_fd_sc_hd__buf_1 _34419_ (.A(_18501_),
    .X(_04317_));
 sky130_fd_sc_hd__o21a_4 _34420_ (.A1(_04294_),
    .A2(\pcpi_mul.rd[22] ),
    .B1(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__o21a_4 _34421_ (.A1(_04293_),
    .A2(\pcpi_mul.rd[54] ),
    .B1(_04318_),
    .X(_04319_));
 sky130_fd_sc_hd__a2111oi_4 _34422_ (.A1(_04305_),
    .A2(_04313_),
    .B1(_04314_),
    .C1(_04316_),
    .D1(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__a22oi_4 _34423_ (.A1(_22001_),
    .A2(_04243_),
    .B1(_04302_),
    .B2(_04320_),
    .Y(_24267_));
 sky130_fd_sc_hd__nand2_4 _34424_ (.A(\decoded_imm[23] ),
    .B(_21772_),
    .Y(_04321_));
 sky130_fd_sc_hd__buf_1 _34425_ (.A(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__nand2_4 _34426_ (.A(_21301_),
    .B(_02119_),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2_4 _34427_ (.A(_21296_),
    .B(\reg_pc[22] ),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_4 _34428_ (.A(_04300_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__a21o_4 _34429_ (.A1(_04322_),
    .A2(_04323_),
    .B1(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__nand3_4 _34430_ (.A(_04325_),
    .B(_04322_),
    .C(_04323_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand3_4 _34431_ (.A(_04326_),
    .B(_04246_),
    .C(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__a2111o_4 _34432_ (.A1(_20634_),
    .A2(_20648_),
    .B1(_04278_),
    .C1(_20656_),
    .D1(_04228_),
    .X(_04329_));
 sky130_fd_sc_hd__a22oi_4 _34433_ (.A1(_04252_),
    .A2(\timer[23] ),
    .B1(_04253_),
    .B2(\irq_mask[23] ),
    .Y(_04330_));
 sky130_fd_sc_hd__nand3_4 _34434_ (.A(_04329_),
    .B(_04280_),
    .C(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__buf_1 _34435_ (.A(_04017_),
    .X(_04332_));
 sky130_fd_sc_hd__buf_1 _34436_ (.A(\count_cycle[23] ),
    .X(_04333_));
 sky130_fd_sc_hd__nand4_4 _34437_ (.A(_04306_),
    .B(_04307_),
    .C(_04283_),
    .D(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__nand2_4 _34438_ (.A(_04257_),
    .B(\count_instr[55] ),
    .Y(_04335_));
 sky130_fd_sc_hd__buf_1 _34439_ (.A(\count_cycle[55] ),
    .X(_04336_));
 sky130_fd_sc_hd__a22oi_4 _34440_ (.A1(_04259_),
    .A2(\count_instr[23] ),
    .B1(_04286_),
    .B2(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__a41oi_4 _34441_ (.A1(_04332_),
    .A2(_04334_),
    .A3(_04335_),
    .A4(_04337_),
    .B1(_04289_),
    .Y(_04338_));
 sky130_fd_sc_hd__nand3_4 _34442_ (.A(_04264_),
    .B(_04265_),
    .C(mem_rdata[23]),
    .Y(_04339_));
 sky130_fd_sc_hd__a21oi_4 _34443_ (.A1(_04263_),
    .A2(_04339_),
    .B1(_04267_),
    .Y(_04340_));
 sky130_fd_sc_hd__o21a_4 _34444_ (.A1(_04294_),
    .A2(\pcpi_mul.rd[23] ),
    .B1(_04317_),
    .X(_04341_));
 sky130_fd_sc_hd__o21a_4 _34445_ (.A1(_04293_),
    .A2(\pcpi_mul.rd[55] ),
    .B1(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__a2111oi_4 _34446_ (.A1(_04331_),
    .A2(_04338_),
    .B1(_04314_),
    .C1(_04340_),
    .D1(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__a22oi_4 _34447_ (.A1(_22002_),
    .A2(_04243_),
    .B1(_04328_),
    .B2(_04343_),
    .Y(_24268_));
 sky130_fd_sc_hd__buf_1 _34448_ (.A(_04143_),
    .X(_04344_));
 sky130_fd_sc_hd__xor2_4 _34449_ (.A(\decoded_imm[24] ),
    .B(\reg_pc[24] ),
    .X(_04345_));
 sky130_vsdinv _34450_ (.A(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__a21o_4 _34451_ (.A1(_04327_),
    .A2(_04322_),
    .B1(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__nand3_4 _34452_ (.A(_04327_),
    .B(_04322_),
    .C(_04346_),
    .Y(_04348_));
 sky130_fd_sc_hd__nand3_4 _34453_ (.A(_04347_),
    .B(_04246_),
    .C(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__buf_1 _34454_ (.A(_03715_),
    .X(_04350_));
 sky130_fd_sc_hd__a2111o_4 _34455_ (.A1(_20680_),
    .A2(_20695_),
    .B1(_04278_),
    .C1(_20703_),
    .D1(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__buf_1 _34456_ (.A(_04011_),
    .X(_04352_));
 sky130_fd_sc_hd__buf_1 _34457_ (.A(_04013_),
    .X(_04353_));
 sky130_fd_sc_hd__a22oi_4 _34458_ (.A1(_04352_),
    .A2(\timer[24] ),
    .B1(_04353_),
    .B2(\irq_mask[24] ),
    .Y(_04354_));
 sky130_fd_sc_hd__nand3_4 _34459_ (.A(_04351_),
    .B(_04280_),
    .C(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__buf_1 _34460_ (.A(\count_cycle[24] ),
    .X(_04356_));
 sky130_fd_sc_hd__nand4_4 _34461_ (.A(_04306_),
    .B(_04307_),
    .C(_04283_),
    .D(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__buf_1 _34462_ (.A(_03684_),
    .X(_04358_));
 sky130_fd_sc_hd__nand2_4 _34463_ (.A(_04358_),
    .B(\count_instr[56] ),
    .Y(_04359_));
 sky130_fd_sc_hd__buf_1 _34464_ (.A(_04022_),
    .X(_04360_));
 sky130_fd_sc_hd__buf_1 _34465_ (.A(\count_cycle[56] ),
    .X(_04361_));
 sky130_fd_sc_hd__a22oi_4 _34466_ (.A1(_04360_),
    .A2(_23198_),
    .B1(_04286_),
    .B2(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__a41oi_4 _34467_ (.A1(_04332_),
    .A2(_04357_),
    .A3(_04359_),
    .A4(_04362_),
    .B1(_04289_),
    .Y(_04363_));
 sky130_fd_sc_hd__buf_1 _34468_ (.A(_04166_),
    .X(_04364_));
 sky130_fd_sc_hd__buf_1 _34469_ (.A(_01484_),
    .X(_04365_));
 sky130_fd_sc_hd__buf_1 _34470_ (.A(_24240_),
    .X(_04366_));
 sky130_fd_sc_hd__nand3_4 _34471_ (.A(_04365_),
    .B(_04366_),
    .C(mem_rdata[24]),
    .Y(_04367_));
 sky130_fd_sc_hd__buf_1 _34472_ (.A(_04138_),
    .X(_04368_));
 sky130_fd_sc_hd__a21oi_4 _34473_ (.A1(_04364_),
    .A2(_04367_),
    .B1(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__o21a_4 _34474_ (.A1(_04294_),
    .A2(\pcpi_mul.rd[24] ),
    .B1(_04317_),
    .X(_04370_));
 sky130_fd_sc_hd__o21a_4 _34475_ (.A1(_04293_),
    .A2(\pcpi_mul.rd[56] ),
    .B1(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__a2111oi_4 _34476_ (.A1(_04355_),
    .A2(_04363_),
    .B1(_04314_),
    .C1(_04369_),
    .D1(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__a22oi_4 _34477_ (.A1(_22015_),
    .A2(_04344_),
    .B1(_04349_),
    .B2(_04372_),
    .Y(_24269_));
 sky130_fd_sc_hd__nand2_4 _34478_ (.A(_21305_),
    .B(\reg_pc[24] ),
    .Y(_04373_));
 sky130_fd_sc_hd__xor2_4 _34479_ (.A(_21311_),
    .B(\reg_pc[25] ),
    .X(_04374_));
 sky130_vsdinv _34480_ (.A(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__a21o_4 _34481_ (.A1(_04347_),
    .A2(_04373_),
    .B1(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__nand3_4 _34482_ (.A(_04347_),
    .B(_04373_),
    .C(_04375_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand3_4 _34483_ (.A(_04376_),
    .B(_04246_),
    .C(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__a2111o_4 _34484_ (.A1(_20727_),
    .A2(_20742_),
    .B1(_04278_),
    .C1(_20749_),
    .D1(_04350_),
    .X(_04379_));
 sky130_fd_sc_hd__buf_1 _34485_ (.A(_18515_),
    .X(_04380_));
 sky130_fd_sc_hd__a22oi_4 _34486_ (.A1(_04352_),
    .A2(\timer[25] ),
    .B1(_04353_),
    .B2(\irq_mask[25] ),
    .Y(_04381_));
 sky130_fd_sc_hd__nand3_4 _34487_ (.A(_04379_),
    .B(_04380_),
    .C(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__buf_1 _34488_ (.A(_24093_),
    .X(_04383_));
 sky130_fd_sc_hd__nand4_4 _34489_ (.A(_04306_),
    .B(_04307_),
    .C(_04383_),
    .D(\count_cycle[25] ),
    .Y(_04384_));
 sky130_fd_sc_hd__nand2_4 _34490_ (.A(_04358_),
    .B(_23415_),
    .Y(_04385_));
 sky130_fd_sc_hd__buf_1 _34491_ (.A(_04073_),
    .X(_04386_));
 sky130_fd_sc_hd__buf_1 _34492_ (.A(\count_cycle[57] ),
    .X(_04387_));
 sky130_fd_sc_hd__a22oi_4 _34493_ (.A1(_04360_),
    .A2(_23205_),
    .B1(_04386_),
    .B2(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__buf_1 _34494_ (.A(_21214_),
    .X(_04389_));
 sky130_fd_sc_hd__a41oi_4 _34495_ (.A1(_04332_),
    .A2(_04384_),
    .A3(_04385_),
    .A4(_04388_),
    .B1(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand3_4 _34496_ (.A(_04365_),
    .B(_04366_),
    .C(mem_rdata[25]),
    .Y(_04391_));
 sky130_fd_sc_hd__a21oi_4 _34497_ (.A1(_04364_),
    .A2(_04391_),
    .B1(_04368_),
    .Y(_04392_));
 sky130_fd_sc_hd__buf_1 _34498_ (.A(_03740_),
    .X(_04393_));
 sky130_fd_sc_hd__buf_1 _34499_ (.A(_03742_),
    .X(_04394_));
 sky130_fd_sc_hd__o21a_4 _34500_ (.A1(_04394_),
    .A2(\pcpi_mul.rd[25] ),
    .B1(_04317_),
    .X(_04395_));
 sky130_fd_sc_hd__o21a_4 _34501_ (.A1(_04393_),
    .A2(\pcpi_mul.rd[57] ),
    .B1(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__a2111oi_4 _34502_ (.A1(_04382_),
    .A2(_04390_),
    .B1(_04314_),
    .C1(_04392_),
    .D1(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__a22oi_4 _34503_ (.A1(_22016_),
    .A2(_04344_),
    .B1(_04378_),
    .B2(_04397_),
    .Y(_24270_));
 sky130_fd_sc_hd__xor2_4 _34504_ (.A(_21318_),
    .B(\reg_pc[26] ),
    .X(_04398_));
 sky130_fd_sc_hd__and2_4 _34505_ (.A(_04345_),
    .B(_04374_),
    .X(_04399_));
 sky130_vsdinv _34506_ (.A(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__a21boi_4 _34507_ (.A1(_04325_),
    .A2(_04323_),
    .B1_N(_04321_),
    .Y(_04401_));
 sky130_fd_sc_hd__maj3_4 _34508_ (.A(_21312_),
    .B(_04373_),
    .C(_02150_),
    .X(_04402_));
 sky130_fd_sc_hd__o21ai_4 _34509_ (.A1(_04400_),
    .A2(_04401_),
    .B1(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__or2_4 _34510_ (.A(_04398_),
    .B(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__buf_1 _34511_ (.A(_18400_),
    .X(_04405_));
 sky130_fd_sc_hd__nand2_4 _34512_ (.A(_04403_),
    .B(_04398_),
    .Y(_04406_));
 sky130_fd_sc_hd__nand3_4 _34513_ (.A(_04404_),
    .B(_04405_),
    .C(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__buf_1 _34514_ (.A(_20029_),
    .X(_04408_));
 sky130_fd_sc_hd__a2111o_4 _34515_ (.A1(_20770_),
    .A2(_20784_),
    .B1(_04408_),
    .C1(_20792_),
    .D1(_04350_),
    .X(_04409_));
 sky130_fd_sc_hd__a22oi_4 _34516_ (.A1(_04352_),
    .A2(\timer[26] ),
    .B1(_04353_),
    .B2(\irq_mask[26] ),
    .Y(_04410_));
 sky130_fd_sc_hd__nand3_4 _34517_ (.A(_04409_),
    .B(_04380_),
    .C(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__buf_1 _34518_ (.A(_24085_),
    .X(_04412_));
 sky130_fd_sc_hd__buf_1 _34519_ (.A(_24072_),
    .X(_04413_));
 sky130_fd_sc_hd__buf_1 _34520_ (.A(\count_cycle[26] ),
    .X(_04414_));
 sky130_fd_sc_hd__nand4_4 _34521_ (.A(_04412_),
    .B(_04413_),
    .C(_04383_),
    .D(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__nand2_4 _34522_ (.A(_04358_),
    .B(_23419_),
    .Y(_04416_));
 sky130_fd_sc_hd__buf_1 _34523_ (.A(\count_cycle[58] ),
    .X(_04417_));
 sky130_fd_sc_hd__a22oi_4 _34524_ (.A1(_04360_),
    .A2(_23213_),
    .B1(_04386_),
    .B2(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__a41oi_4 _34525_ (.A1(_04332_),
    .A2(_04415_),
    .A3(_04416_),
    .A4(_04418_),
    .B1(_04389_),
    .Y(_04419_));
 sky130_fd_sc_hd__buf_1 _34526_ (.A(_03641_),
    .X(_04420_));
 sky130_fd_sc_hd__nand3_4 _34527_ (.A(_04365_),
    .B(_04366_),
    .C(mem_rdata[26]),
    .Y(_04421_));
 sky130_fd_sc_hd__a21oi_4 _34528_ (.A1(_04364_),
    .A2(_04421_),
    .B1(_04368_),
    .Y(_04422_));
 sky130_fd_sc_hd__buf_1 _34529_ (.A(_18501_),
    .X(_04423_));
 sky130_fd_sc_hd__o21a_4 _34530_ (.A1(_04394_),
    .A2(\pcpi_mul.rd[26] ),
    .B1(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__o21a_4 _34531_ (.A1(_04393_),
    .A2(\pcpi_mul.rd[58] ),
    .B1(_04424_),
    .X(_04425_));
 sky130_fd_sc_hd__a2111oi_4 _34532_ (.A1(_04411_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04422_),
    .D1(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__a22oi_4 _34533_ (.A1(_22017_),
    .A2(_04344_),
    .B1(_04407_),
    .B2(_04426_),
    .Y(_24271_));
 sky130_fd_sc_hd__nand2_4 _34534_ (.A(\decoded_imm[26] ),
    .B(\reg_pc[26] ),
    .Y(_04427_));
 sky130_fd_sc_hd__xor2_4 _34535_ (.A(_21321_),
    .B(\reg_pc[27] ),
    .X(_04428_));
 sky130_vsdinv _34536_ (.A(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__a21o_4 _34537_ (.A1(_04406_),
    .A2(_04427_),
    .B1(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__nand3_4 _34538_ (.A(_04406_),
    .B(_04427_),
    .C(_04429_),
    .Y(_04431_));
 sky130_fd_sc_hd__nand3_4 _34539_ (.A(_04430_),
    .B(_04405_),
    .C(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__a21o_4 _34540_ (.A1(_24050_),
    .A2(_18511_),
    .B1(_20842_),
    .X(_04433_));
 sky130_fd_sc_hd__a22oi_4 _34541_ (.A1(_04352_),
    .A2(\timer[27] ),
    .B1(_04353_),
    .B2(\irq_mask[27] ),
    .Y(_04434_));
 sky130_fd_sc_hd__nand3_4 _34542_ (.A(_04433_),
    .B(_04380_),
    .C(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__buf_1 _34543_ (.A(_03680_),
    .X(_04436_));
 sky130_fd_sc_hd__nand4_4 _34544_ (.A(_04412_),
    .B(_04413_),
    .C(_04383_),
    .D(\count_cycle[27] ),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_4 _34545_ (.A(_04358_),
    .B(\count_instr[59] ),
    .Y(_04438_));
 sky130_fd_sc_hd__a22oi_4 _34546_ (.A1(_04360_),
    .A2(\count_instr[27] ),
    .B1(_04386_),
    .B2(\count_cycle[59] ),
    .Y(_04439_));
 sky130_fd_sc_hd__a41oi_4 _34547_ (.A1(_04436_),
    .A2(_04437_),
    .A3(_04438_),
    .A4(_04439_),
    .B1(_04389_),
    .Y(_04440_));
 sky130_fd_sc_hd__nand3_4 _34548_ (.A(_04365_),
    .B(_04366_),
    .C(mem_rdata[27]),
    .Y(_04441_));
 sky130_fd_sc_hd__a21oi_4 _34549_ (.A1(_04364_),
    .A2(_04441_),
    .B1(_04368_),
    .Y(_04442_));
 sky130_fd_sc_hd__o21a_4 _34550_ (.A1(_04394_),
    .A2(\pcpi_mul.rd[27] ),
    .B1(_04423_),
    .X(_04443_));
 sky130_fd_sc_hd__o21a_4 _34551_ (.A1(_04393_),
    .A2(\pcpi_mul.rd[59] ),
    .B1(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__a2111oi_4 _34552_ (.A1(_04435_),
    .A2(_04440_),
    .B1(_04420_),
    .C1(_04442_),
    .D1(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__a22oi_4 _34553_ (.A1(_22018_),
    .A2(_04344_),
    .B1(_04432_),
    .B2(_04445_),
    .Y(_24272_));
 sky130_fd_sc_hd__buf_1 _34554_ (.A(_04143_),
    .X(_04446_));
 sky130_fd_sc_hd__xnor2_4 _34555_ (.A(_21326_),
    .B(_21850_),
    .Y(_04447_));
 sky130_fd_sc_hd__and2_4 _34556_ (.A(_04428_),
    .B(_04398_),
    .X(_04448_));
 sky130_vsdinv _34557_ (.A(_04427_),
    .Y(_04449_));
 sky130_fd_sc_hd__maj3_4 _34558_ (.A(_21321_),
    .B(_04449_),
    .C(_21828_),
    .X(_04450_));
 sky130_fd_sc_hd__a21oi_4 _34559_ (.A1(_04403_),
    .A2(_04448_),
    .B1(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__o21ai_4 _34560_ (.A1(_04447_),
    .A2(_04451_),
    .B1(_04055_),
    .Y(_04452_));
 sky130_fd_sc_hd__a21o_4 _34561_ (.A1(_04447_),
    .A2(_04451_),
    .B1(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__a2111o_4 _34562_ (.A1(_20859_),
    .A2(_20873_),
    .B1(_04408_),
    .C1(_20882_),
    .D1(_04350_),
    .X(_04454_));
 sky130_fd_sc_hd__buf_1 _34563_ (.A(_19163_),
    .X(_04455_));
 sky130_fd_sc_hd__buf_1 _34564_ (.A(_21016_),
    .X(_04456_));
 sky130_fd_sc_hd__a22oi_4 _34565_ (.A1(_04455_),
    .A2(_20884_),
    .B1(_04456_),
    .B2(\irq_mask[28] ),
    .Y(_04457_));
 sky130_fd_sc_hd__nand3_4 _34566_ (.A(_04454_),
    .B(_04380_),
    .C(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand4_4 _34567_ (.A(_04412_),
    .B(_04413_),
    .C(_04383_),
    .D(\count_cycle[28] ),
    .Y(_04459_));
 sky130_fd_sc_hd__buf_1 _34568_ (.A(_03684_),
    .X(_04460_));
 sky130_fd_sc_hd__nand2_4 _34569_ (.A(_04460_),
    .B(\count_instr[60] ),
    .Y(_04461_));
 sky130_fd_sc_hd__buf_1 _34570_ (.A(_03688_),
    .X(_04462_));
 sky130_fd_sc_hd__a22oi_4 _34571_ (.A1(_04462_),
    .A2(\count_instr[28] ),
    .B1(_04386_),
    .B2(\count_cycle[60] ),
    .Y(_04463_));
 sky130_fd_sc_hd__a41oi_4 _34572_ (.A1(_04436_),
    .A2(_04459_),
    .A3(_04461_),
    .A4(_04463_),
    .B1(_04389_),
    .Y(_04464_));
 sky130_fd_sc_hd__buf_1 _34573_ (.A(_04166_),
    .X(_04465_));
 sky130_fd_sc_hd__buf_1 _34574_ (.A(_01484_),
    .X(_04466_));
 sky130_fd_sc_hd__buf_1 _34575_ (.A(_24240_),
    .X(_04467_));
 sky130_fd_sc_hd__nand3_4 _34576_ (.A(_04466_),
    .B(_04467_),
    .C(mem_rdata[28]),
    .Y(_04468_));
 sky130_fd_sc_hd__buf_1 _34577_ (.A(_04137_),
    .X(_04469_));
 sky130_fd_sc_hd__a21oi_4 _34578_ (.A1(_04465_),
    .A2(_04468_),
    .B1(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__o21a_4 _34579_ (.A1(_04394_),
    .A2(\pcpi_mul.rd[28] ),
    .B1(_04423_),
    .X(_04471_));
 sky130_fd_sc_hd__o21a_4 _34580_ (.A1(_04393_),
    .A2(\pcpi_mul.rd[60] ),
    .B1(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__a2111oi_4 _34581_ (.A1(_04458_),
    .A2(_04464_),
    .B1(_04420_),
    .C1(_04470_),
    .D1(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__a22oi_4 _34582_ (.A1(_22010_),
    .A2(_04446_),
    .B1(_04453_),
    .B2(_04473_),
    .Y(_24273_));
 sky130_fd_sc_hd__xor2_4 _34583_ (.A(_21331_),
    .B(_21865_),
    .X(_04474_));
 sky130_fd_sc_hd__nor2_4 _34584_ (.A(\decoded_imm[28] ),
    .B(_02194_),
    .Y(_04475_));
 sky130_fd_sc_hd__nand2_4 _34585_ (.A(_21326_),
    .B(_02194_),
    .Y(_04476_));
 sky130_fd_sc_hd__o21ai_4 _34586_ (.A1(_04475_),
    .A2(_04451_),
    .B1(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__a21oi_4 _34587_ (.A1(_04477_),
    .A2(_04474_),
    .B1(_19038_),
    .Y(_04478_));
 sky130_fd_sc_hd__o21ai_4 _34588_ (.A1(_04474_),
    .A2(_04477_),
    .B1(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__a2111o_4 _34589_ (.A1(_20908_),
    .A2(_20922_),
    .B1(_04408_),
    .C1(_20929_),
    .D1(_03780_),
    .X(_04480_));
 sky130_fd_sc_hd__a22oi_4 _34590_ (.A1(_04455_),
    .A2(_20890_),
    .B1(_04456_),
    .B2(\irq_mask[29] ),
    .Y(_04481_));
 sky130_fd_sc_hd__nand3_4 _34591_ (.A(_04480_),
    .B(_03782_),
    .C(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__nand4_4 _34592_ (.A(_04412_),
    .B(_04413_),
    .C(_24094_),
    .D(\count_cycle[29] ),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_4 _34593_ (.A(_04460_),
    .B(_23439_),
    .Y(_04484_));
 sky130_fd_sc_hd__a22oi_4 _34594_ (.A1(_04462_),
    .A2(\count_instr[29] ),
    .B1(_03691_),
    .B2(\count_cycle[61] ),
    .Y(_04485_));
 sky130_fd_sc_hd__a41oi_4 _34595_ (.A1(_04436_),
    .A2(_04483_),
    .A3(_04484_),
    .A4(_04485_),
    .B1(_21215_),
    .Y(_04486_));
 sky130_fd_sc_hd__nand3_4 _34596_ (.A(_04466_),
    .B(_04467_),
    .C(mem_rdata[29]),
    .Y(_04487_));
 sky130_fd_sc_hd__a21oi_4 _34597_ (.A1(_04465_),
    .A2(_04487_),
    .B1(_04469_),
    .Y(_04488_));
 sky130_fd_sc_hd__o21a_4 _34598_ (.A1(_03743_),
    .A2(\pcpi_mul.rd[29] ),
    .B1(_04423_),
    .X(_04489_));
 sky130_fd_sc_hd__o21a_4 _34599_ (.A1(_03741_),
    .A2(\pcpi_mul.rd[61] ),
    .B1(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__a2111oi_4 _34600_ (.A1(_04482_),
    .A2(_04486_),
    .B1(_04420_),
    .C1(_04488_),
    .D1(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__a22oi_4 _34601_ (.A1(_22011_),
    .A2(_04446_),
    .B1(_04479_),
    .B2(_04491_),
    .Y(_24274_));
 sky130_fd_sc_hd__nor2_4 _34602_ (.A(_21330_),
    .B(_21864_),
    .Y(_04492_));
 sky130_vsdinv _34603_ (.A(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2_4 _34604_ (.A(_04477_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__nand2_4 _34605_ (.A(_21331_),
    .B(_21865_),
    .Y(_04495_));
 sky130_fd_sc_hd__xnor2_4 _34606_ (.A(\decoded_imm[30] ),
    .B(_21887_),
    .Y(_04496_));
 sky130_fd_sc_hd__a21o_4 _34607_ (.A1(_04494_),
    .A2(_04495_),
    .B1(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__nand3_4 _34608_ (.A(_04494_),
    .B(_04495_),
    .C(_04496_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand3_4 _34609_ (.A(_04497_),
    .B(_04405_),
    .C(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__a2111o_4 _34610_ (.A1(_20948_),
    .A2(_20962_),
    .B1(_04408_),
    .C1(_20969_),
    .D1(_03780_),
    .X(_04500_));
 sky130_fd_sc_hd__a22oi_4 _34611_ (.A1(_04455_),
    .A2(\timer[30] ),
    .B1(_04456_),
    .B2(\irq_mask[30] ),
    .Y(_04501_));
 sky130_fd_sc_hd__nand3_4 _34612_ (.A(_04500_),
    .B(_03782_),
    .C(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand4_4 _34613_ (.A(_24086_),
    .B(_24073_),
    .C(_24094_),
    .D(\count_cycle[30] ),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_4 _34614_ (.A(_04460_),
    .B(\count_instr[62] ),
    .Y(_04504_));
 sky130_fd_sc_hd__a22oi_4 _34615_ (.A1(_04462_),
    .A2(\count_instr[30] ),
    .B1(_03691_),
    .B2(\count_cycle[62] ),
    .Y(_04505_));
 sky130_fd_sc_hd__a41oi_4 _34616_ (.A1(_04436_),
    .A2(_04503_),
    .A3(_04504_),
    .A4(_04505_),
    .B1(_21215_),
    .Y(_04506_));
 sky130_fd_sc_hd__nand3_4 _34617_ (.A(_04466_),
    .B(_04467_),
    .C(mem_rdata[30]),
    .Y(_04507_));
 sky130_fd_sc_hd__a21oi_4 _34618_ (.A1(_04465_),
    .A2(_04507_),
    .B1(_04469_),
    .Y(_04508_));
 sky130_fd_sc_hd__o21a_4 _34619_ (.A1(_03743_),
    .A2(\pcpi_mul.rd[30] ),
    .B1(_18502_),
    .X(_04509_));
 sky130_fd_sc_hd__o21a_4 _34620_ (.A1(_03741_),
    .A2(\pcpi_mul.rd[62] ),
    .B1(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__a2111oi_4 _34621_ (.A1(_04502_),
    .A2(_04506_),
    .B1(_03866_),
    .C1(_04508_),
    .D1(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__a22oi_4 _34622_ (.A1(_22012_),
    .A2(_04446_),
    .B1(_04499_),
    .B2(_04511_),
    .Y(_24276_));
 sky130_fd_sc_hd__nand2_4 _34623_ (.A(_21336_),
    .B(_21887_),
    .Y(_04512_));
 sky130_vsdinv _34624_ (.A(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__a21oi_4 _34625_ (.A1(_04494_),
    .A2(_04495_),
    .B1(_04496_),
    .Y(_04514_));
 sky130_fd_sc_hd__xor2_4 _34626_ (.A(\decoded_imm[31] ),
    .B(_21900_),
    .X(_04515_));
 sky130_fd_sc_hd__o21ai_4 _34627_ (.A1(_04513_),
    .A2(_04514_),
    .B1(_04515_),
    .Y(_04516_));
 sky130_vsdinv _34628_ (.A(_04515_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand3_4 _34629_ (.A(_04497_),
    .B(_04512_),
    .C(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__nand3_4 _34630_ (.A(_04516_),
    .B(_04405_),
    .C(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__a2111o_4 _34631_ (.A1(_20991_),
    .A2(_21005_),
    .B1(_20030_),
    .C1(_21012_),
    .D1(_03780_),
    .X(_04520_));
 sky130_fd_sc_hd__a22oi_4 _34632_ (.A1(_04455_),
    .A2(\timer[31] ),
    .B1(_04456_),
    .B2(\irq_mask[31] ),
    .Y(_04521_));
 sky130_fd_sc_hd__nand3_4 _34633_ (.A(_04520_),
    .B(_03782_),
    .C(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__buf_1 _34634_ (.A(\count_cycle[31] ),
    .X(_04523_));
 sky130_fd_sc_hd__nand4_4 _34635_ (.A(_24086_),
    .B(_24073_),
    .C(_24094_),
    .D(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__nand2_4 _34636_ (.A(_04460_),
    .B(\count_instr[63] ),
    .Y(_04525_));
 sky130_fd_sc_hd__a22oi_4 _34637_ (.A1(_04462_),
    .A2(\count_instr[31] ),
    .B1(_03691_),
    .B2(\count_cycle[63] ),
    .Y(_04526_));
 sky130_fd_sc_hd__a41oi_4 _34638_ (.A1(_03681_),
    .A2(_04524_),
    .A3(_04525_),
    .A4(_04526_),
    .B1(_21215_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand3_4 _34639_ (.A(_04466_),
    .B(_04467_),
    .C(mem_rdata[31]),
    .Y(_04528_));
 sky130_fd_sc_hd__a21oi_4 _34640_ (.A1(_04465_),
    .A2(_04528_),
    .B1(_04469_),
    .Y(_04529_));
 sky130_fd_sc_hd__o21a_4 _34641_ (.A1(_03743_),
    .A2(\pcpi_mul.rd[31] ),
    .B1(_18502_),
    .X(_04530_));
 sky130_fd_sc_hd__o21a_4 _34642_ (.A1(_03741_),
    .A2(\pcpi_mul.rd[63] ),
    .B1(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__a2111oi_4 _34643_ (.A1(_04522_),
    .A2(_04527_),
    .B1(_03866_),
    .C1(_04529_),
    .D1(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__a22oi_4 _34644_ (.A1(_22013_),
    .A2(_04446_),
    .B1(_04519_),
    .B2(_04532_),
    .Y(_24277_));
 sky130_fd_sc_hd__nor4_4 _34645_ (.A(instr_xor),
    .B(instr_xori),
    .C(is_compare),
    .D(_18338_),
    .Y(_04533_));
 sky130_fd_sc_hd__nor2_4 _34646_ (.A(instr_sll),
    .B(instr_slli),
    .Y(_04534_));
 sky130_fd_sc_hd__nor2_4 _34647_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04535_));
 sky130_fd_sc_hd__nor2_4 _34648_ (.A(instr_and),
    .B(instr_andi),
    .Y(_04536_));
 sky130_fd_sc_hd__nand3_4 _34649_ (.A(_04534_),
    .B(_04535_),
    .C(_04536_),
    .Y(_04537_));
 sky130_vsdinv _34650_ (.A(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__and2_4 _34651_ (.A(_04533_),
    .B(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__buf_1 _34652_ (.A(_04539_),
    .X(_04540_));
 sky130_vsdinv _34653_ (.A(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_4 _34654_ (.A(\alu_add_sub[0] ),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__buf_1 _34655_ (.A(_18338_),
    .X(_04543_));
 sky130_fd_sc_hd__buf_1 _34656_ (.A(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__buf_1 _34657_ (.A(_18333_),
    .X(_04545_));
 sky130_fd_sc_hd__buf_1 _34658_ (.A(_18634_),
    .X(_04546_));
 sky130_fd_sc_hd__buf_1 _34659_ (.A(_04535_),
    .X(_04547_));
 sky130_fd_sc_hd__o21a_4 _34660_ (.A1(_04545_),
    .A2(_04546_),
    .B1(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__nor2_4 _34661_ (.A(_18632_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__buf_1 _34662_ (.A(_04536_),
    .X(_04550_));
 sky130_vsdinv _34663_ (.A(_04534_),
    .Y(_04551_));
 sky130_fd_sc_hd__a2bb2o_4 _34664_ (.A1_N(_18633_),
    .A2_N(_04550_),
    .B1(\alu_shl[0] ),
    .B2(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__a2111o_4 _34665_ (.A1(\alu_shr[0] ),
    .A2(_04544_),
    .B1(_04549_),
    .C1(_04552_),
    .D1(_04540_),
    .X(_04553_));
 sky130_fd_sc_hd__a21oi_4 _34666_ (.A1(is_compare),
    .A2(_19046_),
    .B1(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__nor2_4 _34667_ (.A(_04542_),
    .B(_04554_),
    .Y(\alu_out[0] ));
 sky130_fd_sc_hd__buf_1 _34668_ (.A(_18338_),
    .X(_04555_));
 sky130_fd_sc_hd__buf_1 _34669_ (.A(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__buf_1 _34670_ (.A(_04536_),
    .X(_04557_));
 sky130_fd_sc_hd__buf_1 _34671_ (.A(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__nor2_4 _34672_ (.A(_18625_),
    .B(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__buf_1 _34673_ (.A(instr_sll),
    .X(_04560_));
 sky130_fd_sc_hd__buf_1 _34674_ (.A(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__buf_1 _34675_ (.A(instr_slli),
    .X(_04562_));
 sky130_fd_sc_hd__buf_1 _34676_ (.A(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__o21a_4 _34677_ (.A1(_04561_),
    .A2(_04563_),
    .B1(\alu_shl[1] ),
    .X(_04564_));
 sky130_fd_sc_hd__buf_1 _34678_ (.A(_04545_),
    .X(_04565_));
 sky130_fd_sc_hd__buf_1 _34679_ (.A(_04547_),
    .X(_04566_));
 sky130_fd_sc_hd__o21a_4 _34680_ (.A1(_04565_),
    .A2(_18626_),
    .B1(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__nor2_4 _34681_ (.A(_18624_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__a2111oi_4 _34682_ (.A1(_04556_),
    .A2(\alu_shr[1] ),
    .B1(_04559_),
    .C1(_04564_),
    .D1(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__buf_1 _34683_ (.A(_04539_),
    .X(_04570_));
 sky130_fd_sc_hd__buf_1 _34684_ (.A(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__buf_1 _34685_ (.A(_04533_),
    .X(_04572_));
 sky130_fd_sc_hd__buf_1 _34686_ (.A(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__buf_1 _34687_ (.A(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__buf_1 _34688_ (.A(_04538_),
    .X(_04575_));
 sky130_fd_sc_hd__buf_1 _34689_ (.A(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__buf_1 _34690_ (.A(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__nand3_4 _34691_ (.A(_04574_),
    .B(\alu_add_sub[1] ),
    .C(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__o21ai_4 _34692_ (.A1(_04569_),
    .A2(_04571_),
    .B1(_04578_),
    .Y(\alu_out[1] ));
 sky130_fd_sc_hd__nor2_4 _34693_ (.A(_18616_),
    .B(_04558_),
    .Y(_04579_));
 sky130_fd_sc_hd__o21a_4 _34694_ (.A1(_04561_),
    .A2(_04563_),
    .B1(\alu_shl[2] ),
    .X(_04580_));
 sky130_fd_sc_hd__o21a_4 _34695_ (.A1(_04565_),
    .A2(_18617_),
    .B1(_04566_),
    .X(_04581_));
 sky130_fd_sc_hd__nor2_4 _34696_ (.A(_18615_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__a2111oi_4 _34697_ (.A1(_04556_),
    .A2(\alu_shr[2] ),
    .B1(_04579_),
    .C1(_04580_),
    .D1(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand3_4 _34698_ (.A(_04574_),
    .B(\alu_add_sub[2] ),
    .C(_04577_),
    .Y(_04584_));
 sky130_fd_sc_hd__o21ai_4 _34699_ (.A1(_04583_),
    .A2(_04571_),
    .B1(_04584_),
    .Y(\alu_out[2] ));
 sky130_fd_sc_hd__nor2_4 _34700_ (.A(_18610_),
    .B(_04558_),
    .Y(_04585_));
 sky130_fd_sc_hd__buf_1 _34701_ (.A(_04560_),
    .X(_04586_));
 sky130_fd_sc_hd__buf_1 _34702_ (.A(_04562_),
    .X(_04587_));
 sky130_fd_sc_hd__o21a_4 _34703_ (.A1(_04586_),
    .A2(_04587_),
    .B1(\alu_shl[3] ),
    .X(_04588_));
 sky130_fd_sc_hd__o21a_4 _34704_ (.A1(_04565_),
    .A2(_18611_),
    .B1(_04566_),
    .X(_04589_));
 sky130_fd_sc_hd__nor2_4 _34705_ (.A(_18609_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__a2111oi_4 _34706_ (.A1(_04556_),
    .A2(\alu_shr[3] ),
    .B1(_04585_),
    .C1(_04588_),
    .D1(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand3_4 _34707_ (.A(_04574_),
    .B(\alu_add_sub[3] ),
    .C(_04577_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_4 _34708_ (.A1(_04591_),
    .A2(_04571_),
    .B1(_04592_),
    .Y(\alu_out[3] ));
 sky130_fd_sc_hd__nor2_4 _34709_ (.A(_18604_),
    .B(_04558_),
    .Y(_04593_));
 sky130_fd_sc_hd__o21a_4 _34710_ (.A1(_04586_),
    .A2(_04587_),
    .B1(\alu_shl[4] ),
    .X(_04594_));
 sky130_fd_sc_hd__buf_1 _34711_ (.A(_04547_),
    .X(_04595_));
 sky130_fd_sc_hd__o21a_4 _34712_ (.A1(_04565_),
    .A2(_18605_),
    .B1(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__nor2_4 _34713_ (.A(_18603_),
    .B(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__a2111oi_4 _34714_ (.A1(_04556_),
    .A2(\alu_shr[4] ),
    .B1(_04593_),
    .C1(_04594_),
    .D1(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand3_4 _34715_ (.A(_04574_),
    .B(\alu_add_sub[4] ),
    .C(_04577_),
    .Y(_04599_));
 sky130_fd_sc_hd__o21ai_4 _34716_ (.A1(_04598_),
    .A2(_04571_),
    .B1(_04599_),
    .Y(\alu_out[4] ));
 sky130_fd_sc_hd__buf_1 _34717_ (.A(_04555_),
    .X(_04600_));
 sky130_fd_sc_hd__buf_1 _34718_ (.A(_04550_),
    .X(_04601_));
 sky130_fd_sc_hd__buf_1 _34719_ (.A(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__nor2_4 _34720_ (.A(_18585_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__buf_1 _34721_ (.A(instr_xor),
    .X(_04604_));
 sky130_fd_sc_hd__buf_1 _34722_ (.A(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__buf_1 _34723_ (.A(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__buf_1 _34724_ (.A(instr_xori),
    .X(_04607_));
 sky130_fd_sc_hd__buf_1 _34725_ (.A(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__buf_1 _34726_ (.A(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__o21ai_4 _34727_ (.A1(_04606_),
    .A2(_04609_),
    .B1(_18585_),
    .Y(_04610_));
 sky130_fd_sc_hd__buf_1 _34728_ (.A(_04535_),
    .X(_04611_));
 sky130_fd_sc_hd__buf_1 _34729_ (.A(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__a21oi_4 _34730_ (.A1(_04610_),
    .A2(_04612_),
    .B1(_18584_),
    .Y(_04613_));
 sky130_fd_sc_hd__buf_1 _34731_ (.A(instr_sll),
    .X(_04614_));
 sky130_fd_sc_hd__buf_1 _34732_ (.A(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__o21a_4 _34733_ (.A1(_04615_),
    .A2(_24110_),
    .B1(\alu_shl[5] ),
    .X(_04616_));
 sky130_fd_sc_hd__a2111oi_4 _34734_ (.A1(_04600_),
    .A2(\alu_shr[5] ),
    .B1(_04603_),
    .C1(_04613_),
    .D1(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__buf_1 _34735_ (.A(_04539_),
    .X(_04618_));
 sky130_fd_sc_hd__buf_1 _34736_ (.A(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__buf_1 _34737_ (.A(_04572_),
    .X(_04620_));
 sky130_fd_sc_hd__buf_1 _34738_ (.A(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__buf_1 _34739_ (.A(_04575_),
    .X(_04622_));
 sky130_fd_sc_hd__buf_1 _34740_ (.A(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__nand3_4 _34741_ (.A(_04621_),
    .B(\alu_add_sub[5] ),
    .C(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__o21ai_4 _34742_ (.A1(_04617_),
    .A2(_04619_),
    .B1(_04624_),
    .Y(\alu_out[5] ));
 sky130_fd_sc_hd__nor2_4 _34743_ (.A(_18597_),
    .B(_04602_),
    .Y(_04625_));
 sky130_fd_sc_hd__o21ai_4 _34744_ (.A1(_04606_),
    .A2(_04609_),
    .B1(_18597_),
    .Y(_04626_));
 sky130_fd_sc_hd__buf_1 _34745_ (.A(_04547_),
    .X(_04627_));
 sky130_fd_sc_hd__buf_1 _34746_ (.A(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__a21oi_4 _34747_ (.A1(_04626_),
    .A2(_04628_),
    .B1(_18596_),
    .Y(_04629_));
 sky130_fd_sc_hd__o21a_4 _34748_ (.A1(_04615_),
    .A2(_24110_),
    .B1(\alu_shl[6] ),
    .X(_04630_));
 sky130_fd_sc_hd__a2111oi_4 _34749_ (.A1(_04600_),
    .A2(\alu_shr[6] ),
    .B1(_04625_),
    .C1(_04629_),
    .D1(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__nand3_4 _34750_ (.A(_04621_),
    .B(\alu_add_sub[6] ),
    .C(_04623_),
    .Y(_04632_));
 sky130_fd_sc_hd__o21ai_4 _34751_ (.A1(_04631_),
    .A2(_04619_),
    .B1(_04632_),
    .Y(\alu_out[6] ));
 sky130_fd_sc_hd__nor2_4 _34752_ (.A(_18590_),
    .B(_04602_),
    .Y(_04633_));
 sky130_fd_sc_hd__o21a_4 _34753_ (.A1(_04586_),
    .A2(_04587_),
    .B1(\alu_shl[7] ),
    .X(_04634_));
 sky130_fd_sc_hd__buf_1 _34754_ (.A(_18333_),
    .X(_04635_));
 sky130_fd_sc_hd__o21a_4 _34755_ (.A1(_04635_),
    .A2(_18591_),
    .B1(_04595_),
    .X(_04636_));
 sky130_fd_sc_hd__nor2_4 _34756_ (.A(_18592_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__a2111oi_4 _34757_ (.A1(_04600_),
    .A2(\alu_shr[7] ),
    .B1(_04633_),
    .C1(_04634_),
    .D1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand3_4 _34758_ (.A(_04621_),
    .B(\alu_add_sub[7] ),
    .C(_04623_),
    .Y(_04639_));
 sky130_fd_sc_hd__o21ai_4 _34759_ (.A1(_04638_),
    .A2(_04619_),
    .B1(_04639_),
    .Y(\alu_out[7] ));
 sky130_fd_sc_hd__nand2_4 _34760_ (.A(_21507_),
    .B(_24236_),
    .Y(_04640_));
 sky130_fd_sc_hd__nor2_4 _34761_ (.A(_04640_),
    .B(_04602_),
    .Y(_04641_));
 sky130_fd_sc_hd__o21a_4 _34762_ (.A1(_04586_),
    .A2(_04587_),
    .B1(\alu_shl[8] ),
    .X(_04642_));
 sky130_fd_sc_hd__buf_1 _34763_ (.A(_04605_),
    .X(_04643_));
 sky130_fd_sc_hd__buf_1 _34764_ (.A(_04608_),
    .X(_04644_));
 sky130_fd_sc_hd__o21ai_4 _34765_ (.A1(_04643_),
    .A2(_04644_),
    .B1(_04640_),
    .Y(_04645_));
 sky130_fd_sc_hd__a22oi_4 _34766_ (.A1(_21506_),
    .A2(_21204_),
    .B1(_04645_),
    .B2(_04612_),
    .Y(_04646_));
 sky130_fd_sc_hd__a2111oi_4 _34767_ (.A1(_04600_),
    .A2(\alu_shr[8] ),
    .B1(_04641_),
    .C1(_04642_),
    .D1(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__nand3_4 _34768_ (.A(_04621_),
    .B(\alu_add_sub[8] ),
    .C(_04623_),
    .Y(_04648_));
 sky130_fd_sc_hd__o21ai_4 _34769_ (.A1(_04647_),
    .A2(_04619_),
    .B1(_04648_),
    .Y(\alu_out[8] ));
 sky130_fd_sc_hd__buf_1 _34770_ (.A(_04555_),
    .X(_04649_));
 sky130_fd_sc_hd__nand2_4 _34771_ (.A(_21530_),
    .B(_24243_),
    .Y(_04650_));
 sky130_fd_sc_hd__buf_1 _34772_ (.A(_04601_),
    .X(_04651_));
 sky130_fd_sc_hd__nor2_4 _34773_ (.A(_04650_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__buf_1 _34774_ (.A(_04604_),
    .X(_04653_));
 sky130_fd_sc_hd__buf_1 _34775_ (.A(_04607_),
    .X(_04654_));
 sky130_fd_sc_hd__o21ai_4 _34776_ (.A1(_04653_),
    .A2(_04654_),
    .B1(_04650_),
    .Y(_04655_));
 sky130_fd_sc_hd__buf_1 _34777_ (.A(_04627_),
    .X(_04656_));
 sky130_fd_sc_hd__a22oi_4 _34778_ (.A1(_21529_),
    .A2(_21211_),
    .B1(_04655_),
    .B2(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__o21a_4 _34779_ (.A1(_04615_),
    .A2(_24110_),
    .B1(\alu_shl[9] ),
    .X(_04658_));
 sky130_fd_sc_hd__a2111oi_4 _34780_ (.A1(_04649_),
    .A2(\alu_shr[9] ),
    .B1(_04652_),
    .C1(_04657_),
    .D1(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__buf_1 _34781_ (.A(_04618_),
    .X(_04660_));
 sky130_fd_sc_hd__buf_1 _34782_ (.A(_04620_),
    .X(_04661_));
 sky130_fd_sc_hd__buf_1 _34783_ (.A(_04622_),
    .X(_04662_));
 sky130_fd_sc_hd__nand3_4 _34784_ (.A(_04661_),
    .B(\alu_add_sub[9] ),
    .C(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__o21ai_4 _34785_ (.A1(_04659_),
    .A2(_04660_),
    .B1(_04663_),
    .Y(\alu_out[9] ));
 sky130_fd_sc_hd__nand2_4 _34786_ (.A(_01611_),
    .B(_21227_),
    .Y(_04664_));
 sky130_fd_sc_hd__nor2_4 _34787_ (.A(_04664_),
    .B(_04651_),
    .Y(_04665_));
 sky130_fd_sc_hd__buf_1 _34788_ (.A(_04560_),
    .X(_04666_));
 sky130_fd_sc_hd__buf_1 _34789_ (.A(_04562_),
    .X(_04667_));
 sky130_fd_sc_hd__o21a_4 _34790_ (.A1(_04666_),
    .A2(_04667_),
    .B1(\alu_shl[10] ),
    .X(_04668_));
 sky130_fd_sc_hd__o21ai_4 _34791_ (.A1(_04605_),
    .A2(_04608_),
    .B1(_04664_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand2_4 _34792_ (.A(_04669_),
    .B(_04566_),
    .Y(_04670_));
 sky130_fd_sc_hd__o21a_4 _34793_ (.A1(_01611_),
    .A2(_21228_),
    .B1(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__a2111oi_4 _34794_ (.A1(_04649_),
    .A2(\alu_shr[10] ),
    .B1(_04665_),
    .C1(_04668_),
    .D1(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__nand3_4 _34795_ (.A(_04661_),
    .B(\alu_add_sub[10] ),
    .C(_04662_),
    .Y(_04673_));
 sky130_fd_sc_hd__o21ai_4 _34796_ (.A1(_04672_),
    .A2(_04660_),
    .B1(_04673_),
    .Y(\alu_out[10] ));
 sky130_fd_sc_hd__nand2_4 _34797_ (.A(_21565_),
    .B(_24248_),
    .Y(_04674_));
 sky130_fd_sc_hd__nor2_4 _34798_ (.A(_04674_),
    .B(_04651_),
    .Y(_04675_));
 sky130_fd_sc_hd__o21a_4 _34799_ (.A1(_04666_),
    .A2(_04667_),
    .B1(\alu_shl[11] ),
    .X(_04676_));
 sky130_fd_sc_hd__o21ai_4 _34800_ (.A1(_04643_),
    .A2(_04644_),
    .B1(_04674_),
    .Y(_04677_));
 sky130_fd_sc_hd__a22oi_4 _34801_ (.A1(_21564_),
    .A2(_21230_),
    .B1(_04677_),
    .B2(_04612_),
    .Y(_04678_));
 sky130_fd_sc_hd__a2111oi_4 _34802_ (.A1(_04649_),
    .A2(\alu_shr[11] ),
    .B1(_04675_),
    .C1(_04676_),
    .D1(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__nand3_4 _34803_ (.A(_04661_),
    .B(\alu_add_sub[11] ),
    .C(_04662_),
    .Y(_04680_));
 sky130_fd_sc_hd__o21ai_4 _34804_ (.A1(_04679_),
    .A2(_04660_),
    .B1(_04680_),
    .Y(\alu_out[11] ));
 sky130_fd_sc_hd__nand2_4 _34805_ (.A(_21590_),
    .B(_24252_),
    .Y(_04681_));
 sky130_fd_sc_hd__nor2_4 _34806_ (.A(_04681_),
    .B(_04651_),
    .Y(_04682_));
 sky130_fd_sc_hd__buf_1 _34807_ (.A(_04604_),
    .X(_04683_));
 sky130_fd_sc_hd__buf_1 _34808_ (.A(_04607_),
    .X(_04684_));
 sky130_fd_sc_hd__o21ai_4 _34809_ (.A1(_04683_),
    .A2(_04684_),
    .B1(_04681_),
    .Y(_04685_));
 sky130_fd_sc_hd__a22oi_4 _34810_ (.A1(_21580_),
    .A2(_21236_),
    .B1(_04685_),
    .B2(_04656_),
    .Y(_04686_));
 sky130_fd_sc_hd__buf_1 _34811_ (.A(_04614_),
    .X(_04687_));
 sky130_fd_sc_hd__buf_1 _34812_ (.A(_24109_),
    .X(_04688_));
 sky130_fd_sc_hd__o21a_4 _34813_ (.A1(_04687_),
    .A2(_04688_),
    .B1(\alu_shl[12] ),
    .X(_04689_));
 sky130_fd_sc_hd__a2111oi_4 _34814_ (.A1(_04649_),
    .A2(\alu_shr[12] ),
    .B1(_04682_),
    .C1(_04686_),
    .D1(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand3_4 _34815_ (.A(_04661_),
    .B(\alu_add_sub[12] ),
    .C(_04662_),
    .Y(_04691_));
 sky130_fd_sc_hd__o21ai_4 _34816_ (.A1(_04690_),
    .A2(_04660_),
    .B1(_04691_),
    .Y(\alu_out[12] ));
 sky130_fd_sc_hd__buf_1 _34817_ (.A(_04555_),
    .X(_04692_));
 sky130_fd_sc_hd__nand2_4 _34818_ (.A(_21605_),
    .B(_01476_),
    .Y(_04693_));
 sky130_fd_sc_hd__buf_1 _34819_ (.A(_04601_),
    .X(_04694_));
 sky130_fd_sc_hd__nor2_4 _34820_ (.A(_04693_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__o21ai_4 _34821_ (.A1(_04683_),
    .A2(_04684_),
    .B1(_04693_),
    .Y(_04696_));
 sky130_fd_sc_hd__buf_1 _34822_ (.A(_04627_),
    .X(_04697_));
 sky130_fd_sc_hd__a22oi_4 _34823_ (.A1(_21602_),
    .A2(_21244_),
    .B1(_04696_),
    .B2(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__o21a_4 _34824_ (.A1(_04687_),
    .A2(_04688_),
    .B1(\alu_shl[13] ),
    .X(_04699_));
 sky130_fd_sc_hd__a2111oi_4 _34825_ (.A1(_04692_),
    .A2(\alu_shr[13] ),
    .B1(_04695_),
    .C1(_04698_),
    .D1(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__buf_1 _34826_ (.A(_04618_),
    .X(_04701_));
 sky130_fd_sc_hd__buf_1 _34827_ (.A(_04620_),
    .X(_04702_));
 sky130_fd_sc_hd__buf_1 _34828_ (.A(_04622_),
    .X(_04703_));
 sky130_fd_sc_hd__nand3_4 _34829_ (.A(_04702_),
    .B(\alu_add_sub[13] ),
    .C(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__o21ai_4 _34830_ (.A1(_04700_),
    .A2(_04701_),
    .B1(_04704_),
    .Y(\alu_out[13] ));
 sky130_fd_sc_hd__nand2_4 _34831_ (.A(_01630_),
    .B(_01478_),
    .Y(_04705_));
 sky130_fd_sc_hd__nor2_4 _34832_ (.A(_04705_),
    .B(_04694_),
    .Y(_04706_));
 sky130_fd_sc_hd__o21ai_4 _34833_ (.A1(_04683_),
    .A2(_04684_),
    .B1(_04705_),
    .Y(_04707_));
 sky130_fd_sc_hd__a22oi_4 _34834_ (.A1(_21622_),
    .A2(_21250_),
    .B1(_04707_),
    .B2(_04697_),
    .Y(_04708_));
 sky130_fd_sc_hd__o21a_4 _34835_ (.A1(_04687_),
    .A2(_04688_),
    .B1(\alu_shl[14] ),
    .X(_04709_));
 sky130_fd_sc_hd__a2111oi_4 _34836_ (.A1(_04692_),
    .A2(\alu_shr[14] ),
    .B1(_04706_),
    .C1(_04708_),
    .D1(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand3_4 _34837_ (.A(_04702_),
    .B(\alu_add_sub[14] ),
    .C(_04703_),
    .Y(_04711_));
 sky130_fd_sc_hd__o21ai_4 _34838_ (.A1(_04710_),
    .A2(_04701_),
    .B1(_04711_),
    .Y(\alu_out[14] ));
 sky130_fd_sc_hd__nand2_4 _34839_ (.A(_01636_),
    .B(_01480_),
    .Y(_04712_));
 sky130_fd_sc_hd__nor2_4 _34840_ (.A(_04712_),
    .B(_04694_),
    .Y(_04713_));
 sky130_fd_sc_hd__o21ai_4 _34841_ (.A1(_04683_),
    .A2(_04684_),
    .B1(_04712_),
    .Y(_04714_));
 sky130_fd_sc_hd__a22oi_4 _34842_ (.A1(_21640_),
    .A2(_21257_),
    .B1(_04714_),
    .B2(_04697_),
    .Y(_04715_));
 sky130_fd_sc_hd__o21a_4 _34843_ (.A1(_04687_),
    .A2(_04688_),
    .B1(\alu_shl[15] ),
    .X(_04716_));
 sky130_fd_sc_hd__a2111oi_4 _34844_ (.A1(_04692_),
    .A2(\alu_shr[15] ),
    .B1(_04713_),
    .C1(_04715_),
    .D1(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__nand3_4 _34845_ (.A(_04702_),
    .B(\alu_add_sub[15] ),
    .C(_04703_),
    .Y(_04718_));
 sky130_fd_sc_hd__o21ai_4 _34846_ (.A1(_04717_),
    .A2(_04701_),
    .B1(_04718_),
    .Y(\alu_out[15] ));
 sky130_fd_sc_hd__nand2_4 _34847_ (.A(_21678_),
    .B(_18712_),
    .Y(_04719_));
 sky130_fd_sc_hd__nor2_4 _34848_ (.A(_04719_),
    .B(_04694_),
    .Y(_04720_));
 sky130_fd_sc_hd__o21a_4 _34849_ (.A1(_04666_),
    .A2(_04667_),
    .B1(\alu_shl[16] ),
    .X(_04721_));
 sky130_fd_sc_hd__o21ai_4 _34850_ (.A1(_04643_),
    .A2(_04644_),
    .B1(_04719_),
    .Y(_04722_));
 sky130_fd_sc_hd__a22oi_4 _34851_ (.A1(_21654_),
    .A2(_21262_),
    .B1(_04722_),
    .B2(_04612_),
    .Y(_04723_));
 sky130_fd_sc_hd__a2111oi_4 _34852_ (.A1(_04692_),
    .A2(\alu_shr[16] ),
    .B1(_04720_),
    .C1(_04721_),
    .D1(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__nand3_4 _34853_ (.A(_04702_),
    .B(\alu_add_sub[16] ),
    .C(_04703_),
    .Y(_04725_));
 sky130_fd_sc_hd__o21ai_4 _34854_ (.A1(_04724_),
    .A2(_04701_),
    .B1(_04725_),
    .Y(\alu_out[16] ));
 sky130_fd_sc_hd__buf_1 _34855_ (.A(_04543_),
    .X(_04726_));
 sky130_fd_sc_hd__nand2_4 _34856_ (.A(_18715_),
    .B(_18717_),
    .Y(_04727_));
 sky130_fd_sc_hd__buf_1 _34857_ (.A(_04601_),
    .X(_04728_));
 sky130_fd_sc_hd__nor2_4 _34858_ (.A(_04727_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__o21ai_4 _34859_ (.A1(_04605_),
    .A2(_04608_),
    .B1(_04727_),
    .Y(_04730_));
 sky130_fd_sc_hd__a22oi_4 _34860_ (.A1(_21671_),
    .A2(_21267_),
    .B1(_04730_),
    .B2(_04697_),
    .Y(_04731_));
 sky130_fd_sc_hd__buf_1 _34861_ (.A(_04614_),
    .X(_04732_));
 sky130_fd_sc_hd__buf_1 _34862_ (.A(_24109_),
    .X(_04733_));
 sky130_fd_sc_hd__o21a_4 _34863_ (.A1(_04732_),
    .A2(_04733_),
    .B1(\alu_shl[17] ),
    .X(_04734_));
 sky130_fd_sc_hd__a2111oi_4 _34864_ (.A1(_04726_),
    .A2(\alu_shr[17] ),
    .B1(_04729_),
    .C1(_04731_),
    .D1(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__buf_1 _34865_ (.A(_04618_),
    .X(_04736_));
 sky130_fd_sc_hd__buf_1 _34866_ (.A(_04620_),
    .X(_04737_));
 sky130_fd_sc_hd__buf_1 _34867_ (.A(_04622_),
    .X(_04738_));
 sky130_fd_sc_hd__nand3_4 _34868_ (.A(_04737_),
    .B(\alu_add_sub[17] ),
    .C(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__o21ai_4 _34869_ (.A1(_04735_),
    .A2(_04736_),
    .B1(_04739_),
    .Y(\alu_out[17] ));
 sky130_fd_sc_hd__nor2_4 _34870_ (.A(_18707_),
    .B(_04728_),
    .Y(_04740_));
 sky130_fd_sc_hd__buf_1 _34871_ (.A(_04604_),
    .X(_04741_));
 sky130_fd_sc_hd__buf_1 _34872_ (.A(_04607_),
    .X(_04742_));
 sky130_fd_sc_hd__o21ai_4 _34873_ (.A1(_04741_),
    .A2(_04742_),
    .B1(_18707_),
    .Y(_04743_));
 sky130_fd_sc_hd__buf_1 _34874_ (.A(_04627_),
    .X(_04744_));
 sky130_fd_sc_hd__a21boi_4 _34875_ (.A1(_04743_),
    .A2(_04744_),
    .B1_N(_18704_),
    .Y(_04745_));
 sky130_fd_sc_hd__o21a_4 _34876_ (.A1(_04732_),
    .A2(_04733_),
    .B1(\alu_shl[18] ),
    .X(_04746_));
 sky130_fd_sc_hd__a2111oi_4 _34877_ (.A1(_04726_),
    .A2(\alu_shr[18] ),
    .B1(_04740_),
    .C1(_04745_),
    .D1(_04746_),
    .Y(_04747_));
 sky130_fd_sc_hd__nand3_4 _34878_ (.A(_04737_),
    .B(\alu_add_sub[18] ),
    .C(_04738_),
    .Y(_04748_));
 sky130_fd_sc_hd__o21ai_4 _34879_ (.A1(_04747_),
    .A2(_04736_),
    .B1(_04748_),
    .Y(\alu_out[18] ));
 sky130_fd_sc_hd__nor2_4 _34880_ (.A(_18698_),
    .B(_04728_),
    .Y(_04749_));
 sky130_fd_sc_hd__o21a_4 _34881_ (.A1(_04666_),
    .A2(_04667_),
    .B1(\alu_shl[19] ),
    .X(_04750_));
 sky130_fd_sc_hd__o21a_4 _34882_ (.A1(_04635_),
    .A2(_18699_),
    .B1(_04595_),
    .X(_04751_));
 sky130_fd_sc_hd__nor2_4 _34883_ (.A(_18697_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__a2111oi_4 _34884_ (.A1(_04726_),
    .A2(\alu_shr[19] ),
    .B1(_04749_),
    .C1(_04750_),
    .D1(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand3_4 _34885_ (.A(_04737_),
    .B(\alu_add_sub[19] ),
    .C(_04738_),
    .Y(_04754_));
 sky130_fd_sc_hd__o21ai_4 _34886_ (.A1(_04753_),
    .A2(_04736_),
    .B1(_04754_),
    .Y(\alu_out[19] ));
 sky130_fd_sc_hd__nor2_4 _34887_ (.A(_18670_),
    .B(_04728_),
    .Y(_04755_));
 sky130_fd_sc_hd__buf_1 _34888_ (.A(_04560_),
    .X(_04756_));
 sky130_fd_sc_hd__buf_1 _34889_ (.A(_04562_),
    .X(_04757_));
 sky130_fd_sc_hd__o21a_4 _34890_ (.A1(_04756_),
    .A2(_04757_),
    .B1(\alu_shl[20] ),
    .X(_04758_));
 sky130_fd_sc_hd__o21a_4 _34891_ (.A1(_04635_),
    .A2(_18671_),
    .B1(_04595_),
    .X(_04759_));
 sky130_fd_sc_hd__nor2_4 _34892_ (.A(_18669_),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__a2111oi_4 _34893_ (.A1(_04726_),
    .A2(\alu_shr[20] ),
    .B1(_04755_),
    .C1(_04758_),
    .D1(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__nand3_4 _34894_ (.A(_04737_),
    .B(\alu_add_sub[20] ),
    .C(_04738_),
    .Y(_04762_));
 sky130_fd_sc_hd__o21ai_4 _34895_ (.A1(_04761_),
    .A2(_04736_),
    .B1(_04762_),
    .Y(\alu_out[20] ));
 sky130_fd_sc_hd__buf_1 _34896_ (.A(_04543_),
    .X(_04763_));
 sky130_fd_sc_hd__buf_1 _34897_ (.A(_04550_),
    .X(_04764_));
 sky130_fd_sc_hd__nor2_4 _34898_ (.A(_18684_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__o21ai_4 _34899_ (.A1(_04606_),
    .A2(_04609_),
    .B1(_18684_),
    .Y(_04766_));
 sky130_fd_sc_hd__a21oi_4 _34900_ (.A1(_04766_),
    .A2(_04628_),
    .B1(_18683_),
    .Y(_04767_));
 sky130_fd_sc_hd__o21a_4 _34901_ (.A1(_04732_),
    .A2(_04733_),
    .B1(\alu_shl[21] ),
    .X(_04768_));
 sky130_fd_sc_hd__a2111oi_4 _34902_ (.A1(_04763_),
    .A2(\alu_shr[21] ),
    .B1(_04765_),
    .C1(_04767_),
    .D1(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__buf_1 _34903_ (.A(_04540_),
    .X(_04770_));
 sky130_fd_sc_hd__buf_1 _34904_ (.A(_04572_),
    .X(_04771_));
 sky130_fd_sc_hd__buf_1 _34905_ (.A(_04575_),
    .X(_04772_));
 sky130_fd_sc_hd__nand3_4 _34906_ (.A(_04771_),
    .B(\alu_add_sub[21] ),
    .C(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__o21ai_4 _34907_ (.A1(_04769_),
    .A2(_04770_),
    .B1(_04773_),
    .Y(\alu_out[21] ));
 sky130_fd_sc_hd__nor2_4 _34908_ (.A(_18678_),
    .B(_04764_),
    .Y(_04774_));
 sky130_fd_sc_hd__o21ai_4 _34909_ (.A1(_04653_),
    .A2(_04654_),
    .B1(_18678_),
    .Y(_04775_));
 sky130_fd_sc_hd__a21boi_4 _34910_ (.A1(_04775_),
    .A2(_04744_),
    .B1_N(_18675_),
    .Y(_04776_));
 sky130_fd_sc_hd__o21a_4 _34911_ (.A1(_04732_),
    .A2(_04733_),
    .B1(\alu_shl[22] ),
    .X(_04777_));
 sky130_fd_sc_hd__a2111oi_4 _34912_ (.A1(_04763_),
    .A2(\alu_shr[22] ),
    .B1(_04774_),
    .C1(_04776_),
    .D1(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand3_4 _34913_ (.A(_04771_),
    .B(\alu_add_sub[22] ),
    .C(_04772_),
    .Y(_04779_));
 sky130_fd_sc_hd__o21ai_4 _34914_ (.A1(_04778_),
    .A2(_04770_),
    .B1(_04779_),
    .Y(\alu_out[22] ));
 sky130_fd_sc_hd__nor2_4 _34915_ (.A(_18686_),
    .B(_04764_),
    .Y(_04780_));
 sky130_fd_sc_hd__o21a_4 _34916_ (.A1(_04756_),
    .A2(_04757_),
    .B1(\alu_shl[23] ),
    .X(_04781_));
 sky130_fd_sc_hd__o21a_4 _34917_ (.A1(_04635_),
    .A2(_18687_),
    .B1(_04611_),
    .X(_04782_));
 sky130_fd_sc_hd__nor2_4 _34918_ (.A(_18690_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__a2111oi_4 _34919_ (.A1(_04763_),
    .A2(\alu_shr[23] ),
    .B1(_04780_),
    .C1(_04781_),
    .D1(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__nand3_4 _34920_ (.A(_04771_),
    .B(\alu_add_sub[23] ),
    .C(_04772_),
    .Y(_04785_));
 sky130_fd_sc_hd__o21ai_4 _34921_ (.A1(_04784_),
    .A2(_04770_),
    .B1(_04785_),
    .Y(\alu_out[23] ));
 sky130_fd_sc_hd__nor2_4 _34922_ (.A(_18735_),
    .B(_04764_),
    .Y(_04786_));
 sky130_fd_sc_hd__o21ai_4 _34923_ (.A1(_04653_),
    .A2(_04654_),
    .B1(_18735_),
    .Y(_04787_));
 sky130_fd_sc_hd__a21boi_4 _34924_ (.A1(_04787_),
    .A2(_04656_),
    .B1_N(_18730_),
    .Y(_04788_));
 sky130_fd_sc_hd__buf_1 _34925_ (.A(_04614_),
    .X(_04789_));
 sky130_fd_sc_hd__buf_1 _34926_ (.A(_24109_),
    .X(_04790_));
 sky130_fd_sc_hd__o21a_4 _34927_ (.A1(_04789_),
    .A2(_04790_),
    .B1(\alu_shl[24] ),
    .X(_04791_));
 sky130_fd_sc_hd__a2111oi_4 _34928_ (.A1(_04763_),
    .A2(\alu_shr[24] ),
    .B1(_04786_),
    .C1(_04788_),
    .D1(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand3_4 _34929_ (.A(_04771_),
    .B(\alu_add_sub[24] ),
    .C(_04772_),
    .Y(_04793_));
 sky130_fd_sc_hd__o21ai_4 _34930_ (.A1(_04792_),
    .A2(_04770_),
    .B1(_04793_),
    .Y(\alu_out[24] ));
 sky130_fd_sc_hd__buf_1 _34931_ (.A(_04543_),
    .X(_04794_));
 sky130_fd_sc_hd__buf_1 _34932_ (.A(_04550_),
    .X(_04795_));
 sky130_fd_sc_hd__nor2_4 _34933_ (.A(_18770_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__o21ai_4 _34934_ (.A1(_04606_),
    .A2(_04609_),
    .B1(_18770_),
    .Y(_04797_));
 sky130_fd_sc_hd__a21oi_4 _34935_ (.A1(_04797_),
    .A2(_04628_),
    .B1(_18768_),
    .Y(_04798_));
 sky130_fd_sc_hd__o21a_4 _34936_ (.A1(_04789_),
    .A2(_04790_),
    .B1(\alu_shl[25] ),
    .X(_04799_));
 sky130_fd_sc_hd__a2111oi_4 _34937_ (.A1(_04794_),
    .A2(\alu_shr[25] ),
    .B1(_04796_),
    .C1(_04798_),
    .D1(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__buf_1 _34938_ (.A(_04540_),
    .X(_04801_));
 sky130_fd_sc_hd__buf_1 _34939_ (.A(_04572_),
    .X(_04802_));
 sky130_fd_sc_hd__buf_1 _34940_ (.A(_04575_),
    .X(_04803_));
 sky130_fd_sc_hd__nand3_4 _34941_ (.A(_04802_),
    .B(\alu_add_sub[25] ),
    .C(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__o21ai_4 _34942_ (.A1(_04800_),
    .A2(_04801_),
    .B1(_04804_),
    .Y(\alu_out[25] ));
 sky130_fd_sc_hd__nor2_4 _34943_ (.A(_18725_),
    .B(_04795_),
    .Y(_04805_));
 sky130_fd_sc_hd__o21ai_4 _34944_ (.A1(_04741_),
    .A2(_04742_),
    .B1(_18725_),
    .Y(_04806_));
 sky130_fd_sc_hd__a21oi_4 _34945_ (.A1(_04806_),
    .A2(_04628_),
    .B1(_18723_),
    .Y(_04807_));
 sky130_fd_sc_hd__o21a_4 _34946_ (.A1(_04789_),
    .A2(_04790_),
    .B1(\alu_shl[26] ),
    .X(_04808_));
 sky130_fd_sc_hd__a2111oi_4 _34947_ (.A1(_04794_),
    .A2(\alu_shr[26] ),
    .B1(_04805_),
    .C1(_04807_),
    .D1(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__nand3_4 _34948_ (.A(_04802_),
    .B(\alu_add_sub[26] ),
    .C(_04803_),
    .Y(_04810_));
 sky130_fd_sc_hd__o21ai_4 _34949_ (.A1(_04809_),
    .A2(_04801_),
    .B1(_04810_),
    .Y(\alu_out[26] ));
 sky130_fd_sc_hd__nor2_4 _34950_ (.A(_18763_),
    .B(_04795_),
    .Y(_04811_));
 sky130_fd_sc_hd__o21ai_4 _34951_ (.A1(_04653_),
    .A2(_04654_),
    .B1(_18763_),
    .Y(_04812_));
 sky130_fd_sc_hd__a21boi_4 _34952_ (.A1(_04812_),
    .A2(_04656_),
    .B1_N(_18761_),
    .Y(_04813_));
 sky130_fd_sc_hd__o21a_4 _34953_ (.A1(_04789_),
    .A2(_04790_),
    .B1(\alu_shl[27] ),
    .X(_04814_));
 sky130_fd_sc_hd__a2111oi_4 _34954_ (.A1(_04794_),
    .A2(\alu_shr[27] ),
    .B1(_04811_),
    .C1(_04813_),
    .D1(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand3_4 _34955_ (.A(_04802_),
    .B(\alu_add_sub[27] ),
    .C(_04803_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21ai_4 _34956_ (.A1(_04815_),
    .A2(_04801_),
    .B1(_04816_),
    .Y(\alu_out[27] ));
 sky130_fd_sc_hd__nor2_4 _34957_ (.A(_18749_),
    .B(_04795_),
    .Y(_04817_));
 sky130_fd_sc_hd__o21a_4 _34958_ (.A1(_04756_),
    .A2(_04757_),
    .B1(\alu_shl[28] ),
    .X(_04818_));
 sky130_fd_sc_hd__o21a_4 _34959_ (.A1(_04545_),
    .A2(_18750_),
    .B1(_04611_),
    .X(_04819_));
 sky130_fd_sc_hd__nor2_4 _34960_ (.A(_18748_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__a2111oi_4 _34961_ (.A1(_04794_),
    .A2(\alu_shr[28] ),
    .B1(_04817_),
    .C1(_04818_),
    .D1(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__nand3_4 _34962_ (.A(_04802_),
    .B(\alu_add_sub[28] ),
    .C(_04803_),
    .Y(_04822_));
 sky130_fd_sc_hd__o21ai_4 _34963_ (.A1(_04821_),
    .A2(_04801_),
    .B1(_04822_),
    .Y(\alu_out[28] ));
 sky130_fd_sc_hd__nor2_4 _34964_ (.A(_18753_),
    .B(_04557_),
    .Y(_04823_));
 sky130_fd_sc_hd__o21ai_4 _34965_ (.A1(_04741_),
    .A2(_04742_),
    .B1(_18753_),
    .Y(_04824_));
 sky130_fd_sc_hd__a21oi_4 _34966_ (.A1(_04824_),
    .A2(_04744_),
    .B1(_18755_),
    .Y(_04825_));
 sky130_fd_sc_hd__o21a_4 _34967_ (.A1(_04561_),
    .A2(_04563_),
    .B1(\alu_shl[29] ),
    .X(_04826_));
 sky130_fd_sc_hd__a2111oi_4 _34968_ (.A1(_04544_),
    .A2(\alu_shr[29] ),
    .B1(_04823_),
    .C1(_04825_),
    .D1(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__nand3_4 _34969_ (.A(_04573_),
    .B(\alu_add_sub[29] ),
    .C(_04576_),
    .Y(_04828_));
 sky130_fd_sc_hd__o21ai_4 _34970_ (.A1(_04827_),
    .A2(_04570_),
    .B1(_04828_),
    .Y(\alu_out[29] ));
 sky130_fd_sc_hd__nor2_4 _34971_ (.A(_18739_),
    .B(_04557_),
    .Y(_04829_));
 sky130_fd_sc_hd__o21a_4 _34972_ (.A1(_04756_),
    .A2(_04757_),
    .B1(\alu_shl[30] ),
    .X(_04830_));
 sky130_fd_sc_hd__o21a_4 _34973_ (.A1(_04545_),
    .A2(_18740_),
    .B1(_04611_),
    .X(_04831_));
 sky130_fd_sc_hd__nor2_4 _34974_ (.A(_18738_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__a2111oi_4 _34975_ (.A1(_04544_),
    .A2(\alu_shr[30] ),
    .B1(_04829_),
    .C1(_04830_),
    .D1(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__nand3_4 _34976_ (.A(_04573_),
    .B(\alu_add_sub[30] ),
    .C(_04576_),
    .Y(_04834_));
 sky130_fd_sc_hd__o21ai_4 _34977_ (.A1(_04833_),
    .A2(_04570_),
    .B1(_04834_),
    .Y(\alu_out[30] ));
 sky130_fd_sc_hd__nor2_4 _34978_ (.A(_18742_),
    .B(_04557_),
    .Y(_04835_));
 sky130_fd_sc_hd__o21ai_4 _34979_ (.A1(_04741_),
    .A2(_04742_),
    .B1(_18742_),
    .Y(_04836_));
 sky130_fd_sc_hd__a21oi_4 _34980_ (.A1(_04836_),
    .A2(_04744_),
    .B1(_18744_),
    .Y(_04837_));
 sky130_fd_sc_hd__o21a_4 _34981_ (.A1(_04561_),
    .A2(_04563_),
    .B1(\alu_shl[31] ),
    .X(_04838_));
 sky130_fd_sc_hd__a2111oi_4 _34982_ (.A1(_04544_),
    .A2(\alu_shr[31] ),
    .B1(_04835_),
    .C1(_04837_),
    .D1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand3_4 _34983_ (.A(_04573_),
    .B(\alu_add_sub[31] ),
    .C(_04576_),
    .Y(_04840_));
 sky130_fd_sc_hd__o21ai_4 _34984_ (.A1(_04839_),
    .A2(_04570_),
    .B1(_04840_),
    .Y(\alu_out[31] ));
 sky130_fd_sc_hd__nor4_4 _34985_ (.A(_19068_),
    .B(_01786_),
    .C(_02530_),
    .D(_02818_),
    .Y(_04841_));
 sky130_vsdinv _34986_ (.A(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__buf_1 _34987_ (.A(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__buf_1 _34988_ (.A(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__nor3_4 _34989_ (.A(_02535_),
    .B(_02248_),
    .C(_02393_),
    .Y(_04845_));
 sky130_fd_sc_hd__a21o_4 _34990_ (.A1(\cpuregs[13][0] ),
    .A2(_04844_),
    .B1(_04845_),
    .X(_00865_));
 sky130_fd_sc_hd__and2_4 _34991_ (.A(_04841_),
    .B(_02253_),
    .X(_04846_));
 sky130_fd_sc_hd__a21o_4 _34992_ (.A1(\cpuregs[13][1] ),
    .A2(_04844_),
    .B1(_04846_),
    .X(_00876_));
 sky130_fd_sc_hd__buf_1 _34993_ (.A(_04842_),
    .X(_04847_));
 sky130_fd_sc_hd__buf_1 _34994_ (.A(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__nor2_4 _34995_ (.A(_04848_),
    .B(_02827_),
    .Y(_04849_));
 sky130_fd_sc_hd__a21o_4 _34996_ (.A1(\cpuregs[13][2] ),
    .A2(_04844_),
    .B1(_04849_),
    .X(_00887_));
 sky130_fd_sc_hd__nor2_4 _34997_ (.A(_04848_),
    .B(_03183_),
    .Y(_04850_));
 sky130_fd_sc_hd__a21o_4 _34998_ (.A1(\cpuregs[13][3] ),
    .A2(_04844_),
    .B1(_04850_),
    .X(_00890_));
 sky130_fd_sc_hd__buf_1 _34999_ (.A(_04843_),
    .X(_04851_));
 sky130_fd_sc_hd__a41oi_4 _35000_ (.A1(_02831_),
    .A2(_02832_),
    .A3(_02833_),
    .A4(_02834_),
    .B1(_04848_),
    .Y(_04852_));
 sky130_fd_sc_hd__a21o_4 _35001_ (.A1(\cpuregs[13][4] ),
    .A2(_04851_),
    .B1(_04852_),
    .X(_00891_));
 sky130_fd_sc_hd__a41oi_4 _35002_ (.A1(_02836_),
    .A2(_02837_),
    .A3(_02838_),
    .A4(_02839_),
    .B1(_04848_),
    .Y(_04853_));
 sky130_fd_sc_hd__a21o_4 _35003_ (.A1(\cpuregs[13][5] ),
    .A2(_04851_),
    .B1(_04853_),
    .X(_00892_));
 sky130_fd_sc_hd__buf_1 _35004_ (.A(_04842_),
    .X(_04854_));
 sky130_fd_sc_hd__buf_1 _35005_ (.A(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__a41oi_4 _35006_ (.A1(_02841_),
    .A2(_02842_),
    .A3(_02843_),
    .A4(_02844_),
    .B1(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__a21o_4 _35007_ (.A1(\cpuregs[13][6] ),
    .A2(_04851_),
    .B1(_04856_),
    .X(_00893_));
 sky130_fd_sc_hd__a41oi_4 _35008_ (.A1(_02848_),
    .A2(_02849_),
    .A3(_02850_),
    .A4(_02851_),
    .B1(_04855_),
    .Y(_04857_));
 sky130_fd_sc_hd__a21o_4 _35009_ (.A1(\cpuregs[13][7] ),
    .A2(_04851_),
    .B1(_04857_),
    .X(_00894_));
 sky130_fd_sc_hd__buf_1 _35010_ (.A(_04843_),
    .X(_04858_));
 sky130_fd_sc_hd__a41oi_4 _35011_ (.A1(_02854_),
    .A2(_02855_),
    .A3(_02856_),
    .A4(_02857_),
    .B1(_04855_),
    .Y(_04859_));
 sky130_fd_sc_hd__a21o_4 _35012_ (.A1(\cpuregs[13][8] ),
    .A2(_04858_),
    .B1(_04859_),
    .X(_00895_));
 sky130_fd_sc_hd__a41oi_4 _35013_ (.A1(_02859_),
    .A2(_02860_),
    .A3(_02861_),
    .A4(_02862_),
    .B1(_04855_),
    .Y(_04860_));
 sky130_fd_sc_hd__a21o_4 _35014_ (.A1(\cpuregs[13][9] ),
    .A2(_04858_),
    .B1(_04860_),
    .X(_00896_));
 sky130_fd_sc_hd__buf_1 _35015_ (.A(_04854_),
    .X(_04861_));
 sky130_fd_sc_hd__a41oi_4 _35016_ (.A1(_02864_),
    .A2(_02865_),
    .A3(_02866_),
    .A4(_02867_),
    .B1(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__a21o_4 _35017_ (.A1(\cpuregs[13][10] ),
    .A2(_04858_),
    .B1(_04862_),
    .X(_00866_));
 sky130_fd_sc_hd__a41oi_4 _35018_ (.A1(_02870_),
    .A2(_02871_),
    .A3(_02872_),
    .A4(_02873_),
    .B1(_04861_),
    .Y(_04863_));
 sky130_fd_sc_hd__a21o_4 _35019_ (.A1(\cpuregs[13][11] ),
    .A2(_04858_),
    .B1(_04863_),
    .X(_00867_));
 sky130_fd_sc_hd__buf_1 _35020_ (.A(_04842_),
    .X(_04864_));
 sky130_fd_sc_hd__buf_1 _35021_ (.A(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__a41oi_4 _35022_ (.A1(_02877_),
    .A2(_02878_),
    .A3(_02879_),
    .A4(_02880_),
    .B1(_04861_),
    .Y(_04866_));
 sky130_fd_sc_hd__a21o_4 _35023_ (.A1(\cpuregs[13][12] ),
    .A2(_04865_),
    .B1(_04866_),
    .X(_00868_));
 sky130_fd_sc_hd__a41oi_4 _35024_ (.A1(_02882_),
    .A2(_02883_),
    .A3(_02884_),
    .A4(_02885_),
    .B1(_04861_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21o_4 _35025_ (.A1(\cpuregs[13][13] ),
    .A2(_04865_),
    .B1(_04867_),
    .X(_00869_));
 sky130_fd_sc_hd__buf_1 _35026_ (.A(_04854_),
    .X(_04868_));
 sky130_fd_sc_hd__a41oi_4 _35027_ (.A1(_02887_),
    .A2(_02888_),
    .A3(_02889_),
    .A4(_02890_),
    .B1(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__a21o_4 _35028_ (.A1(\cpuregs[13][14] ),
    .A2(_04865_),
    .B1(_04869_),
    .X(_00870_));
 sky130_fd_sc_hd__a41oi_4 _35029_ (.A1(_02893_),
    .A2(_02894_),
    .A3(_02895_),
    .A4(_02896_),
    .B1(_04868_),
    .Y(_04870_));
 sky130_fd_sc_hd__a21o_4 _35030_ (.A1(\cpuregs[13][15] ),
    .A2(_04865_),
    .B1(_04870_),
    .X(_00871_));
 sky130_fd_sc_hd__buf_1 _35031_ (.A(_04864_),
    .X(_04871_));
 sky130_fd_sc_hd__a41oi_4 _35032_ (.A1(_02899_),
    .A2(_02900_),
    .A3(_02901_),
    .A4(_02902_),
    .B1(_04868_),
    .Y(_04872_));
 sky130_fd_sc_hd__a21o_4 _35033_ (.A1(\cpuregs[13][16] ),
    .A2(_04871_),
    .B1(_04872_),
    .X(_00872_));
 sky130_fd_sc_hd__a41oi_4 _35034_ (.A1(_02904_),
    .A2(_02905_),
    .A3(_02906_),
    .A4(_02907_),
    .B1(_04868_),
    .Y(_04873_));
 sky130_fd_sc_hd__a21o_4 _35035_ (.A1(\cpuregs[13][17] ),
    .A2(_04871_),
    .B1(_04873_),
    .X(_00873_));
 sky130_fd_sc_hd__buf_1 _35036_ (.A(_04847_),
    .X(_04874_));
 sky130_fd_sc_hd__a41oi_4 _35037_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_02911_),
    .A4(_02912_),
    .B1(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__a21o_4 _35038_ (.A1(\cpuregs[13][18] ),
    .A2(_04871_),
    .B1(_04875_),
    .X(_00874_));
 sky130_fd_sc_hd__a41oi_4 _35039_ (.A1(_02915_),
    .A2(_02916_),
    .A3(_02917_),
    .A4(_02918_),
    .B1(_04874_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21o_4 _35040_ (.A1(\cpuregs[13][19] ),
    .A2(_04871_),
    .B1(_04876_),
    .X(_00875_));
 sky130_fd_sc_hd__buf_1 _35041_ (.A(_04864_),
    .X(_04877_));
 sky130_fd_sc_hd__a41oi_4 _35042_ (.A1(_02921_),
    .A2(_02922_),
    .A3(_02923_),
    .A4(_02924_),
    .B1(_04874_),
    .Y(_04878_));
 sky130_fd_sc_hd__a21o_4 _35043_ (.A1(\cpuregs[13][20] ),
    .A2(_04877_),
    .B1(_04878_),
    .X(_00877_));
 sky130_fd_sc_hd__a41oi_4 _35044_ (.A1(_02926_),
    .A2(_02927_),
    .A3(_02928_),
    .A4(_02929_),
    .B1(_04874_),
    .Y(_04879_));
 sky130_fd_sc_hd__a21o_4 _35045_ (.A1(\cpuregs[13][21] ),
    .A2(_04877_),
    .B1(_04879_),
    .X(_00878_));
 sky130_fd_sc_hd__buf_1 _35046_ (.A(_04847_),
    .X(_04880_));
 sky130_fd_sc_hd__a41oi_4 _35047_ (.A1(_02931_),
    .A2(_02932_),
    .A3(_02933_),
    .A4(_02934_),
    .B1(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__a21o_4 _35048_ (.A1(\cpuregs[13][22] ),
    .A2(_04877_),
    .B1(_04881_),
    .X(_00879_));
 sky130_fd_sc_hd__a41oi_4 _35049_ (.A1(_02937_),
    .A2(_02938_),
    .A3(_02939_),
    .A4(_02940_),
    .B1(_04880_),
    .Y(_04882_));
 sky130_fd_sc_hd__a21o_4 _35050_ (.A1(\cpuregs[13][23] ),
    .A2(_04877_),
    .B1(_04882_),
    .X(_00880_));
 sky130_fd_sc_hd__buf_1 _35051_ (.A(_04864_),
    .X(_04883_));
 sky130_fd_sc_hd__a41oi_4 _35052_ (.A1(_02943_),
    .A2(_02944_),
    .A3(_02945_),
    .A4(_02946_),
    .B1(_04880_),
    .Y(_04884_));
 sky130_fd_sc_hd__a21o_4 _35053_ (.A1(\cpuregs[13][24] ),
    .A2(_04883_),
    .B1(_04884_),
    .X(_00881_));
 sky130_fd_sc_hd__a41oi_4 _35054_ (.A1(_02948_),
    .A2(_02949_),
    .A3(_02950_),
    .A4(_02951_),
    .B1(_04880_),
    .Y(_04885_));
 sky130_fd_sc_hd__a21o_4 _35055_ (.A1(\cpuregs[13][25] ),
    .A2(_04883_),
    .B1(_04885_),
    .X(_00882_));
 sky130_fd_sc_hd__buf_1 _35056_ (.A(_04847_),
    .X(_04886_));
 sky130_fd_sc_hd__a41oi_4 _35057_ (.A1(_02953_),
    .A2(_02954_),
    .A3(_02955_),
    .A4(_02956_),
    .B1(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__a21o_4 _35058_ (.A1(\cpuregs[13][26] ),
    .A2(_04883_),
    .B1(_04887_),
    .X(_00883_));
 sky130_fd_sc_hd__a41oi_4 _35059_ (.A1(_02959_),
    .A2(_02960_),
    .A3(_02961_),
    .A4(_02962_),
    .B1(_04886_),
    .Y(_04888_));
 sky130_fd_sc_hd__a21o_4 _35060_ (.A1(\cpuregs[13][27] ),
    .A2(_04883_),
    .B1(_04888_),
    .X(_00884_));
 sky130_fd_sc_hd__buf_1 _35061_ (.A(_04854_),
    .X(_04889_));
 sky130_fd_sc_hd__and2_4 _35062_ (.A(_02375_),
    .B(_04841_),
    .X(_04890_));
 sky130_fd_sc_hd__a21o_4 _35063_ (.A1(\cpuregs[13][28] ),
    .A2(_04889_),
    .B1(_04890_),
    .X(_00885_));
 sky130_fd_sc_hd__a41oi_4 _35064_ (.A1(_02966_),
    .A2(_02967_),
    .A3(_02968_),
    .A4(_02969_),
    .B1(_04886_),
    .Y(_04891_));
 sky130_fd_sc_hd__a21o_4 _35065_ (.A1(\cpuregs[13][29] ),
    .A2(_04889_),
    .B1(_04891_),
    .X(_00886_));
 sky130_fd_sc_hd__a41oi_4 _35066_ (.A1(_02971_),
    .A2(_02972_),
    .A3(_02973_),
    .A4(_02974_),
    .B1(_04886_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21o_4 _35067_ (.A1(\cpuregs[13][30] ),
    .A2(_04889_),
    .B1(_04892_),
    .X(_00888_));
 sky130_fd_sc_hd__a41oi_4 _35068_ (.A1(_02976_),
    .A2(_02977_),
    .A3(_02978_),
    .A4(_02979_),
    .B1(_04843_),
    .Y(_04893_));
 sky130_fd_sc_hd__a21o_4 _35069_ (.A1(\cpuregs[13][31] ),
    .A2(_04889_),
    .B1(_04893_),
    .X(_00889_));
 sky130_fd_sc_hd__nor2_4 _35070_ (.A(_02535_),
    .B(_02445_),
    .Y(_04894_));
 sky130_vsdinv _35071_ (.A(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__buf_1 _35072_ (.A(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__buf_1 _35073_ (.A(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__nor3_4 _35074_ (.A(_02450_),
    .B(_02535_),
    .C(_01783_),
    .Y(_04898_));
 sky130_fd_sc_hd__a21o_4 _35075_ (.A1(\cpuregs[12][0] ),
    .A2(_04897_),
    .B1(_04898_),
    .X(_00833_));
 sky130_fd_sc_hd__buf_1 _35076_ (.A(_04894_),
    .X(_04899_));
 sky130_fd_sc_hd__buf_1 _35077_ (.A(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__buf_1 _35078_ (.A(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__buf_1 _35079_ (.A(_04899_),
    .X(_04902_));
 sky130_fd_sc_hd__nand2_4 _35080_ (.A(_02989_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__o21ai_4 _35081_ (.A1(_19300_),
    .A2(_04901_),
    .B1(_04903_),
    .Y(_00844_));
 sky130_fd_sc_hd__buf_1 _35082_ (.A(_04896_),
    .X(_04904_));
 sky130_fd_sc_hd__a41oi_4 _35083_ (.A1(_02458_),
    .A2(_02460_),
    .A3(_02462_),
    .A4(_02464_),
    .B1(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21o_4 _35084_ (.A1(\cpuregs[12][2] ),
    .A2(_04897_),
    .B1(_04905_),
    .X(_00855_));
 sky130_fd_sc_hd__nor2_4 _35085_ (.A(_04897_),
    .B(_03183_),
    .Y(_04906_));
 sky130_fd_sc_hd__a21o_4 _35086_ (.A1(\cpuregs[12][3] ),
    .A2(_04897_),
    .B1(_04906_),
    .X(_00858_));
 sky130_fd_sc_hd__a41o_4 _35087_ (.A1(_01837_),
    .A2(_03112_),
    .A3(_01840_),
    .A4(_01843_),
    .B1(_04904_),
    .X(_04907_));
 sky130_fd_sc_hd__o21ai_4 _35088_ (.A1(_19579_),
    .A2(_04901_),
    .B1(_04907_),
    .Y(_00859_));
 sky130_fd_sc_hd__a41o_4 _35089_ (.A1(_01850_),
    .A2(_03117_),
    .A3(_01853_),
    .A4(_01857_),
    .B1(_04904_),
    .X(_04908_));
 sky130_fd_sc_hd__o21ai_4 _35090_ (.A1(_19658_),
    .A2(_04901_),
    .B1(_04908_),
    .Y(_00860_));
 sky130_fd_sc_hd__a41o_4 _35091_ (.A1(_01865_),
    .A2(_03119_),
    .A3(_01868_),
    .A4(_01871_),
    .B1(_04904_),
    .X(_04909_));
 sky130_fd_sc_hd__o21ai_4 _35092_ (.A1(_19703_),
    .A2(_04901_),
    .B1(_04909_),
    .Y(_00861_));
 sky130_fd_sc_hd__buf_1 _35093_ (.A(_04900_),
    .X(_04910_));
 sky130_fd_sc_hd__buf_1 _35094_ (.A(_04895_),
    .X(_04911_));
 sky130_fd_sc_hd__buf_1 _35095_ (.A(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__a41o_4 _35096_ (.A1(_01881_),
    .A2(_03121_),
    .A3(_01885_),
    .A4(_01888_),
    .B1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__o21ai_4 _35097_ (.A1(_19757_),
    .A2(_04910_),
    .B1(_04913_),
    .Y(_00862_));
 sky130_fd_sc_hd__a41o_4 _35098_ (.A1(_01895_),
    .A2(_03123_),
    .A3(_01898_),
    .A4(_01901_),
    .B1(_04912_),
    .X(_04914_));
 sky130_fd_sc_hd__o21ai_4 _35099_ (.A1(_19811_),
    .A2(_04910_),
    .B1(_04914_),
    .Y(_00863_));
 sky130_fd_sc_hd__a41o_4 _35100_ (.A1(_01908_),
    .A2(_03127_),
    .A3(_01911_),
    .A4(_01916_),
    .B1(_04912_),
    .X(_04915_));
 sky130_fd_sc_hd__o21ai_4 _35101_ (.A1(_19872_),
    .A2(_04910_),
    .B1(_04915_),
    .Y(_00864_));
 sky130_fd_sc_hd__a41o_4 _35102_ (.A1(_01923_),
    .A2(_03129_),
    .A3(_01926_),
    .A4(_01929_),
    .B1(_04912_),
    .X(_04916_));
 sky130_fd_sc_hd__o21ai_4 _35103_ (.A1(_19953_),
    .A2(_04910_),
    .B1(_04916_),
    .Y(_00834_));
 sky130_fd_sc_hd__buf_1 _35104_ (.A(_04900_),
    .X(_04917_));
 sky130_fd_sc_hd__buf_1 _35105_ (.A(_04911_),
    .X(_04918_));
 sky130_fd_sc_hd__a41o_4 _35106_ (.A1(_01938_),
    .A2(_03131_),
    .A3(_01942_),
    .A4(_01945_),
    .B1(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__o21ai_4 _35107_ (.A1(_19989_),
    .A2(_04917_),
    .B1(_04919_),
    .Y(_00835_));
 sky130_fd_sc_hd__a41o_4 _35108_ (.A1(_01953_),
    .A2(_03133_),
    .A3(_01956_),
    .A4(_01959_),
    .B1(_04918_),
    .X(_04920_));
 sky130_fd_sc_hd__o21ai_4 _35109_ (.A1(_20062_),
    .A2(_04917_),
    .B1(_04920_),
    .Y(_00836_));
 sky130_fd_sc_hd__a41o_4 _35110_ (.A1(_01967_),
    .A2(_03137_),
    .A3(_01970_),
    .A4(_01974_),
    .B1(_04918_),
    .X(_04921_));
 sky130_fd_sc_hd__o21ai_4 _35111_ (.A1(_20120_),
    .A2(_04917_),
    .B1(_04921_),
    .Y(_00837_));
 sky130_fd_sc_hd__a41o_4 _35112_ (.A1(_01983_),
    .A2(_03139_),
    .A3(_01986_),
    .A4(_01989_),
    .B1(_04918_),
    .X(_04922_));
 sky130_fd_sc_hd__o21ai_4 _35113_ (.A1(_20184_),
    .A2(_04917_),
    .B1(_04922_),
    .Y(_00838_));
 sky130_fd_sc_hd__buf_1 _35114_ (.A(_04899_),
    .X(_04923_));
 sky130_fd_sc_hd__buf_1 _35115_ (.A(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__buf_1 _35116_ (.A(_04911_),
    .X(_04925_));
 sky130_fd_sc_hd__a41o_4 _35117_ (.A1(_01999_),
    .A2(_03141_),
    .A3(_02003_),
    .A4(_02006_),
    .B1(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__o21ai_4 _35118_ (.A1(_20239_),
    .A2(_04924_),
    .B1(_04926_),
    .Y(_00839_));
 sky130_fd_sc_hd__a41o_4 _35119_ (.A1(_02016_),
    .A2(_03143_),
    .A3(_02019_),
    .A4(_02022_),
    .B1(_04925_),
    .X(_04927_));
 sky130_fd_sc_hd__o21ai_4 _35120_ (.A1(_20284_),
    .A2(_04924_),
    .B1(_04927_),
    .Y(_00840_));
 sky130_fd_sc_hd__a41o_4 _35121_ (.A1(_02031_),
    .A2(_03147_),
    .A3(_02034_),
    .A4(_02038_),
    .B1(_04925_),
    .X(_04928_));
 sky130_fd_sc_hd__o21ai_4 _35122_ (.A1(_20339_),
    .A2(_04924_),
    .B1(_04928_),
    .Y(_00841_));
 sky130_fd_sc_hd__nand2_4 _35123_ (.A(_03017_),
    .B(_04902_),
    .Y(_04929_));
 sky130_fd_sc_hd__o21ai_4 _35124_ (.A1(_20394_),
    .A2(_04924_),
    .B1(_04929_),
    .Y(_00842_));
 sky130_fd_sc_hd__buf_1 _35125_ (.A(_04923_),
    .X(_04930_));
 sky130_fd_sc_hd__a41o_4 _35126_ (.A1(_02061_),
    .A2(_03151_),
    .A3(_02064_),
    .A4(_02067_),
    .B1(_04925_),
    .X(_04931_));
 sky130_fd_sc_hd__o21ai_4 _35127_ (.A1(_20442_),
    .A2(_04930_),
    .B1(_04931_),
    .Y(_00843_));
 sky130_fd_sc_hd__buf_1 _35128_ (.A(_04911_),
    .X(_04932_));
 sky130_fd_sc_hd__a41o_4 _35129_ (.A1(_02077_),
    .A2(_03153_),
    .A3(_02081_),
    .A4(_02084_),
    .B1(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__o21ai_4 _35130_ (.A1(_20485_),
    .A2(_04930_),
    .B1(_04933_),
    .Y(_00845_));
 sky130_fd_sc_hd__a41o_4 _35131_ (.A1(_02092_),
    .A2(_03156_),
    .A3(_02095_),
    .A4(_02098_),
    .B1(_04932_),
    .X(_04934_));
 sky130_fd_sc_hd__o21ai_4 _35132_ (.A1(_20539_),
    .A2(_04930_),
    .B1(_04934_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_4 _35133_ (.A(_03024_),
    .B(_04902_),
    .Y(_04935_));
 sky130_fd_sc_hd__o21ai_4 _35134_ (.A1(_20595_),
    .A2(_04930_),
    .B1(_04935_),
    .Y(_00847_));
 sky130_fd_sc_hd__buf_1 _35135_ (.A(_04923_),
    .X(_04936_));
 sky130_fd_sc_hd__a41o_4 _35136_ (.A1(_02122_),
    .A2(_03160_),
    .A3(_02125_),
    .A4(_02129_),
    .B1(_04932_),
    .X(_04937_));
 sky130_fd_sc_hd__o21ai_4 _35137_ (.A1(_20622_),
    .A2(_04936_),
    .B1(_04937_),
    .Y(_00848_));
 sky130_fd_sc_hd__a41o_4 _35138_ (.A1(_02139_),
    .A2(_03162_),
    .A3(_02142_),
    .A4(_02145_),
    .B1(_04932_),
    .X(_04938_));
 sky130_fd_sc_hd__o21ai_4 _35139_ (.A1(_20667_),
    .A2(_04936_),
    .B1(_04938_),
    .Y(_00849_));
 sky130_fd_sc_hd__a41o_4 _35140_ (.A1(_02154_),
    .A2(_03165_),
    .A3(_02157_),
    .A4(_02160_),
    .B1(_04896_),
    .X(_04939_));
 sky130_fd_sc_hd__o21ai_4 _35141_ (.A1(_20715_),
    .A2(_04936_),
    .B1(_04939_),
    .Y(_00850_));
 sky130_fd_sc_hd__a41o_4 _35142_ (.A1(_02168_),
    .A2(_03167_),
    .A3(_02171_),
    .A4(_02174_),
    .B1(_04896_),
    .X(_04940_));
 sky130_fd_sc_hd__o21ai_4 _35143_ (.A1(_20758_),
    .A2(_04936_),
    .B1(_04940_),
    .Y(_00851_));
 sky130_fd_sc_hd__buf_1 _35144_ (.A(_04923_),
    .X(_04941_));
 sky130_fd_sc_hd__buf_1 _35145_ (.A(_04899_),
    .X(_04942_));
 sky130_fd_sc_hd__nand2_4 _35146_ (.A(_03032_),
    .B(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__o21ai_4 _35147_ (.A1(_20821_),
    .A2(_04941_),
    .B1(_04943_),
    .Y(_00852_));
 sky130_fd_sc_hd__nand2_4 _35148_ (.A(_03035_),
    .B(_04942_),
    .Y(_04944_));
 sky130_fd_sc_hd__o21ai_4 _35149_ (.A1(_20847_),
    .A2(_04941_),
    .B1(_04944_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_4 _35150_ (.A(_03037_),
    .B(_04942_),
    .Y(_04945_));
 sky130_fd_sc_hd__o21ai_4 _35151_ (.A1(_20896_),
    .A2(_04941_),
    .B1(_04945_),
    .Y(_00854_));
 sky130_fd_sc_hd__nand2_4 _35152_ (.A(_03039_),
    .B(_04942_),
    .Y(_04946_));
 sky130_fd_sc_hd__o21ai_4 _35153_ (.A1(_20936_),
    .A2(_04941_),
    .B1(_04946_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand2_4 _35154_ (.A(_03041_),
    .B(_04900_),
    .Y(_04947_));
 sky130_fd_sc_hd__o21ai_4 _35155_ (.A1(_20979_),
    .A2(_04902_),
    .B1(_04947_),
    .Y(_00857_));
 sky130_fd_sc_hd__and4_4 _35156_ (.A(_01784_),
    .B(_01785_),
    .C(_01786_),
    .D(_01764_),
    .X(_04948_));
 sky130_vsdinv _35157_ (.A(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__buf_1 _35158_ (.A(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__buf_1 _35159_ (.A(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__buf_1 _35160_ (.A(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__buf_1 _35161_ (.A(_04950_),
    .X(_04953_));
 sky130_fd_sc_hd__nor2_4 _35162_ (.A(_02451_),
    .B(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__a21o_4 _35163_ (.A1(\cpuregs[3][0] ),
    .A2(_04952_),
    .B1(_04954_),
    .X(_01153_));
 sky130_fd_sc_hd__and2_4 _35164_ (.A(_01803_),
    .B(_04948_),
    .X(_04955_));
 sky130_fd_sc_hd__a21o_4 _35165_ (.A1(\cpuregs[3][1] ),
    .A2(_04952_),
    .B1(_04955_),
    .X(_01164_));
 sky130_fd_sc_hd__a41oi_4 _35166_ (.A1(_02458_),
    .A2(_02460_),
    .A3(_02462_),
    .A4(_02464_),
    .B1(_04953_),
    .Y(_04956_));
 sky130_fd_sc_hd__a21o_4 _35167_ (.A1(\cpuregs[3][2] ),
    .A2(_04952_),
    .B1(_04956_),
    .X(_01175_));
 sky130_fd_sc_hd__a41oi_4 _35168_ (.A1(_23478_),
    .A2(_02263_),
    .A3(_02265_),
    .A4(_02267_),
    .B1(_04953_),
    .Y(_04957_));
 sky130_fd_sc_hd__a21o_4 _35169_ (.A1(\cpuregs[3][3] ),
    .A2(_04952_),
    .B1(_04957_),
    .X(_01178_));
 sky130_fd_sc_hd__buf_1 _35170_ (.A(_04951_),
    .X(_04958_));
 sky130_fd_sc_hd__a41oi_4 _35171_ (.A1(_23488_),
    .A2(_02269_),
    .A3(_02270_),
    .A4(_02271_),
    .B1(_04953_),
    .Y(_04959_));
 sky130_fd_sc_hd__a21o_4 _35172_ (.A1(\cpuregs[3][4] ),
    .A2(_04958_),
    .B1(_04959_),
    .X(_01179_));
 sky130_fd_sc_hd__buf_1 _35173_ (.A(_04949_),
    .X(_04960_));
 sky130_fd_sc_hd__buf_1 _35174_ (.A(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__a41oi_4 _35175_ (.A1(_23495_),
    .A2(_02276_),
    .A3(_02277_),
    .A4(_02278_),
    .B1(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__a21o_4 _35176_ (.A1(\cpuregs[3][5] ),
    .A2(_04958_),
    .B1(_04962_),
    .X(_01180_));
 sky130_fd_sc_hd__a41oi_4 _35177_ (.A1(_23505_),
    .A2(_02280_),
    .A3(_02281_),
    .A4(_02282_),
    .B1(_04961_),
    .Y(_04963_));
 sky130_fd_sc_hd__a21o_4 _35178_ (.A1(\cpuregs[3][6] ),
    .A2(_04958_),
    .B1(_04963_),
    .X(_01181_));
 sky130_fd_sc_hd__a41oi_4 _35179_ (.A1(_23511_),
    .A2(_02284_),
    .A3(_02285_),
    .A4(_02286_),
    .B1(_04961_),
    .Y(_04964_));
 sky130_fd_sc_hd__a21o_4 _35180_ (.A1(\cpuregs[3][7] ),
    .A2(_04958_),
    .B1(_04964_),
    .X(_01182_));
 sky130_fd_sc_hd__buf_1 _35181_ (.A(_04950_),
    .X(_04965_));
 sky130_fd_sc_hd__buf_1 _35182_ (.A(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__a41oi_4 _35183_ (.A1(_23520_),
    .A2(_02288_),
    .A3(_02289_),
    .A4(_02290_),
    .B1(_04961_),
    .Y(_04967_));
 sky130_fd_sc_hd__a21o_4 _35184_ (.A1(\cpuregs[3][8] ),
    .A2(_04966_),
    .B1(_04967_),
    .X(_01183_));
 sky130_fd_sc_hd__buf_1 _35185_ (.A(_04960_),
    .X(_04968_));
 sky130_fd_sc_hd__a41oi_4 _35186_ (.A1(_23527_),
    .A2(_02294_),
    .A3(_02295_),
    .A4(_02296_),
    .B1(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__a21o_4 _35187_ (.A1(\cpuregs[3][9] ),
    .A2(_04966_),
    .B1(_04969_),
    .X(_01184_));
 sky130_fd_sc_hd__a41oi_4 _35188_ (.A1(_23537_),
    .A2(_02298_),
    .A3(_02299_),
    .A4(_02300_),
    .B1(_04968_),
    .Y(_04970_));
 sky130_fd_sc_hd__a21o_4 _35189_ (.A1(\cpuregs[3][10] ),
    .A2(_04966_),
    .B1(_04970_),
    .X(_01154_));
 sky130_fd_sc_hd__a41oi_4 _35190_ (.A1(_23543_),
    .A2(_02302_),
    .A3(_02303_),
    .A4(_02304_),
    .B1(_04968_),
    .Y(_04971_));
 sky130_fd_sc_hd__a21o_4 _35191_ (.A1(\cpuregs[3][11] ),
    .A2(_04966_),
    .B1(_04971_),
    .X(_01155_));
 sky130_fd_sc_hd__buf_1 _35192_ (.A(_04965_),
    .X(_04972_));
 sky130_fd_sc_hd__a41oi_4 _35193_ (.A1(_23551_),
    .A2(_02306_),
    .A3(_02307_),
    .A4(_02308_),
    .B1(_04968_),
    .Y(_04973_));
 sky130_fd_sc_hd__a21o_4 _35194_ (.A1(\cpuregs[3][12] ),
    .A2(_04972_),
    .B1(_04973_),
    .X(_01156_));
 sky130_fd_sc_hd__buf_1 _35195_ (.A(_04950_),
    .X(_04974_));
 sky130_fd_sc_hd__buf_1 _35196_ (.A(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__a41oi_4 _35197_ (.A1(_23558_),
    .A2(_02312_),
    .A3(_02313_),
    .A4(_02314_),
    .B1(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__a21o_4 _35198_ (.A1(\cpuregs[3][13] ),
    .A2(_04972_),
    .B1(_04976_),
    .X(_01157_));
 sky130_fd_sc_hd__a41oi_4 _35199_ (.A1(_23568_),
    .A2(_02316_),
    .A3(_02317_),
    .A4(_02318_),
    .B1(_04975_),
    .Y(_04977_));
 sky130_fd_sc_hd__a21o_4 _35200_ (.A1(\cpuregs[3][14] ),
    .A2(_04972_),
    .B1(_04977_),
    .X(_01158_));
 sky130_fd_sc_hd__a41oi_4 _35201_ (.A1(_23574_),
    .A2(_02320_),
    .A3(_02321_),
    .A4(_02322_),
    .B1(_04975_),
    .Y(_04978_));
 sky130_fd_sc_hd__a21o_4 _35202_ (.A1(\cpuregs[3][15] ),
    .A2(_04972_),
    .B1(_04978_),
    .X(_01159_));
 sky130_fd_sc_hd__buf_1 _35203_ (.A(_04965_),
    .X(_04979_));
 sky130_fd_sc_hd__a41oi_4 _35204_ (.A1(_23583_),
    .A2(_02324_),
    .A3(_02325_),
    .A4(_02326_),
    .B1(_04975_),
    .Y(_04980_));
 sky130_fd_sc_hd__a21o_4 _35205_ (.A1(\cpuregs[3][16] ),
    .A2(_04979_),
    .B1(_04980_),
    .X(_01160_));
 sky130_fd_sc_hd__buf_1 _35206_ (.A(_04974_),
    .X(_04981_));
 sky130_fd_sc_hd__a41oi_4 _35207_ (.A1(_23591_),
    .A2(_02330_),
    .A3(_02331_),
    .A4(_02332_),
    .B1(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__a21o_4 _35208_ (.A1(\cpuregs[3][17] ),
    .A2(_04979_),
    .B1(_04982_),
    .X(_01161_));
 sky130_fd_sc_hd__a41oi_4 _35209_ (.A1(_23599_),
    .A2(_02044_),
    .A3(_02048_),
    .A4(_02051_),
    .B1(_04981_),
    .Y(_04983_));
 sky130_fd_sc_hd__a21o_4 _35210_ (.A1(\cpuregs[3][18] ),
    .A2(_04979_),
    .B1(_04983_),
    .X(_01162_));
 sky130_fd_sc_hd__a41oi_4 _35211_ (.A1(_23606_),
    .A2(_02338_),
    .A3(_02339_),
    .A4(_02340_),
    .B1(_04981_),
    .Y(_04984_));
 sky130_fd_sc_hd__a21o_4 _35212_ (.A1(\cpuregs[3][19] ),
    .A2(_04979_),
    .B1(_04984_),
    .X(_01163_));
 sky130_fd_sc_hd__buf_1 _35213_ (.A(_04965_),
    .X(_04985_));
 sky130_fd_sc_hd__a41oi_4 _35214_ (.A1(_23614_),
    .A2(_02342_),
    .A3(_02343_),
    .A4(_02344_),
    .B1(_04981_),
    .Y(_04986_));
 sky130_fd_sc_hd__a21o_4 _35215_ (.A1(\cpuregs[3][20] ),
    .A2(_04985_),
    .B1(_04986_),
    .X(_01165_));
 sky130_fd_sc_hd__buf_1 _35216_ (.A(_04974_),
    .X(_04987_));
 sky130_fd_sc_hd__a41oi_4 _35217_ (.A1(_23621_),
    .A2(_02347_),
    .A3(_02348_),
    .A4(_02349_),
    .B1(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__a21o_4 _35218_ (.A1(\cpuregs[3][21] ),
    .A2(_04985_),
    .B1(_04988_),
    .X(_01166_));
 sky130_fd_sc_hd__a41oi_4 _35219_ (.A1(_23628_),
    .A2(_02105_),
    .A3(_02108_),
    .A4(_02112_),
    .B1(_04987_),
    .Y(_04989_));
 sky130_fd_sc_hd__a21o_4 _35220_ (.A1(\cpuregs[3][22] ),
    .A2(_04985_),
    .B1(_04989_),
    .X(_01167_));
 sky130_fd_sc_hd__a41oi_4 _35221_ (.A1(_23634_),
    .A2(_02355_),
    .A3(_02356_),
    .A4(_02357_),
    .B1(_04987_),
    .Y(_04990_));
 sky130_fd_sc_hd__a21o_4 _35222_ (.A1(\cpuregs[3][23] ),
    .A2(_04985_),
    .B1(_04990_),
    .X(_01168_));
 sky130_fd_sc_hd__buf_1 _35223_ (.A(_04960_),
    .X(_04991_));
 sky130_fd_sc_hd__a41oi_4 _35224_ (.A1(_23642_),
    .A2(_02359_),
    .A3(_02360_),
    .A4(_02361_),
    .B1(_04987_),
    .Y(_04992_));
 sky130_fd_sc_hd__a21o_4 _35225_ (.A1(\cpuregs[3][24] ),
    .A2(_04991_),
    .B1(_04992_),
    .X(_01169_));
 sky130_fd_sc_hd__buf_1 _35226_ (.A(_04974_),
    .X(_04993_));
 sky130_fd_sc_hd__a41oi_4 _35227_ (.A1(_23649_),
    .A2(_02364_),
    .A3(_02365_),
    .A4(_02366_),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__a21o_4 _35228_ (.A1(\cpuregs[3][25] ),
    .A2(_04991_),
    .B1(_04994_),
    .X(_01170_));
 sky130_fd_sc_hd__a41oi_4 _35229_ (.A1(_23657_),
    .A2(_02368_),
    .A3(_02369_),
    .A4(_02370_),
    .B1(_04993_),
    .Y(_04995_));
 sky130_fd_sc_hd__a21o_4 _35230_ (.A1(\cpuregs[3][26] ),
    .A2(_04991_),
    .B1(_04995_),
    .X(_01171_));
 sky130_fd_sc_hd__a41oi_4 _35231_ (.A1(_23662_),
    .A2(_02183_),
    .A3(_02186_),
    .A4(_02189_),
    .B1(_04993_),
    .Y(_04996_));
 sky130_fd_sc_hd__a21o_4 _35232_ (.A1(\cpuregs[3][27] ),
    .A2(_04991_),
    .B1(_04996_),
    .X(_01172_));
 sky130_fd_sc_hd__buf_1 _35233_ (.A(_04960_),
    .X(_04997_));
 sky130_fd_sc_hd__and2_4 _35234_ (.A(_02375_),
    .B(_04948_),
    .X(_04998_));
 sky130_fd_sc_hd__a21o_4 _35235_ (.A1(\cpuregs[3][28] ),
    .A2(_04997_),
    .B1(_04998_),
    .X(_01173_));
 sky130_fd_sc_hd__a41oi_4 _35236_ (.A1(_23674_),
    .A2(_02205_),
    .A3(_02208_),
    .A4(_02211_),
    .B1(_04993_),
    .Y(_04999_));
 sky130_fd_sc_hd__a21o_4 _35237_ (.A1(\cpuregs[3][29] ),
    .A2(_04997_),
    .B1(_04999_),
    .X(_01174_));
 sky130_fd_sc_hd__a41oi_4 _35238_ (.A1(_23681_),
    .A2(_02218_),
    .A3(_02221_),
    .A4(_02224_),
    .B1(_04951_),
    .Y(_05000_));
 sky130_fd_sc_hd__a21o_4 _35239_ (.A1(\cpuregs[3][30] ),
    .A2(_04997_),
    .B1(_05000_),
    .X(_01176_));
 sky130_fd_sc_hd__a41oi_4 _35240_ (.A1(_23686_),
    .A2(_02232_),
    .A3(_02235_),
    .A4(_02238_),
    .B1(_04951_),
    .Y(_05001_));
 sky130_fd_sc_hd__a21o_4 _35241_ (.A1(\cpuregs[3][31] ),
    .A2(_04997_),
    .B1(_05001_),
    .X(_01177_));
 sky130_fd_sc_hd__and4_4 _35242_ (.A(_01763_),
    .B(_19068_),
    .C(_01786_),
    .D(_01764_),
    .X(_05002_));
 sky130_fd_sc_hd__buf_1 _35243_ (.A(_05002_),
    .X(_05003_));
 sky130_vsdinv _35244_ (.A(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__buf_1 _35245_ (.A(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__buf_1 _35246_ (.A(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__nor2_4 _35247_ (.A(_02451_),
    .B(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__a21o_4 _35248_ (.A1(\cpuregs[2][0] ),
    .A2(_05006_),
    .B1(_05007_),
    .X(_01121_));
 sky130_fd_sc_hd__buf_1 _35249_ (.A(_05003_),
    .X(_05008_));
 sky130_fd_sc_hd__buf_1 _35250_ (.A(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__buf_1 _35251_ (.A(_05003_),
    .X(_05010_));
 sky130_fd_sc_hd__buf_1 _35252_ (.A(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__nand2_4 _35253_ (.A(_02989_),
    .B(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__o21ai_4 _35254_ (.A1(_19347_),
    .A2(_05009_),
    .B1(_05012_),
    .Y(_01132_));
 sky130_fd_sc_hd__a41o_4 _35255_ (.A1(_02459_),
    .A2(_02597_),
    .A3(_02461_),
    .A4(_02463_),
    .B1(_05006_),
    .X(_05013_));
 sky130_fd_sc_hd__o21ai_4 _35256_ (.A1(_19467_),
    .A2(_05009_),
    .B1(_05013_),
    .Y(_01143_));
 sky130_fd_sc_hd__a41o_4 _35257_ (.A1(_02599_),
    .A2(_02262_),
    .A3(_02264_),
    .A4(_02266_),
    .B1(_05006_),
    .X(_05014_));
 sky130_fd_sc_hd__o21ai_4 _35258_ (.A1(_19546_),
    .A2(_05009_),
    .B1(_05014_),
    .Y(_01146_));
 sky130_fd_sc_hd__buf_1 _35259_ (.A(_05005_),
    .X(_05015_));
 sky130_fd_sc_hd__a41o_4 _35260_ (.A1(_01837_),
    .A2(_03112_),
    .A3(_01840_),
    .A4(_01843_),
    .B1(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__o21ai_4 _35261_ (.A1(_19611_),
    .A2(_05009_),
    .B1(_05016_),
    .Y(_01147_));
 sky130_fd_sc_hd__buf_1 _35262_ (.A(_05003_),
    .X(_05017_));
 sky130_fd_sc_hd__buf_1 _35263_ (.A(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__a41o_4 _35264_ (.A1(_01850_),
    .A2(_03117_),
    .A3(_01853_),
    .A4(_01857_),
    .B1(_05015_),
    .X(_05019_));
 sky130_fd_sc_hd__o21ai_4 _35265_ (.A1(_19674_),
    .A2(_05018_),
    .B1(_05019_),
    .Y(_01148_));
 sky130_fd_sc_hd__a41o_4 _35266_ (.A1(_01865_),
    .A2(_03119_),
    .A3(_01868_),
    .A4(_01871_),
    .B1(_05015_),
    .X(_05020_));
 sky130_fd_sc_hd__o21ai_4 _35267_ (.A1(_19724_),
    .A2(_05018_),
    .B1(_05020_),
    .Y(_01149_));
 sky130_fd_sc_hd__a41o_4 _35268_ (.A1(_01881_),
    .A2(_03121_),
    .A3(_01885_),
    .A4(_01888_),
    .B1(_05015_),
    .X(_05021_));
 sky130_fd_sc_hd__o21ai_4 _35269_ (.A1(_19774_),
    .A2(_05018_),
    .B1(_05021_),
    .Y(_01150_));
 sky130_fd_sc_hd__buf_1 _35270_ (.A(_05005_),
    .X(_05022_));
 sky130_fd_sc_hd__a41o_4 _35271_ (.A1(_01895_),
    .A2(_03123_),
    .A3(_01898_),
    .A4(_01901_),
    .B1(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__o21ai_4 _35272_ (.A1(_19834_),
    .A2(_05018_),
    .B1(_05023_),
    .Y(_01151_));
 sky130_fd_sc_hd__buf_1 _35273_ (.A(_05017_),
    .X(_05024_));
 sky130_fd_sc_hd__a41o_4 _35274_ (.A1(_01908_),
    .A2(_03127_),
    .A3(_01911_),
    .A4(_01916_),
    .B1(_05022_),
    .X(_05025_));
 sky130_fd_sc_hd__o21ai_4 _35275_ (.A1(_19894_),
    .A2(_05024_),
    .B1(_05025_),
    .Y(_01152_));
 sky130_fd_sc_hd__a41o_4 _35276_ (.A1(_01923_),
    .A2(_03129_),
    .A3(_01926_),
    .A4(_01929_),
    .B1(_05022_),
    .X(_05026_));
 sky130_fd_sc_hd__o21ai_4 _35277_ (.A1(_19937_),
    .A2(_05024_),
    .B1(_05026_),
    .Y(_01122_));
 sky130_fd_sc_hd__a41o_4 _35278_ (.A1(_01938_),
    .A2(_03131_),
    .A3(_01942_),
    .A4(_01945_),
    .B1(_05022_),
    .X(_05027_));
 sky130_fd_sc_hd__o21ai_4 _35279_ (.A1(_20011_),
    .A2(_05024_),
    .B1(_05027_),
    .Y(_01123_));
 sky130_fd_sc_hd__buf_1 _35280_ (.A(_05004_),
    .X(_05028_));
 sky130_fd_sc_hd__a41o_4 _35281_ (.A1(_01953_),
    .A2(_03133_),
    .A3(_01956_),
    .A4(_01959_),
    .B1(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__o21ai_4 _35282_ (.A1(_20088_),
    .A2(_05024_),
    .B1(_05029_),
    .Y(_01124_));
 sky130_fd_sc_hd__buf_1 _35283_ (.A(_05017_),
    .X(_05030_));
 sky130_fd_sc_hd__a41o_4 _35284_ (.A1(_01967_),
    .A2(_03137_),
    .A3(_01970_),
    .A4(_01974_),
    .B1(_05028_),
    .X(_05031_));
 sky130_fd_sc_hd__o21ai_4 _35285_ (.A1(_20139_),
    .A2(_05030_),
    .B1(_05031_),
    .Y(_01125_));
 sky130_fd_sc_hd__a41o_4 _35286_ (.A1(_01983_),
    .A2(_03139_),
    .A3(_01986_),
    .A4(_01989_),
    .B1(_05028_),
    .X(_05032_));
 sky130_fd_sc_hd__o21ai_4 _35287_ (.A1(_20205_),
    .A2(_05030_),
    .B1(_05032_),
    .Y(_01126_));
 sky130_fd_sc_hd__a41o_4 _35288_ (.A1(_01999_),
    .A2(_03141_),
    .A3(_02003_),
    .A4(_02006_),
    .B1(_05028_),
    .X(_05033_));
 sky130_fd_sc_hd__o21ai_4 _35289_ (.A1(_20254_),
    .A2(_05030_),
    .B1(_05033_),
    .Y(_01127_));
 sky130_fd_sc_hd__buf_1 _35290_ (.A(_05004_),
    .X(_05034_));
 sky130_fd_sc_hd__a41o_4 _35291_ (.A1(_02016_),
    .A2(_03143_),
    .A3(_02019_),
    .A4(_02022_),
    .B1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__o21ai_4 _35292_ (.A1(_20302_),
    .A2(_05030_),
    .B1(_05035_),
    .Y(_01128_));
 sky130_fd_sc_hd__buf_1 _35293_ (.A(_05017_),
    .X(_05036_));
 sky130_fd_sc_hd__a41o_4 _35294_ (.A1(_02031_),
    .A2(_03147_),
    .A3(_02034_),
    .A4(_02038_),
    .B1(_05034_),
    .X(_05037_));
 sky130_fd_sc_hd__o21ai_4 _35295_ (.A1(_20354_),
    .A2(_05036_),
    .B1(_05037_),
    .Y(_01129_));
 sky130_fd_sc_hd__buf_1 _35296_ (.A(_05010_),
    .X(_05038_));
 sky130_fd_sc_hd__nand2_4 _35297_ (.A(_03017_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__o21ai_4 _35298_ (.A1(_20409_),
    .A2(_05036_),
    .B1(_05039_),
    .Y(_01130_));
 sky130_fd_sc_hd__a41o_4 _35299_ (.A1(_02061_),
    .A2(_03151_),
    .A3(_02064_),
    .A4(_02067_),
    .B1(_05034_),
    .X(_05040_));
 sky130_fd_sc_hd__o21ai_4 _35300_ (.A1(_20459_),
    .A2(_05036_),
    .B1(_05040_),
    .Y(_01131_));
 sky130_fd_sc_hd__a41o_4 _35301_ (.A1(_02077_),
    .A2(_03153_),
    .A3(_02081_),
    .A4(_02084_),
    .B1(_05034_),
    .X(_05041_));
 sky130_fd_sc_hd__o21ai_4 _35302_ (.A1(_20503_),
    .A2(_05036_),
    .B1(_05041_),
    .Y(_01133_));
 sky130_fd_sc_hd__buf_1 _35303_ (.A(_05010_),
    .X(_05042_));
 sky130_fd_sc_hd__buf_1 _35304_ (.A(_05004_),
    .X(_05043_));
 sky130_fd_sc_hd__a41o_4 _35305_ (.A1(_02092_),
    .A2(_03156_),
    .A3(_02095_),
    .A4(_02098_),
    .B1(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__o21ai_4 _35306_ (.A1(_20554_),
    .A2(_05042_),
    .B1(_05044_),
    .Y(_01134_));
 sky130_fd_sc_hd__nand2_4 _35307_ (.A(_03024_),
    .B(_05038_),
    .Y(_05045_));
 sky130_fd_sc_hd__o21ai_4 _35308_ (.A1(_20580_),
    .A2(_05042_),
    .B1(_05045_),
    .Y(_01135_));
 sky130_fd_sc_hd__a41o_4 _35309_ (.A1(_02122_),
    .A2(_03160_),
    .A3(_02125_),
    .A4(_02129_),
    .B1(_05043_),
    .X(_05046_));
 sky130_fd_sc_hd__o21ai_4 _35310_ (.A1(_20637_),
    .A2(_05042_),
    .B1(_05046_),
    .Y(_01136_));
 sky130_fd_sc_hd__a41o_4 _35311_ (.A1(_02139_),
    .A2(_03162_),
    .A3(_02142_),
    .A4(_02145_),
    .B1(_05043_),
    .X(_05047_));
 sky130_fd_sc_hd__o21ai_4 _35312_ (.A1(_20683_),
    .A2(_05042_),
    .B1(_05047_),
    .Y(_01137_));
 sky130_fd_sc_hd__buf_1 _35313_ (.A(_05010_),
    .X(_05048_));
 sky130_fd_sc_hd__a41o_4 _35314_ (.A1(_02154_),
    .A2(_03165_),
    .A3(_02157_),
    .A4(_02160_),
    .B1(_05043_),
    .X(_05049_));
 sky130_fd_sc_hd__o21ai_4 _35315_ (.A1(_20730_),
    .A2(_05048_),
    .B1(_05049_),
    .Y(_01138_));
 sky130_fd_sc_hd__a41o_4 _35316_ (.A1(_02168_),
    .A2(_03167_),
    .A3(_02171_),
    .A4(_02174_),
    .B1(_05005_),
    .X(_05050_));
 sky130_fd_sc_hd__o21ai_4 _35317_ (.A1(_20773_),
    .A2(_05048_),
    .B1(_05050_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_4 _35318_ (.A(_03032_),
    .B(_05038_),
    .Y(_05051_));
 sky130_fd_sc_hd__o21ai_4 _35319_ (.A1(_20805_),
    .A2(_05048_),
    .B1(_05051_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand2_4 _35320_ (.A(_03035_),
    .B(_05038_),
    .Y(_05052_));
 sky130_fd_sc_hd__o21ai_4 _35321_ (.A1(_20862_),
    .A2(_05048_),
    .B1(_05052_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand2_4 _35322_ (.A(_03037_),
    .B(_05008_),
    .Y(_05053_));
 sky130_fd_sc_hd__o21ai_4 _35323_ (.A1(_20911_),
    .A2(_05011_),
    .B1(_05053_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand2_4 _35324_ (.A(_03039_),
    .B(_05008_),
    .Y(_05054_));
 sky130_fd_sc_hd__o21ai_4 _35325_ (.A1(_20951_),
    .A2(_05011_),
    .B1(_05054_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand2_4 _35326_ (.A(_03041_),
    .B(_05008_),
    .Y(_05055_));
 sky130_fd_sc_hd__o21ai_4 _35327_ (.A1(_20994_),
    .A2(_05011_),
    .B1(_05055_),
    .Y(_01145_));
 sky130_fd_sc_hd__and4_4 _35328_ (.A(_01784_),
    .B(_01785_),
    .C(_19086_),
    .D(_01764_),
    .X(_05056_));
 sky130_vsdinv _35329_ (.A(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__buf_1 _35330_ (.A(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__buf_1 _35331_ (.A(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__buf_1 _35332_ (.A(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__buf_1 _35333_ (.A(_05058_),
    .X(_05061_));
 sky130_fd_sc_hd__nor2_4 _35334_ (.A(_02451_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__a21o_4 _35335_ (.A1(\cpuregs[1][0] ),
    .A2(_05060_),
    .B1(_05062_),
    .X(_01089_));
 sky130_fd_sc_hd__and2_4 _35336_ (.A(_01803_),
    .B(_05056_),
    .X(_05063_));
 sky130_fd_sc_hd__a21o_4 _35337_ (.A1(\cpuregs[1][1] ),
    .A2(_05060_),
    .B1(_05063_),
    .X(_01100_));
 sky130_fd_sc_hd__a41oi_4 _35338_ (.A1(_23473_),
    .A2(_02258_),
    .A3(_02259_),
    .A4(_02260_),
    .B1(_05061_),
    .Y(_05064_));
 sky130_fd_sc_hd__a21o_4 _35339_ (.A1(\cpuregs[1][2] ),
    .A2(_05060_),
    .B1(_05064_),
    .X(_01111_));
 sky130_fd_sc_hd__a41oi_4 _35340_ (.A1(_23478_),
    .A2(_02263_),
    .A3(_02265_),
    .A4(_02267_),
    .B1(_05061_),
    .Y(_05065_));
 sky130_fd_sc_hd__a21o_4 _35341_ (.A1(\cpuregs[1][3] ),
    .A2(_05060_),
    .B1(_05065_),
    .X(_01114_));
 sky130_fd_sc_hd__buf_1 _35342_ (.A(_05059_),
    .X(_05066_));
 sky130_fd_sc_hd__a41oi_4 _35343_ (.A1(_23488_),
    .A2(_02269_),
    .A3(_02270_),
    .A4(_02271_),
    .B1(_05061_),
    .Y(_05067_));
 sky130_fd_sc_hd__a21o_4 _35344_ (.A1(\cpuregs[1][4] ),
    .A2(_05066_),
    .B1(_05067_),
    .X(_01115_));
 sky130_fd_sc_hd__buf_1 _35345_ (.A(_05057_),
    .X(_05068_));
 sky130_fd_sc_hd__buf_1 _35346_ (.A(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__a41oi_4 _35347_ (.A1(_23495_),
    .A2(_02276_),
    .A3(_02277_),
    .A4(_02278_),
    .B1(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__a21o_4 _35348_ (.A1(\cpuregs[1][5] ),
    .A2(_05066_),
    .B1(_05070_),
    .X(_01116_));
 sky130_fd_sc_hd__a41oi_4 _35349_ (.A1(_23505_),
    .A2(_02280_),
    .A3(_02281_),
    .A4(_02282_),
    .B1(_05069_),
    .Y(_05071_));
 sky130_fd_sc_hd__a21o_4 _35350_ (.A1(\cpuregs[1][6] ),
    .A2(_05066_),
    .B1(_05071_),
    .X(_01117_));
 sky130_fd_sc_hd__a41oi_4 _35351_ (.A1(_23511_),
    .A2(_02284_),
    .A3(_02285_),
    .A4(_02286_),
    .B1(_05069_),
    .Y(_05072_));
 sky130_fd_sc_hd__a21o_4 _35352_ (.A1(\cpuregs[1][7] ),
    .A2(_05066_),
    .B1(_05072_),
    .X(_01118_));
 sky130_fd_sc_hd__buf_1 _35353_ (.A(_05058_),
    .X(_05073_));
 sky130_fd_sc_hd__buf_1 _35354_ (.A(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__a41oi_4 _35355_ (.A1(_23520_),
    .A2(_02288_),
    .A3(_02289_),
    .A4(_02290_),
    .B1(_05069_),
    .Y(_05075_));
 sky130_fd_sc_hd__a21o_4 _35356_ (.A1(\cpuregs[1][8] ),
    .A2(_05074_),
    .B1(_05075_),
    .X(_01119_));
 sky130_fd_sc_hd__buf_1 _35357_ (.A(_05068_),
    .X(_05076_));
 sky130_fd_sc_hd__a41oi_4 _35358_ (.A1(_23527_),
    .A2(_02294_),
    .A3(_02295_),
    .A4(_02296_),
    .B1(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__a21o_4 _35359_ (.A1(\cpuregs[1][9] ),
    .A2(_05074_),
    .B1(_05077_),
    .X(_01120_));
 sky130_fd_sc_hd__a41oi_4 _35360_ (.A1(_23537_),
    .A2(_02298_),
    .A3(_02299_),
    .A4(_02300_),
    .B1(_05076_),
    .Y(_05078_));
 sky130_fd_sc_hd__a21o_4 _35361_ (.A1(\cpuregs[1][10] ),
    .A2(_05074_),
    .B1(_05078_),
    .X(_01090_));
 sky130_fd_sc_hd__a41oi_4 _35362_ (.A1(_23543_),
    .A2(_02302_),
    .A3(_02303_),
    .A4(_02304_),
    .B1(_05076_),
    .Y(_05079_));
 sky130_fd_sc_hd__a21o_4 _35363_ (.A1(\cpuregs[1][11] ),
    .A2(_05074_),
    .B1(_05079_),
    .X(_01091_));
 sky130_fd_sc_hd__buf_1 _35364_ (.A(_05073_),
    .X(_05080_));
 sky130_fd_sc_hd__a41oi_4 _35365_ (.A1(_23551_),
    .A2(_02306_),
    .A3(_02307_),
    .A4(_02308_),
    .B1(_05076_),
    .Y(_05081_));
 sky130_fd_sc_hd__a21o_4 _35366_ (.A1(\cpuregs[1][12] ),
    .A2(_05080_),
    .B1(_05081_),
    .X(_01092_));
 sky130_fd_sc_hd__buf_1 _35367_ (.A(_05058_),
    .X(_05082_));
 sky130_fd_sc_hd__buf_1 _35368_ (.A(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__a41oi_4 _35369_ (.A1(_23558_),
    .A2(_02312_),
    .A3(_02313_),
    .A4(_02314_),
    .B1(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__a21o_4 _35370_ (.A1(\cpuregs[1][13] ),
    .A2(_05080_),
    .B1(_05084_),
    .X(_01093_));
 sky130_fd_sc_hd__a41oi_4 _35371_ (.A1(_23568_),
    .A2(_02316_),
    .A3(_02317_),
    .A4(_02318_),
    .B1(_05083_),
    .Y(_05085_));
 sky130_fd_sc_hd__a21o_4 _35372_ (.A1(\cpuregs[1][14] ),
    .A2(_05080_),
    .B1(_05085_),
    .X(_01094_));
 sky130_fd_sc_hd__a41oi_4 _35373_ (.A1(_23574_),
    .A2(_02320_),
    .A3(_02321_),
    .A4(_02322_),
    .B1(_05083_),
    .Y(_05086_));
 sky130_fd_sc_hd__a21o_4 _35374_ (.A1(\cpuregs[1][15] ),
    .A2(_05080_),
    .B1(_05086_),
    .X(_01095_));
 sky130_fd_sc_hd__buf_1 _35375_ (.A(_05073_),
    .X(_05087_));
 sky130_fd_sc_hd__a41oi_4 _35376_ (.A1(_23583_),
    .A2(_02324_),
    .A3(_02325_),
    .A4(_02326_),
    .B1(_05083_),
    .Y(_05088_));
 sky130_fd_sc_hd__a21o_4 _35377_ (.A1(\cpuregs[1][16] ),
    .A2(_05087_),
    .B1(_05088_),
    .X(_01096_));
 sky130_fd_sc_hd__buf_1 _35378_ (.A(_05082_),
    .X(_05089_));
 sky130_fd_sc_hd__a41oi_4 _35379_ (.A1(_23591_),
    .A2(_02330_),
    .A3(_02331_),
    .A4(_02332_),
    .B1(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__a21o_4 _35380_ (.A1(\cpuregs[1][17] ),
    .A2(_05087_),
    .B1(_05090_),
    .X(_01097_));
 sky130_fd_sc_hd__a41oi_4 _35381_ (.A1(_23599_),
    .A2(_02044_),
    .A3(_02048_),
    .A4(_02051_),
    .B1(_05089_),
    .Y(_05091_));
 sky130_fd_sc_hd__a21o_4 _35382_ (.A1(\cpuregs[1][18] ),
    .A2(_05087_),
    .B1(_05091_),
    .X(_01098_));
 sky130_fd_sc_hd__a41oi_4 _35383_ (.A1(_23606_),
    .A2(_02338_),
    .A3(_02339_),
    .A4(_02340_),
    .B1(_05089_),
    .Y(_05092_));
 sky130_fd_sc_hd__a21o_4 _35384_ (.A1(\cpuregs[1][19] ),
    .A2(_05087_),
    .B1(_05092_),
    .X(_01099_));
 sky130_fd_sc_hd__buf_1 _35385_ (.A(_05073_),
    .X(_05093_));
 sky130_fd_sc_hd__a41oi_4 _35386_ (.A1(_23614_),
    .A2(_02342_),
    .A3(_02343_),
    .A4(_02344_),
    .B1(_05089_),
    .Y(_05094_));
 sky130_fd_sc_hd__a21o_4 _35387_ (.A1(\cpuregs[1][20] ),
    .A2(_05093_),
    .B1(_05094_),
    .X(_01101_));
 sky130_fd_sc_hd__buf_1 _35388_ (.A(_05082_),
    .X(_05095_));
 sky130_fd_sc_hd__a41oi_4 _35389_ (.A1(_23621_),
    .A2(_02347_),
    .A3(_02348_),
    .A4(_02349_),
    .B1(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__a21o_4 _35390_ (.A1(\cpuregs[1][21] ),
    .A2(_05093_),
    .B1(_05096_),
    .X(_01102_));
 sky130_fd_sc_hd__a41oi_4 _35391_ (.A1(_23628_),
    .A2(_02105_),
    .A3(_02108_),
    .A4(_02112_),
    .B1(_05095_),
    .Y(_05097_));
 sky130_fd_sc_hd__a21o_4 _35392_ (.A1(\cpuregs[1][22] ),
    .A2(_05093_),
    .B1(_05097_),
    .X(_01103_));
 sky130_fd_sc_hd__a41oi_4 _35393_ (.A1(_23634_),
    .A2(_02355_),
    .A3(_02356_),
    .A4(_02357_),
    .B1(_05095_),
    .Y(_05098_));
 sky130_fd_sc_hd__a21o_4 _35394_ (.A1(\cpuregs[1][23] ),
    .A2(_05093_),
    .B1(_05098_),
    .X(_01104_));
 sky130_fd_sc_hd__buf_1 _35395_ (.A(_05068_),
    .X(_05099_));
 sky130_fd_sc_hd__a41oi_4 _35396_ (.A1(_23642_),
    .A2(_02359_),
    .A3(_02360_),
    .A4(_02361_),
    .B1(_05095_),
    .Y(_05100_));
 sky130_fd_sc_hd__a21o_4 _35397_ (.A1(\cpuregs[1][24] ),
    .A2(_05099_),
    .B1(_05100_),
    .X(_01105_));
 sky130_fd_sc_hd__buf_1 _35398_ (.A(_05082_),
    .X(_05101_));
 sky130_fd_sc_hd__a41oi_4 _35399_ (.A1(_23649_),
    .A2(_02364_),
    .A3(_02365_),
    .A4(_02366_),
    .B1(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__a21o_4 _35400_ (.A1(\cpuregs[1][25] ),
    .A2(_05099_),
    .B1(_05102_),
    .X(_01106_));
 sky130_fd_sc_hd__a41oi_4 _35401_ (.A1(_23657_),
    .A2(_02368_),
    .A3(_02369_),
    .A4(_02370_),
    .B1(_05101_),
    .Y(_05103_));
 sky130_fd_sc_hd__a21o_4 _35402_ (.A1(\cpuregs[1][26] ),
    .A2(_05099_),
    .B1(_05103_),
    .X(_01107_));
 sky130_fd_sc_hd__a41oi_4 _35403_ (.A1(_23662_),
    .A2(_02183_),
    .A3(_02186_),
    .A4(_02189_),
    .B1(_05101_),
    .Y(_05104_));
 sky130_fd_sc_hd__a21o_4 _35404_ (.A1(\cpuregs[1][27] ),
    .A2(_05099_),
    .B1(_05104_),
    .X(_01108_));
 sky130_fd_sc_hd__buf_1 _35405_ (.A(_05068_),
    .X(_05105_));
 sky130_fd_sc_hd__and2_4 _35406_ (.A(_02375_),
    .B(_05056_),
    .X(_05106_));
 sky130_fd_sc_hd__a21o_4 _35407_ (.A1(\cpuregs[1][28] ),
    .A2(_05105_),
    .B1(_05106_),
    .X(_01109_));
 sky130_fd_sc_hd__a41oi_4 _35408_ (.A1(_23674_),
    .A2(_02205_),
    .A3(_02208_),
    .A4(_02211_),
    .B1(_05101_),
    .Y(_05107_));
 sky130_fd_sc_hd__a21o_4 _35409_ (.A1(\cpuregs[1][29] ),
    .A2(_05105_),
    .B1(_05107_),
    .X(_01110_));
 sky130_fd_sc_hd__a41oi_4 _35410_ (.A1(_23681_),
    .A2(_02218_),
    .A3(_02221_),
    .A4(_02224_),
    .B1(_05059_),
    .Y(_05108_));
 sky130_fd_sc_hd__a21o_4 _35411_ (.A1(\cpuregs[1][30] ),
    .A2(_05105_),
    .B1(_05108_),
    .X(_01112_));
 sky130_fd_sc_hd__a41oi_4 _35412_ (.A1(_23686_),
    .A2(_02232_),
    .A3(_02235_),
    .A4(_02238_),
    .B1(_05059_),
    .Y(_05109_));
 sky130_fd_sc_hd__a21o_4 _35413_ (.A1(\cpuregs[1][31] ),
    .A2(_05105_),
    .B1(_05109_),
    .X(_01113_));
 sky130_fd_sc_hd__buf_1 _35414_ (.A(\cpuregs[0][0] ),
    .X(_00737_));
 sky130_fd_sc_hd__buf_1 _35415_ (.A(\cpuregs[0][1] ),
    .X(_00748_));
 sky130_fd_sc_hd__buf_1 _35416_ (.A(\cpuregs[0][2] ),
    .X(_00759_));
 sky130_fd_sc_hd__buf_1 _35417_ (.A(\cpuregs[0][3] ),
    .X(_00762_));
 sky130_fd_sc_hd__buf_1 _35418_ (.A(\cpuregs[0][4] ),
    .X(_00763_));
 sky130_fd_sc_hd__buf_1 _35419_ (.A(\cpuregs[0][5] ),
    .X(_00764_));
 sky130_fd_sc_hd__buf_1 _35420_ (.A(\cpuregs[0][6] ),
    .X(_00765_));
 sky130_fd_sc_hd__buf_1 _35421_ (.A(\cpuregs[0][7] ),
    .X(_00766_));
 sky130_fd_sc_hd__buf_1 _35422_ (.A(\cpuregs[0][8] ),
    .X(_00767_));
 sky130_fd_sc_hd__buf_1 _35423_ (.A(\cpuregs[0][9] ),
    .X(_00768_));
 sky130_fd_sc_hd__buf_1 _35424_ (.A(\cpuregs[0][10] ),
    .X(_00738_));
 sky130_fd_sc_hd__buf_1 _35425_ (.A(\cpuregs[0][11] ),
    .X(_00739_));
 sky130_fd_sc_hd__buf_1 _35426_ (.A(\cpuregs[0][12] ),
    .X(_00740_));
 sky130_fd_sc_hd__buf_1 _35427_ (.A(\cpuregs[0][13] ),
    .X(_00741_));
 sky130_fd_sc_hd__buf_1 _35428_ (.A(\cpuregs[0][14] ),
    .X(_00742_));
 sky130_fd_sc_hd__buf_1 _35429_ (.A(\cpuregs[0][15] ),
    .X(_00743_));
 sky130_fd_sc_hd__buf_1 _35430_ (.A(\cpuregs[0][16] ),
    .X(_00744_));
 sky130_fd_sc_hd__buf_1 _35431_ (.A(\cpuregs[0][17] ),
    .X(_00745_));
 sky130_fd_sc_hd__buf_1 _35432_ (.A(\cpuregs[0][18] ),
    .X(_00746_));
 sky130_fd_sc_hd__buf_1 _35433_ (.A(\cpuregs[0][19] ),
    .X(_00747_));
 sky130_fd_sc_hd__buf_1 _35434_ (.A(\cpuregs[0][20] ),
    .X(_00749_));
 sky130_fd_sc_hd__buf_1 _35435_ (.A(\cpuregs[0][21] ),
    .X(_00750_));
 sky130_fd_sc_hd__buf_1 _35436_ (.A(\cpuregs[0][22] ),
    .X(_00751_));
 sky130_fd_sc_hd__buf_1 _35437_ (.A(\cpuregs[0][23] ),
    .X(_00752_));
 sky130_fd_sc_hd__buf_1 _35438_ (.A(\cpuregs[0][24] ),
    .X(_00753_));
 sky130_fd_sc_hd__buf_1 _35439_ (.A(\cpuregs[0][25] ),
    .X(_00754_));
 sky130_fd_sc_hd__buf_1 _35440_ (.A(\cpuregs[0][26] ),
    .X(_00755_));
 sky130_fd_sc_hd__buf_1 _35441_ (.A(\cpuregs[0][27] ),
    .X(_00756_));
 sky130_fd_sc_hd__buf_1 _35442_ (.A(\cpuregs[0][28] ),
    .X(_00757_));
 sky130_fd_sc_hd__buf_1 _35443_ (.A(\cpuregs[0][29] ),
    .X(_00758_));
 sky130_fd_sc_hd__buf_1 _35444_ (.A(\cpuregs[0][30] ),
    .X(_00760_));
 sky130_fd_sc_hd__buf_1 _35445_ (.A(\cpuregs[0][31] ),
    .X(_00761_));
 sky130_fd_sc_hd__buf_1 _35446_ (.A(\count_cycle[0] ),
    .X(_05110_));
 sky130_fd_sc_hd__nor2_4 _35447_ (.A(_05110_),
    .B(_19427_),
    .Y(_00004_));
 sky130_fd_sc_hd__or2_4 _35448_ (.A(_05110_),
    .B(_03723_),
    .X(_05111_));
 sky130_fd_sc_hd__buf_1 _35449_ (.A(_18861_),
    .X(_05112_));
 sky130_fd_sc_hd__nand2_4 _35450_ (.A(_05110_),
    .B(_03723_),
    .Y(_05113_));
 sky130_fd_sc_hd__and3_4 _35451_ (.A(_05111_),
    .B(_05112_),
    .C(_05113_),
    .X(_00015_));
 sky130_fd_sc_hd__nand2_4 _35452_ (.A(_05113_),
    .B(_03758_),
    .Y(_05114_));
 sky130_fd_sc_hd__nand3_4 _35453_ (.A(_05110_),
    .B(_03723_),
    .C(\count_cycle[2] ),
    .Y(_05115_));
 sky130_fd_sc_hd__and3_4 _35454_ (.A(_05114_),
    .B(_05112_),
    .C(_05115_),
    .X(_00026_));
 sky130_fd_sc_hd__a21oi_4 _35455_ (.A1(_05115_),
    .A2(_03786_),
    .B1(_18530_),
    .Y(_05116_));
 sky130_fd_sc_hd__nand4_4 _35456_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .D(\count_cycle[3] ),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_4 _35457_ (.A(_05116_),
    .B(_05117_),
    .Y(_05118_));
 sky130_vsdinv _35458_ (.A(_05118_),
    .Y(_00037_));
 sky130_fd_sc_hd__buf_1 _35459_ (.A(\count_cycle[4] ),
    .X(_05119_));
 sky130_vsdinv _35460_ (.A(_05117_),
    .Y(_05120_));
 sky130_fd_sc_hd__buf_1 _35461_ (.A(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__buf_1 _35462_ (.A(_18228_),
    .X(_05122_));
 sky130_fd_sc_hd__a21oi_4 _35463_ (.A1(_05121_),
    .A2(_05119_),
    .B1(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__o21a_4 _35464_ (.A1(_05119_),
    .A2(_05121_),
    .B1(_05123_),
    .X(_00048_));
 sky130_fd_sc_hd__a21oi_4 _35465_ (.A1(_05121_),
    .A2(_05119_),
    .B1(_03830_),
    .Y(_05124_));
 sky130_fd_sc_hd__and3_4 _35466_ (.A(_05120_),
    .B(\count_cycle[4] ),
    .C(_03830_),
    .X(_05125_));
 sky130_fd_sc_hd__or3_4 _35467_ (.A(_21022_),
    .B(_05124_),
    .C(_05125_),
    .X(_05126_));
 sky130_vsdinv _35468_ (.A(_05126_),
    .Y(_00059_));
 sky130_fd_sc_hd__a41oi_4 _35469_ (.A1(_05119_),
    .A2(_05121_),
    .A3(_03830_),
    .A4(\count_cycle[6] ),
    .B1(_23372_),
    .Y(_05127_));
 sky130_fd_sc_hd__o21a_4 _35470_ (.A1(\count_cycle[6] ),
    .A2(_05125_),
    .B1(_05127_),
    .X(_00064_));
 sky130_fd_sc_hd__buf_1 _35471_ (.A(\count_cycle[7] ),
    .X(_05128_));
 sky130_fd_sc_hd__and4_4 _35472_ (.A(_05120_),
    .B(\count_cycle[4] ),
    .C(\count_cycle[5] ),
    .D(\count_cycle[6] ),
    .X(_05129_));
 sky130_fd_sc_hd__buf_1 _35473_ (.A(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__o21ai_4 _35474_ (.A1(_05128_),
    .A2(_05130_),
    .B1(_23175_),
    .Y(_05131_));
 sky130_fd_sc_hd__a21o_4 _35475_ (.A1(_05128_),
    .A2(_05130_),
    .B1(_05131_),
    .X(_05132_));
 sky130_vsdinv _35476_ (.A(_05132_),
    .Y(_00065_));
 sky130_fd_sc_hd__a21oi_4 _35477_ (.A1(_05130_),
    .A2(_05128_),
    .B1(_03918_),
    .Y(_05133_));
 sky130_fd_sc_hd__and3_4 _35478_ (.A(_05129_),
    .B(\count_cycle[7] ),
    .C(_03918_),
    .X(_05134_));
 sky130_fd_sc_hd__nor3_4 _35479_ (.A(_18934_),
    .B(_05133_),
    .C(_05134_),
    .Y(_00066_));
 sky130_fd_sc_hd__a41oi_4 _35480_ (.A1(_05128_),
    .A2(_05130_),
    .A3(_03918_),
    .A4(_03957_),
    .B1(_23372_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21a_4 _35481_ (.A1(_03957_),
    .A2(_05134_),
    .B1(_05135_),
    .X(_00067_));
 sky130_fd_sc_hd__buf_1 _35482_ (.A(_03983_),
    .X(_05136_));
 sky130_fd_sc_hd__and4_4 _35483_ (.A(_05129_),
    .B(\count_cycle[7] ),
    .C(\count_cycle[8] ),
    .D(\count_cycle[9] ),
    .X(_05137_));
 sky130_fd_sc_hd__buf_1 _35484_ (.A(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__a21oi_4 _35485_ (.A1(_05138_),
    .A2(_05136_),
    .B1(_05122_),
    .Y(_05139_));
 sky130_fd_sc_hd__o21a_4 _35486_ (.A1(_05136_),
    .A2(_05138_),
    .B1(_05139_),
    .X(_00005_));
 sky130_fd_sc_hd__buf_1 _35487_ (.A(\count_cycle[11] ),
    .X(_05140_));
 sky130_fd_sc_hd__and2_4 _35488_ (.A(_05137_),
    .B(_03983_),
    .X(_05141_));
 sky130_fd_sc_hd__a41oi_4 _35489_ (.A1(_03957_),
    .A2(_05134_),
    .A3(_03983_),
    .A4(_05140_),
    .B1(_18285_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21ai_4 _35490_ (.A1(_05140_),
    .A2(_05141_),
    .B1(_05142_),
    .Y(_05143_));
 sky130_vsdinv _35491_ (.A(_05143_),
    .Y(_00006_));
 sky130_fd_sc_hd__and3_4 _35492_ (.A(_05138_),
    .B(_05136_),
    .C(_05140_),
    .X(_05144_));
 sky130_fd_sc_hd__a41oi_4 _35493_ (.A1(_05136_),
    .A2(_05138_),
    .A3(_05140_),
    .A4(\count_cycle[12] ),
    .B1(_23372_),
    .Y(_05145_));
 sky130_fd_sc_hd__o21a_4 _35494_ (.A1(\count_cycle[12] ),
    .A2(_05144_),
    .B1(_05145_),
    .X(_00007_));
 sky130_fd_sc_hd__buf_1 _35495_ (.A(\count_cycle[13] ),
    .X(_05146_));
 sky130_fd_sc_hd__and4_4 _35496_ (.A(_05137_),
    .B(\count_cycle[10] ),
    .C(\count_cycle[11] ),
    .D(\count_cycle[12] ),
    .X(_05147_));
 sky130_fd_sc_hd__buf_1 _35497_ (.A(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__a21oi_4 _35498_ (.A1(_05148_),
    .A2(_05146_),
    .B1(_05122_),
    .Y(_05149_));
 sky130_fd_sc_hd__o21a_4 _35499_ (.A1(_05146_),
    .A2(_05148_),
    .B1(_05149_),
    .X(_00008_));
 sky130_fd_sc_hd__a21oi_4 _35500_ (.A1(_05148_),
    .A2(_05146_),
    .B1(_04101_),
    .Y(_05150_));
 sky130_fd_sc_hd__and3_4 _35501_ (.A(_05147_),
    .B(\count_cycle[13] ),
    .C(_04101_),
    .X(_05151_));
 sky130_fd_sc_hd__buf_1 _35502_ (.A(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__nor3_4 _35503_ (.A(_18934_),
    .B(_05150_),
    .C(_05152_),
    .Y(_00009_));
 sky130_fd_sc_hd__buf_1 _35504_ (.A(\count_cycle[15] ),
    .X(_05153_));
 sky130_fd_sc_hd__buf_1 _35505_ (.A(_23371_),
    .X(_05154_));
 sky130_fd_sc_hd__a41oi_4 _35506_ (.A1(_05146_),
    .A2(_05148_),
    .A3(_04101_),
    .A4(_05153_),
    .B1(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21a_4 _35507_ (.A1(_05153_),
    .A2(_05152_),
    .B1(_05155_),
    .X(_00010_));
 sky130_fd_sc_hd__buf_1 _35508_ (.A(\count_cycle[16] ),
    .X(_05156_));
 sky130_fd_sc_hd__buf_1 _35509_ (.A(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__and4_4 _35510_ (.A(_05147_),
    .B(\count_cycle[13] ),
    .C(\count_cycle[14] ),
    .D(\count_cycle[15] ),
    .X(_05158_));
 sky130_fd_sc_hd__buf_1 _35511_ (.A(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__buf_1 _35512_ (.A(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__a21oi_4 _35513_ (.A1(_05160_),
    .A2(_05157_),
    .B1(_05122_),
    .Y(_05161_));
 sky130_fd_sc_hd__o21a_4 _35514_ (.A1(_05157_),
    .A2(_05160_),
    .B1(_05161_),
    .X(_00011_));
 sky130_fd_sc_hd__buf_1 _35515_ (.A(\count_cycle[17] ),
    .X(_05162_));
 sky130_fd_sc_hd__and2_4 _35516_ (.A(_05159_),
    .B(_05156_),
    .X(_05163_));
 sky130_fd_sc_hd__a41oi_4 _35517_ (.A1(\count_cycle[15] ),
    .A2(_05151_),
    .A3(_05156_),
    .A4(_05162_),
    .B1(_21056_),
    .Y(_05164_));
 sky130_fd_sc_hd__o21ai_4 _35518_ (.A1(_05162_),
    .A2(_05163_),
    .B1(_05164_),
    .Y(_05165_));
 sky130_vsdinv _35519_ (.A(_05165_),
    .Y(_00012_));
 sky130_fd_sc_hd__buf_1 _35520_ (.A(_05156_),
    .X(_05166_));
 sky130_fd_sc_hd__and3_4 _35521_ (.A(_05160_),
    .B(_05166_),
    .C(_05162_),
    .X(_05167_));
 sky130_fd_sc_hd__nand2_4 _35522_ (.A(_05162_),
    .B(\count_cycle[18] ),
    .Y(_05168_));
 sky130_vsdinv _35523_ (.A(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__a41oi_4 _35524_ (.A1(_05153_),
    .A2(_05152_),
    .A3(_05157_),
    .A4(_05169_),
    .B1(_05154_),
    .Y(_05170_));
 sky130_fd_sc_hd__o21a_4 _35525_ (.A1(\count_cycle[18] ),
    .A2(_05167_),
    .B1(_05170_),
    .X(_00013_));
 sky130_fd_sc_hd__and3_4 _35526_ (.A(_05159_),
    .B(_05166_),
    .C(_05169_),
    .X(_05171_));
 sky130_fd_sc_hd__nand3_4 _35527_ (.A(\count_cycle[17] ),
    .B(\count_cycle[18] ),
    .C(\count_cycle[19] ),
    .Y(_05172_));
 sky130_vsdinv _35528_ (.A(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__a41oi_4 _35529_ (.A1(_05153_),
    .A2(_05152_),
    .A3(_05166_),
    .A4(_05173_),
    .B1(_05154_),
    .Y(_05174_));
 sky130_fd_sc_hd__o21a_4 _35530_ (.A1(\count_cycle[19] ),
    .A2(_05171_),
    .B1(_05174_),
    .X(_00014_));
 sky130_fd_sc_hd__and3_4 _35531_ (.A(_05159_),
    .B(_05166_),
    .C(_05173_),
    .X(_05175_));
 sky130_fd_sc_hd__a41oi_4 _35532_ (.A1(_05157_),
    .A2(_05160_),
    .A3(\count_cycle[20] ),
    .A4(_05173_),
    .B1(_05154_),
    .Y(_05176_));
 sky130_fd_sc_hd__o21a_4 _35533_ (.A1(\count_cycle[20] ),
    .A2(_05175_),
    .B1(_05176_),
    .X(_00016_));
 sky130_fd_sc_hd__buf_1 _35534_ (.A(\count_cycle[21] ),
    .X(_05177_));
 sky130_fd_sc_hd__and4_4 _35535_ (.A(_05158_),
    .B(\count_cycle[16] ),
    .C(\count_cycle[20] ),
    .D(_05173_),
    .X(_05178_));
 sky130_fd_sc_hd__buf_1 _35536_ (.A(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__buf_1 _35537_ (.A(_24215_),
    .X(_05180_));
 sky130_fd_sc_hd__a21oi_4 _35538_ (.A1(_05179_),
    .A2(_05177_),
    .B1(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__o21a_4 _35539_ (.A1(_05177_),
    .A2(_05179_),
    .B1(_05181_),
    .X(_00017_));
 sky130_fd_sc_hd__buf_1 _35540_ (.A(_18783_),
    .X(_05182_));
 sky130_fd_sc_hd__a21oi_4 _35541_ (.A1(_05179_),
    .A2(_05177_),
    .B1(_04308_),
    .Y(_05183_));
 sky130_fd_sc_hd__and3_4 _35542_ (.A(_05178_),
    .B(\count_cycle[21] ),
    .C(_04308_),
    .X(_05184_));
 sky130_fd_sc_hd__nor3_4 _35543_ (.A(_05182_),
    .B(_05183_),
    .C(_05184_),
    .Y(_00018_));
 sky130_fd_sc_hd__buf_1 _35544_ (.A(_23371_),
    .X(_05185_));
 sky130_fd_sc_hd__a41oi_4 _35545_ (.A1(_05177_),
    .A2(_05179_),
    .A3(_04308_),
    .A4(_04333_),
    .B1(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__o21a_4 _35546_ (.A1(_04333_),
    .A2(_05184_),
    .B1(_05186_),
    .X(_00019_));
 sky130_fd_sc_hd__buf_1 _35547_ (.A(_04356_),
    .X(_05187_));
 sky130_fd_sc_hd__and4_4 _35548_ (.A(_05178_),
    .B(\count_cycle[21] ),
    .C(\count_cycle[22] ),
    .D(\count_cycle[23] ),
    .X(_05188_));
 sky130_fd_sc_hd__buf_1 _35549_ (.A(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__a21oi_4 _35550_ (.A1(_05189_),
    .A2(_05187_),
    .B1(_05180_),
    .Y(_05190_));
 sky130_fd_sc_hd__o21a_4 _35551_ (.A1(_05187_),
    .A2(_05189_),
    .B1(_05190_),
    .X(_00020_));
 sky130_fd_sc_hd__buf_1 _35552_ (.A(\count_cycle[25] ),
    .X(_05191_));
 sky130_fd_sc_hd__and2_4 _35553_ (.A(_05189_),
    .B(_04356_),
    .X(_05192_));
 sky130_fd_sc_hd__a41oi_4 _35554_ (.A1(_04333_),
    .A2(_05184_),
    .A3(_05187_),
    .A4(_05191_),
    .B1(_21056_),
    .Y(_05193_));
 sky130_fd_sc_hd__o21ai_4 _35555_ (.A1(_05191_),
    .A2(_05192_),
    .B1(_05193_),
    .Y(_05194_));
 sky130_vsdinv _35556_ (.A(_05194_),
    .Y(_00021_));
 sky130_fd_sc_hd__and3_4 _35557_ (.A(_05188_),
    .B(_04356_),
    .C(_05191_),
    .X(_05195_));
 sky130_fd_sc_hd__a41oi_4 _35558_ (.A1(_05187_),
    .A2(_05189_),
    .A3(_05191_),
    .A4(_04414_),
    .B1(_05185_),
    .Y(_05196_));
 sky130_fd_sc_hd__o21a_4 _35559_ (.A1(_04414_),
    .A2(_05195_),
    .B1(_05196_),
    .X(_00022_));
 sky130_fd_sc_hd__buf_1 _35560_ (.A(\count_cycle[27] ),
    .X(_05197_));
 sky130_fd_sc_hd__buf_1 _35561_ (.A(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__and4_4 _35562_ (.A(_05188_),
    .B(\count_cycle[24] ),
    .C(\count_cycle[25] ),
    .D(\count_cycle[26] ),
    .X(_05199_));
 sky130_fd_sc_hd__buf_1 _35563_ (.A(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__a21oi_4 _35564_ (.A1(_05200_),
    .A2(_05198_),
    .B1(_05180_),
    .Y(_05201_));
 sky130_fd_sc_hd__o21a_4 _35565_ (.A1(_05198_),
    .A2(_05200_),
    .B1(_05201_),
    .X(_00023_));
 sky130_fd_sc_hd__a21oi_4 _35566_ (.A1(_05200_),
    .A2(_05198_),
    .B1(\count_cycle[28] ),
    .Y(_05202_));
 sky130_fd_sc_hd__and3_4 _35567_ (.A(_05199_),
    .B(_05197_),
    .C(\count_cycle[28] ),
    .X(_05203_));
 sky130_fd_sc_hd__nor3_4 _35568_ (.A(_05182_),
    .B(_05202_),
    .C(_05203_),
    .Y(_00024_));
 sky130_fd_sc_hd__nand2_4 _35569_ (.A(\count_cycle[28] ),
    .B(\count_cycle[29] ),
    .Y(_05204_));
 sky130_vsdinv _35570_ (.A(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__a41oi_4 _35571_ (.A1(_04414_),
    .A2(_05195_),
    .A3(_05197_),
    .A4(_05205_),
    .B1(_05185_),
    .Y(_05206_));
 sky130_fd_sc_hd__o21a_4 _35572_ (.A1(\count_cycle[29] ),
    .A2(_05203_),
    .B1(_05206_),
    .X(_00025_));
 sky130_fd_sc_hd__buf_1 _35573_ (.A(\count_cycle[30] ),
    .X(_05207_));
 sky130_fd_sc_hd__and3_4 _35574_ (.A(_05199_),
    .B(_05197_),
    .C(_05205_),
    .X(_05208_));
 sky130_fd_sc_hd__a41oi_4 _35575_ (.A1(_05198_),
    .A2(_05200_),
    .A3(_05207_),
    .A4(_05205_),
    .B1(_05185_),
    .Y(_05209_));
 sky130_fd_sc_hd__o21a_4 _35576_ (.A1(_05207_),
    .A2(_05208_),
    .B1(_05209_),
    .X(_00027_));
 sky130_fd_sc_hd__buf_1 _35577_ (.A(_04523_),
    .X(_05210_));
 sky130_fd_sc_hd__buf_1 _35578_ (.A(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__and4_4 _35579_ (.A(_05199_),
    .B(\count_cycle[27] ),
    .C(\count_cycle[30] ),
    .D(_05205_),
    .X(_05212_));
 sky130_fd_sc_hd__buf_1 _35580_ (.A(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__buf_1 _35581_ (.A(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__buf_1 _35582_ (.A(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__a21oi_4 _35583_ (.A1(_05215_),
    .A2(_05211_),
    .B1(_05180_),
    .Y(_05216_));
 sky130_fd_sc_hd__o21a_4 _35584_ (.A1(_05211_),
    .A2(_05215_),
    .B1(_05216_),
    .X(_00028_));
 sky130_fd_sc_hd__a21o_4 _35585_ (.A1(_05214_),
    .A2(_05210_),
    .B1(_03693_),
    .X(_05217_));
 sky130_fd_sc_hd__nand3_4 _35586_ (.A(_05215_),
    .B(_03693_),
    .C(_05210_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand3_4 _35587_ (.A(_05217_),
    .B(_23097_),
    .C(_05218_),
    .Y(_05219_));
 sky130_vsdinv _35588_ (.A(_05219_),
    .Y(_00029_));
 sky130_fd_sc_hd__nand2_4 _35589_ (.A(_03693_),
    .B(\count_cycle[33] ),
    .Y(_05220_));
 sky130_vsdinv _35590_ (.A(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__a41o_4 _35591_ (.A1(_05208_),
    .A2(_05207_),
    .A3(_05210_),
    .A4(_05221_),
    .B1(_18530_),
    .X(_05222_));
 sky130_fd_sc_hd__a21oi_4 _35592_ (.A1(_03727_),
    .A2(_05218_),
    .B1(_05222_),
    .Y(_00030_));
 sky130_fd_sc_hd__buf_1 _35593_ (.A(_04523_),
    .X(_05223_));
 sky130_fd_sc_hd__and3_4 _35594_ (.A(_05213_),
    .B(_05223_),
    .C(_05221_),
    .X(_05224_));
 sky130_fd_sc_hd__o21a_4 _35595_ (.A1(\count_cycle[34] ),
    .A2(_05224_),
    .B1(_23410_),
    .X(_05225_));
 sky130_fd_sc_hd__and4_4 _35596_ (.A(_05214_),
    .B(\count_cycle[34] ),
    .C(_05223_),
    .D(_05221_),
    .X(_05226_));
 sky130_vsdinv _35597_ (.A(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__nand2_4 _35598_ (.A(_05225_),
    .B(_05227_),
    .Y(_05228_));
 sky130_vsdinv _35599_ (.A(_05228_),
    .Y(_00031_));
 sky130_fd_sc_hd__and4_4 _35600_ (.A(\count_cycle[32] ),
    .B(\count_cycle[33] ),
    .C(\count_cycle[34] ),
    .D(\count_cycle[35] ),
    .X(_05229_));
 sky130_fd_sc_hd__buf_1 _35601_ (.A(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__buf_1 _35602_ (.A(_23371_),
    .X(_05231_));
 sky130_fd_sc_hd__a41oi_4 _35603_ (.A1(_05207_),
    .A2(_05208_),
    .A3(_05211_),
    .A4(_05230_),
    .B1(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__o21a_4 _35604_ (.A1(\count_cycle[35] ),
    .A2(_05226_),
    .B1(_05232_),
    .X(_00032_));
 sky130_fd_sc_hd__and3_4 _35605_ (.A(_05213_),
    .B(_05223_),
    .C(_05230_),
    .X(_05233_));
 sky130_fd_sc_hd__o21a_4 _35606_ (.A1(\count_cycle[36] ),
    .A2(_05233_),
    .B1(_23410_),
    .X(_05234_));
 sky130_fd_sc_hd__and4_4 _35607_ (.A(_05214_),
    .B(\count_cycle[36] ),
    .C(_05223_),
    .D(_05230_),
    .X(_05235_));
 sky130_vsdinv _35608_ (.A(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_4 _35609_ (.A(_05234_),
    .B(_05236_),
    .Y(_05237_));
 sky130_vsdinv _35610_ (.A(_05237_),
    .Y(_00033_));
 sky130_fd_sc_hd__nand2_4 _35611_ (.A(\count_cycle[36] ),
    .B(\count_cycle[37] ),
    .Y(_05238_));
 sky130_vsdinv _35612_ (.A(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__a41oi_4 _35613_ (.A1(_05211_),
    .A2(_05215_),
    .A3(_05230_),
    .A4(_05239_),
    .B1(_05231_),
    .Y(_05240_));
 sky130_fd_sc_hd__o21a_4 _35614_ (.A1(\count_cycle[37] ),
    .A2(_05235_),
    .B1(_05240_),
    .X(_00034_));
 sky130_fd_sc_hd__and4_4 _35615_ (.A(_05212_),
    .B(\count_cycle[31] ),
    .C(_05229_),
    .D(_05239_),
    .X(_05241_));
 sky130_fd_sc_hd__and2_4 _35616_ (.A(_05241_),
    .B(_03863_),
    .X(_05242_));
 sky130_vsdinv _35617_ (.A(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__o21a_4 _35618_ (.A1(_03863_),
    .A2(_05241_),
    .B1(_23007_),
    .X(_05244_));
 sky130_fd_sc_hd__nand2_4 _35619_ (.A(_05243_),
    .B(_05244_),
    .Y(_05245_));
 sky130_vsdinv _35620_ (.A(_05245_),
    .Y(_00035_));
 sky130_fd_sc_hd__and2_4 _35621_ (.A(_05213_),
    .B(_04523_),
    .X(_05246_));
 sky130_fd_sc_hd__nand2_4 _35622_ (.A(\count_cycle[38] ),
    .B(\count_cycle[39] ),
    .Y(_05247_));
 sky130_vsdinv _35623_ (.A(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__nand4_4 _35624_ (.A(_05246_),
    .B(_05229_),
    .C(_05239_),
    .D(_05248_),
    .Y(_05249_));
 sky130_vsdinv _35625_ (.A(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__a21oi_4 _35626_ (.A1(_05241_),
    .A2(_03863_),
    .B1(\count_cycle[39] ),
    .Y(_05251_));
 sky130_fd_sc_hd__nor3_4 _35627_ (.A(_05182_),
    .B(_05250_),
    .C(_05251_),
    .Y(_00036_));
 sky130_vsdinv _35628_ (.A(\count_cycle[40] ),
    .Y(_05252_));
 sky130_fd_sc_hd__nor2_4 _35629_ (.A(_05252_),
    .B(_05249_),
    .Y(_05253_));
 sky130_vsdinv _35630_ (.A(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__a21oi_4 _35631_ (.A1(_05249_),
    .A2(_05252_),
    .B1(_18805_),
    .Y(_05255_));
 sky130_fd_sc_hd__nand2_4 _35632_ (.A(_05254_),
    .B(_05255_),
    .Y(_05256_));
 sky130_vsdinv _35633_ (.A(_05256_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_4 _35634_ (.A(\count_cycle[40] ),
    .B(\count_cycle[41] ),
    .Y(_05257_));
 sky130_vsdinv _35635_ (.A(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__a41oi_4 _35636_ (.A1(_05233_),
    .A2(_05239_),
    .A3(_05248_),
    .A4(_05258_),
    .B1(_05231_),
    .Y(_05259_));
 sky130_fd_sc_hd__o21a_4 _35637_ (.A1(\count_cycle[41] ),
    .A2(_05253_),
    .B1(_05259_),
    .X(_00039_));
 sky130_fd_sc_hd__nor2_4 _35638_ (.A(_05257_),
    .B(_05249_),
    .Y(_05260_));
 sky130_fd_sc_hd__buf_1 _35639_ (.A(_23262_),
    .X(_05261_));
 sky130_fd_sc_hd__o21a_4 _35640_ (.A1(_03986_),
    .A2(_05260_),
    .B1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__and4_4 _35641_ (.A(_05241_),
    .B(\count_cycle[42] ),
    .C(_05248_),
    .D(_05258_),
    .X(_05263_));
 sky130_fd_sc_hd__buf_1 _35642_ (.A(_05263_),
    .X(_05264_));
 sky130_vsdinv _35643_ (.A(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_4 _35644_ (.A(_05262_),
    .B(_05265_),
    .Y(_05266_));
 sky130_vsdinv _35645_ (.A(_05266_),
    .Y(_00040_));
 sky130_fd_sc_hd__buf_1 _35646_ (.A(_04024_),
    .X(_05267_));
 sky130_fd_sc_hd__a21oi_4 _35647_ (.A1(_05264_),
    .A2(_05267_),
    .B1(_18805_),
    .Y(_05268_));
 sky130_fd_sc_hd__o21ai_4 _35648_ (.A1(_05267_),
    .A2(_05264_),
    .B1(_05268_),
    .Y(_05269_));
 sky130_vsdinv _35649_ (.A(_05269_),
    .Y(_00041_));
 sky130_fd_sc_hd__and4_4 _35650_ (.A(_05250_),
    .B(\count_cycle[42] ),
    .C(\count_cycle[43] ),
    .D(_05258_),
    .X(_05270_));
 sky130_fd_sc_hd__o21a_4 _35651_ (.A1(\count_cycle[44] ),
    .A2(_05270_),
    .B1(_05261_),
    .X(_05271_));
 sky130_fd_sc_hd__and4_4 _35652_ (.A(_05260_),
    .B(_03986_),
    .C(_04024_),
    .D(\count_cycle[44] ),
    .X(_05272_));
 sky130_vsdinv _35653_ (.A(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__nand2_4 _35654_ (.A(_05271_),
    .B(_05273_),
    .Y(_05274_));
 sky130_vsdinv _35655_ (.A(_05274_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand2_4 _35656_ (.A(\count_cycle[44] ),
    .B(\count_cycle[45] ),
    .Y(_05275_));
 sky130_vsdinv _35657_ (.A(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__buf_1 _35658_ (.A(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__a41oi_4 _35659_ (.A1(_03986_),
    .A2(_05260_),
    .A3(_05267_),
    .A4(_05277_),
    .B1(_05231_),
    .Y(_05278_));
 sky130_fd_sc_hd__o21a_4 _35660_ (.A1(\count_cycle[45] ),
    .A2(_05272_),
    .B1(_05278_),
    .X(_00043_));
 sky130_fd_sc_hd__buf_1 _35661_ (.A(\count_cycle[46] ),
    .X(_05279_));
 sky130_fd_sc_hd__and4_4 _35662_ (.A(_05260_),
    .B(\count_cycle[42] ),
    .C(_04024_),
    .D(_05277_),
    .X(_05280_));
 sky130_fd_sc_hd__o21a_4 _35663_ (.A1(_05279_),
    .A2(_05280_),
    .B1(_05261_),
    .X(_05281_));
 sky130_fd_sc_hd__and4_4 _35664_ (.A(_05263_),
    .B(\count_cycle[43] ),
    .C(\count_cycle[46] ),
    .D(_05276_),
    .X(_05282_));
 sky130_vsdinv _35665_ (.A(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__nand2_4 _35666_ (.A(_05281_),
    .B(_05283_),
    .Y(_05284_));
 sky130_vsdinv _35667_ (.A(_05284_),
    .Y(_00044_));
 sky130_fd_sc_hd__buf_1 _35668_ (.A(_04128_),
    .X(_05285_));
 sky130_fd_sc_hd__a41oi_4 _35669_ (.A1(_05267_),
    .A2(_05264_),
    .A3(_05279_),
    .A4(_05277_),
    .B1(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__and4_4 _35670_ (.A(_05270_),
    .B(\count_cycle[46] ),
    .C(_04128_),
    .D(_05277_),
    .X(_05287_));
 sky130_fd_sc_hd__nor3_4 _35671_ (.A(_05182_),
    .B(_05286_),
    .C(_05287_),
    .Y(_00045_));
 sky130_fd_sc_hd__o21a_4 _35672_ (.A1(\count_cycle[48] ),
    .A2(_05287_),
    .B1(_05261_),
    .X(_05288_));
 sky130_fd_sc_hd__and4_4 _35673_ (.A(_05280_),
    .B(_05279_),
    .C(_05285_),
    .D(\count_cycle[48] ),
    .X(_05289_));
 sky130_vsdinv _35674_ (.A(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand2_4 _35675_ (.A(_05288_),
    .B(_05290_),
    .Y(_05291_));
 sky130_vsdinv _35676_ (.A(_05291_),
    .Y(_00046_));
 sky130_fd_sc_hd__nand2_4 _35677_ (.A(\count_cycle[48] ),
    .B(\count_cycle[49] ),
    .Y(_05292_));
 sky130_vsdinv _35678_ (.A(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__a41oi_4 _35679_ (.A1(_05279_),
    .A2(_05280_),
    .A3(_05285_),
    .A4(_05293_),
    .B1(_19131_),
    .Y(_05294_));
 sky130_fd_sc_hd__o21a_4 _35680_ (.A1(\count_cycle[49] ),
    .A2(_05289_),
    .B1(_05294_),
    .X(_00047_));
 sky130_fd_sc_hd__and4_4 _35681_ (.A(_05282_),
    .B(\count_cycle[47] ),
    .C(\count_cycle[50] ),
    .D(_05293_),
    .X(_05295_));
 sky130_vsdinv _35682_ (.A(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__nand3_4 _35683_ (.A(_05282_),
    .B(_04128_),
    .C(_05293_),
    .Y(_05297_));
 sky130_vsdinv _35684_ (.A(\count_cycle[50] ),
    .Y(_05298_));
 sky130_fd_sc_hd__a21oi_4 _35685_ (.A1(_05297_),
    .A2(_05298_),
    .B1(_18894_),
    .Y(_05299_));
 sky130_fd_sc_hd__nand2_4 _35686_ (.A(_05296_),
    .B(_05299_),
    .Y(_05300_));
 sky130_vsdinv _35687_ (.A(_05300_),
    .Y(_00049_));
 sky130_vsdinv _35688_ (.A(\count_cycle[51] ),
    .Y(_05301_));
 sky130_fd_sc_hd__nor3_4 _35689_ (.A(_05298_),
    .B(_05301_),
    .C(_05297_),
    .Y(_05302_));
 sky130_vsdinv _35690_ (.A(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__a41o_4 _35691_ (.A1(_05282_),
    .A2(_05285_),
    .A3(\count_cycle[50] ),
    .A4(_05293_),
    .B1(_04235_),
    .X(_05304_));
 sky130_fd_sc_hd__nand3_4 _35692_ (.A(_05303_),
    .B(_23739_),
    .C(_05304_),
    .Y(_05305_));
 sky130_vsdinv _35693_ (.A(_05305_),
    .Y(_00050_));
 sky130_fd_sc_hd__buf_1 _35694_ (.A(_23262_),
    .X(_05306_));
 sky130_fd_sc_hd__o21a_4 _35695_ (.A1(_04260_),
    .A2(_05302_),
    .B1(_05306_),
    .X(_05307_));
 sky130_vsdinv _35696_ (.A(\count_cycle[52] ),
    .Y(_05308_));
 sky130_fd_sc_hd__nor4_4 _35697_ (.A(_05298_),
    .B(_05301_),
    .C(_05308_),
    .D(_05297_),
    .Y(_05309_));
 sky130_vsdinv _35698_ (.A(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__nand2_4 _35699_ (.A(_05307_),
    .B(_05310_),
    .Y(_05311_));
 sky130_vsdinv _35700_ (.A(_05311_),
    .Y(_00051_));
 sky130_fd_sc_hd__a41oi_4 _35701_ (.A1(_04235_),
    .A2(_05295_),
    .A3(_04260_),
    .A4(_04287_),
    .B1(_19131_),
    .Y(_05312_));
 sky130_fd_sc_hd__o21a_4 _35702_ (.A1(_04287_),
    .A2(_05309_),
    .B1(_05312_),
    .X(_00052_));
 sky130_fd_sc_hd__and4_4 _35703_ (.A(_05295_),
    .B(_04235_),
    .C(\count_cycle[52] ),
    .D(\count_cycle[53] ),
    .X(_05313_));
 sky130_fd_sc_hd__o21a_4 _35704_ (.A1(_04311_),
    .A2(_05313_),
    .B1(_05306_),
    .X(_05314_));
 sky130_fd_sc_hd__and4_4 _35705_ (.A(_05302_),
    .B(_04260_),
    .C(\count_cycle[53] ),
    .D(\count_cycle[54] ),
    .X(_05315_));
 sky130_vsdinv _35706_ (.A(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_4 _35707_ (.A(_05314_),
    .B(_05316_),
    .Y(_05317_));
 sky130_vsdinv _35708_ (.A(_05317_),
    .Y(_00053_));
 sky130_fd_sc_hd__a41oi_4 _35709_ (.A1(_04287_),
    .A2(_05309_),
    .A3(_04311_),
    .A4(_04336_),
    .B1(_19131_),
    .Y(_05318_));
 sky130_fd_sc_hd__o21a_4 _35710_ (.A1(_04336_),
    .A2(_05315_),
    .B1(_05318_),
    .X(_00054_));
 sky130_fd_sc_hd__and4_4 _35711_ (.A(_05309_),
    .B(\count_cycle[53] ),
    .C(\count_cycle[54] ),
    .D(\count_cycle[55] ),
    .X(_05319_));
 sky130_fd_sc_hd__o21a_4 _35712_ (.A1(_04361_),
    .A2(_05319_),
    .B1(_05306_),
    .X(_05320_));
 sky130_fd_sc_hd__and4_4 _35713_ (.A(_05313_),
    .B(_04311_),
    .C(\count_cycle[55] ),
    .D(\count_cycle[56] ),
    .X(_05321_));
 sky130_vsdinv _35714_ (.A(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand2_4 _35715_ (.A(_05320_),
    .B(_05322_),
    .Y(_05323_));
 sky130_vsdinv _35716_ (.A(_05323_),
    .Y(_00055_));
 sky130_fd_sc_hd__a41oi_4 _35717_ (.A1(_04336_),
    .A2(_05315_),
    .A3(_04361_),
    .A4(_04387_),
    .B1(_21056_),
    .Y(_05324_));
 sky130_fd_sc_hd__o21ai_4 _35718_ (.A1(_04387_),
    .A2(_05321_),
    .B1(_05324_),
    .Y(_05325_));
 sky130_vsdinv _35719_ (.A(_05325_),
    .Y(_00056_));
 sky130_fd_sc_hd__and4_4 _35720_ (.A(_05315_),
    .B(\count_cycle[55] ),
    .C(\count_cycle[56] ),
    .D(\count_cycle[57] ),
    .X(_05326_));
 sky130_fd_sc_hd__o21a_4 _35721_ (.A1(_04417_),
    .A2(_05326_),
    .B1(_05306_),
    .X(_05327_));
 sky130_fd_sc_hd__nand4_4 _35722_ (.A(_04361_),
    .B(_05319_),
    .C(_04387_),
    .D(_04417_),
    .Y(_05328_));
 sky130_fd_sc_hd__nand2_4 _35723_ (.A(_05327_),
    .B(_05328_),
    .Y(_05329_));
 sky130_vsdinv _35724_ (.A(_05329_),
    .Y(_00057_));
 sky130_fd_sc_hd__buf_1 _35725_ (.A(\count_cycle[59] ),
    .X(_05330_));
 sky130_fd_sc_hd__and4_4 _35726_ (.A(_05319_),
    .B(\count_cycle[56] ),
    .C(\count_cycle[57] ),
    .D(\count_cycle[58] ),
    .X(_05331_));
 sky130_fd_sc_hd__buf_1 _35727_ (.A(_18548_),
    .X(_05332_));
 sky130_fd_sc_hd__o21a_4 _35728_ (.A1(_05330_),
    .A2(_05331_),
    .B1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__and4_4 _35729_ (.A(_05321_),
    .B(\count_cycle[57] ),
    .C(\count_cycle[58] ),
    .D(\count_cycle[59] ),
    .X(_05334_));
 sky130_vsdinv _35730_ (.A(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand2_4 _35731_ (.A(_05333_),
    .B(_05335_),
    .Y(_05336_));
 sky130_vsdinv _35732_ (.A(_05336_),
    .Y(_00058_));
 sky130_fd_sc_hd__buf_1 _35733_ (.A(\count_cycle[60] ),
    .X(_05337_));
 sky130_fd_sc_hd__o21a_4 _35734_ (.A1(_05337_),
    .A2(_05334_),
    .B1(_05332_),
    .X(_05338_));
 sky130_fd_sc_hd__and4_4 _35735_ (.A(_05326_),
    .B(_04417_),
    .C(_05330_),
    .D(\count_cycle[60] ),
    .X(_05339_));
 sky130_vsdinv _35736_ (.A(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__nand2_4 _35737_ (.A(_05338_),
    .B(_05340_),
    .Y(_05341_));
 sky130_vsdinv _35738_ (.A(_05341_),
    .Y(_00060_));
 sky130_fd_sc_hd__buf_1 _35739_ (.A(\count_cycle[61] ),
    .X(_05342_));
 sky130_fd_sc_hd__o21a_4 _35740_ (.A1(_05342_),
    .A2(_05339_),
    .B1(_05332_),
    .X(_05343_));
 sky130_fd_sc_hd__nand4_4 _35741_ (.A(_05330_),
    .B(_05331_),
    .C(_05337_),
    .D(_05342_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand2_4 _35742_ (.A(_05343_),
    .B(_05344_),
    .Y(_05345_));
 sky130_vsdinv _35743_ (.A(_05345_),
    .Y(_00061_));
 sky130_fd_sc_hd__buf_1 _35744_ (.A(\count_cycle[62] ),
    .X(_05346_));
 sky130_fd_sc_hd__and4_4 _35745_ (.A(_05331_),
    .B(_05330_),
    .C(\count_cycle[60] ),
    .D(\count_cycle[61] ),
    .X(_05347_));
 sky130_fd_sc_hd__o21a_4 _35746_ (.A1(_05346_),
    .A2(_05347_),
    .B1(_05332_),
    .X(_05348_));
 sky130_fd_sc_hd__nand4_4 _35747_ (.A(_05337_),
    .B(_05334_),
    .C(_05342_),
    .D(_05346_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_4 _35748_ (.A(_05348_),
    .B(_05349_),
    .Y(_05350_));
 sky130_vsdinv _35749_ (.A(_05350_),
    .Y(_00062_));
 sky130_fd_sc_hd__and4_4 _35750_ (.A(_05334_),
    .B(_05337_),
    .C(\count_cycle[61] ),
    .D(_05346_),
    .X(_05351_));
 sky130_fd_sc_hd__o21a_4 _35751_ (.A1(\count_cycle[63] ),
    .A2(_05351_),
    .B1(_23719_),
    .X(_05352_));
 sky130_fd_sc_hd__nand4_4 _35752_ (.A(_05342_),
    .B(_05339_),
    .C(_05346_),
    .D(\count_cycle[63] ),
    .Y(_05353_));
 sky130_fd_sc_hd__nand2_4 _35753_ (.A(_05352_),
    .B(_05353_),
    .Y(_05354_));
 sky130_vsdinv _35754_ (.A(_05354_),
    .Y(_00063_));
 sky130_fd_sc_hd__nor2_4 _35755_ (.A(_03049_),
    .B(_02444_),
    .Y(_05355_));
 sky130_vsdinv _35756_ (.A(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__buf_1 _35757_ (.A(_05356_),
    .X(_05357_));
 sky130_fd_sc_hd__buf_1 _35758_ (.A(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__nor3_4 _35759_ (.A(_02450_),
    .B(_03049_),
    .C(_01783_),
    .Y(_05359_));
 sky130_fd_sc_hd__a21o_4 _35760_ (.A1(\cpuregs[4][0] ),
    .A2(_05358_),
    .B1(_05359_),
    .X(_01185_));
 sky130_fd_sc_hd__buf_1 _35761_ (.A(_05355_),
    .X(_05360_));
 sky130_fd_sc_hd__buf_1 _35762_ (.A(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__buf_1 _35763_ (.A(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__buf_1 _35764_ (.A(_05360_),
    .X(_05363_));
 sky130_fd_sc_hd__nand2_4 _35765_ (.A(_01803_),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__o21ai_4 _35766_ (.A1(_19372_),
    .A2(_05362_),
    .B1(_05364_),
    .Y(_01196_));
 sky130_fd_sc_hd__buf_1 _35767_ (.A(_05357_),
    .X(_05365_));
 sky130_fd_sc_hd__a41oi_4 _35768_ (.A1(_23473_),
    .A2(_02258_),
    .A3(_02259_),
    .A4(_02260_),
    .B1(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__a21o_4 _35769_ (.A1(\cpuregs[4][2] ),
    .A2(_05358_),
    .B1(_05366_),
    .X(_01207_));
 sky130_fd_sc_hd__nor2_4 _35770_ (.A(_05358_),
    .B(_03183_),
    .Y(_05367_));
 sky130_fd_sc_hd__a21o_4 _35771_ (.A1(\cpuregs[4][3] ),
    .A2(_05358_),
    .B1(_05367_),
    .X(_01210_));
 sky130_fd_sc_hd__a41o_4 _35772_ (.A1(_01837_),
    .A2(_03112_),
    .A3(_01840_),
    .A4(_01843_),
    .B1(_05365_),
    .X(_05368_));
 sky130_fd_sc_hd__o21ai_4 _35773_ (.A1(_19622_),
    .A2(_05362_),
    .B1(_05368_),
    .Y(_01211_));
 sky130_fd_sc_hd__a41o_4 _35774_ (.A1(_01850_),
    .A2(_03117_),
    .A3(_01853_),
    .A4(_01857_),
    .B1(_05365_),
    .X(_05369_));
 sky130_fd_sc_hd__o21ai_4 _35775_ (.A1(_19682_),
    .A2(_05362_),
    .B1(_05369_),
    .Y(_01212_));
 sky130_fd_sc_hd__a41o_4 _35776_ (.A1(_01865_),
    .A2(_03119_),
    .A3(_01868_),
    .A4(_01871_),
    .B1(_05365_),
    .X(_05370_));
 sky130_fd_sc_hd__o21ai_4 _35777_ (.A1(_19734_),
    .A2(_05362_),
    .B1(_05370_),
    .Y(_01213_));
 sky130_fd_sc_hd__buf_1 _35778_ (.A(_05361_),
    .X(_05371_));
 sky130_fd_sc_hd__buf_1 _35779_ (.A(_05356_),
    .X(_05372_));
 sky130_fd_sc_hd__buf_1 _35780_ (.A(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__a41o_4 _35781_ (.A1(_01881_),
    .A2(_03121_),
    .A3(_01885_),
    .A4(_01888_),
    .B1(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__o21ai_4 _35782_ (.A1(_19781_),
    .A2(_05371_),
    .B1(_05374_),
    .Y(_01214_));
 sky130_fd_sc_hd__a41o_4 _35783_ (.A1(_01895_),
    .A2(_03123_),
    .A3(_01898_),
    .A4(_01901_),
    .B1(_05373_),
    .X(_05375_));
 sky130_fd_sc_hd__o21ai_4 _35784_ (.A1(_19847_),
    .A2(_05371_),
    .B1(_05375_),
    .Y(_01215_));
 sky130_fd_sc_hd__a41o_4 _35785_ (.A1(_01908_),
    .A2(_03127_),
    .A3(_01911_),
    .A4(_01916_),
    .B1(_05373_),
    .X(_05376_));
 sky130_fd_sc_hd__o21ai_4 _35786_ (.A1(_19903_),
    .A2(_05371_),
    .B1(_05376_),
    .Y(_01216_));
 sky130_fd_sc_hd__a41o_4 _35787_ (.A1(_01923_),
    .A2(_03129_),
    .A3(_01926_),
    .A4(_01929_),
    .B1(_05373_),
    .X(_05377_));
 sky130_fd_sc_hd__o21ai_4 _35788_ (.A1(_19945_),
    .A2(_05371_),
    .B1(_05377_),
    .Y(_01186_));
 sky130_fd_sc_hd__buf_1 _35789_ (.A(_05361_),
    .X(_05378_));
 sky130_fd_sc_hd__buf_1 _35790_ (.A(_05372_),
    .X(_05379_));
 sky130_fd_sc_hd__a41o_4 _35791_ (.A1(_01938_),
    .A2(_03131_),
    .A3(_01942_),
    .A4(_01945_),
    .B1(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__o21ai_4 _35792_ (.A1(_20023_),
    .A2(_05378_),
    .B1(_05380_),
    .Y(_01187_));
 sky130_fd_sc_hd__a41o_4 _35793_ (.A1(_01953_),
    .A2(_03133_),
    .A3(_01956_),
    .A4(_01959_),
    .B1(_05379_),
    .X(_05381_));
 sky130_fd_sc_hd__o21ai_4 _35794_ (.A1(_20097_),
    .A2(_05378_),
    .B1(_05381_),
    .Y(_01188_));
 sky130_fd_sc_hd__a41o_4 _35795_ (.A1(_01967_),
    .A2(_03137_),
    .A3(_01970_),
    .A4(_01974_),
    .B1(_05379_),
    .X(_05382_));
 sky130_fd_sc_hd__o21ai_4 _35796_ (.A1(_20149_),
    .A2(_05378_),
    .B1(_05382_),
    .Y(_01189_));
 sky130_fd_sc_hd__a41o_4 _35797_ (.A1(_01983_),
    .A2(_03139_),
    .A3(_01986_),
    .A4(_01989_),
    .B1(_05379_),
    .X(_05383_));
 sky130_fd_sc_hd__o21ai_4 _35798_ (.A1(_20214_),
    .A2(_05378_),
    .B1(_05383_),
    .Y(_01190_));
 sky130_fd_sc_hd__buf_1 _35799_ (.A(_05360_),
    .X(_05384_));
 sky130_fd_sc_hd__buf_1 _35800_ (.A(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__buf_1 _35801_ (.A(_05372_),
    .X(_05386_));
 sky130_fd_sc_hd__a41o_4 _35802_ (.A1(_01999_),
    .A2(_03141_),
    .A3(_02003_),
    .A4(_02006_),
    .B1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__o21ai_4 _35803_ (.A1(_20262_),
    .A2(_05385_),
    .B1(_05387_),
    .Y(_01191_));
 sky130_fd_sc_hd__a41o_4 _35804_ (.A1(_02016_),
    .A2(_03143_),
    .A3(_02019_),
    .A4(_02022_),
    .B1(_05386_),
    .X(_05388_));
 sky130_fd_sc_hd__o21ai_4 _35805_ (.A1(_20312_),
    .A2(_05385_),
    .B1(_05388_),
    .Y(_01192_));
 sky130_fd_sc_hd__a41o_4 _35806_ (.A1(_02031_),
    .A2(_03147_),
    .A3(_02034_),
    .A4(_02038_),
    .B1(_05386_),
    .X(_05389_));
 sky130_fd_sc_hd__o21ai_4 _35807_ (.A1(_20361_),
    .A2(_05385_),
    .B1(_05389_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_4 _35808_ (.A(_02334_),
    .B(_05363_),
    .Y(_05390_));
 sky130_fd_sc_hd__o21ai_4 _35809_ (.A1(_20416_),
    .A2(_05385_),
    .B1(_05390_),
    .Y(_01194_));
 sky130_fd_sc_hd__buf_1 _35810_ (.A(_05384_),
    .X(_05391_));
 sky130_fd_sc_hd__a41o_4 _35811_ (.A1(_02061_),
    .A2(_03151_),
    .A3(_02064_),
    .A4(_02067_),
    .B1(_05386_),
    .X(_05392_));
 sky130_fd_sc_hd__o21ai_4 _35812_ (.A1(_20466_),
    .A2(_05391_),
    .B1(_05392_),
    .Y(_01195_));
 sky130_fd_sc_hd__buf_1 _35813_ (.A(_05372_),
    .X(_05393_));
 sky130_fd_sc_hd__a41o_4 _35814_ (.A1(_02077_),
    .A2(_03153_),
    .A3(_02081_),
    .A4(_02084_),
    .B1(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__o21ai_4 _35815_ (.A1(_20510_),
    .A2(_05391_),
    .B1(_05394_),
    .Y(_01197_));
 sky130_fd_sc_hd__a41o_4 _35816_ (.A1(_02092_),
    .A2(_03156_),
    .A3(_02095_),
    .A4(_02098_),
    .B1(_05393_),
    .X(_05395_));
 sky130_fd_sc_hd__o21ai_4 _35817_ (.A1(_20561_),
    .A2(_05391_),
    .B1(_05395_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_4 _35818_ (.A(_02352_),
    .B(_05363_),
    .Y(_05396_));
 sky130_fd_sc_hd__o21ai_4 _35819_ (.A1(_20587_),
    .A2(_05391_),
    .B1(_05396_),
    .Y(_01199_));
 sky130_fd_sc_hd__buf_1 _35820_ (.A(_05384_),
    .X(_05397_));
 sky130_fd_sc_hd__a41o_4 _35821_ (.A1(_02122_),
    .A2(_03160_),
    .A3(_02125_),
    .A4(_02129_),
    .B1(_05393_),
    .X(_05398_));
 sky130_fd_sc_hd__o21ai_4 _35822_ (.A1(_20644_),
    .A2(_05397_),
    .B1(_05398_),
    .Y(_01200_));
 sky130_fd_sc_hd__a41o_4 _35823_ (.A1(_02139_),
    .A2(_03162_),
    .A3(_02142_),
    .A4(_02145_),
    .B1(_05393_),
    .X(_05399_));
 sky130_fd_sc_hd__o21ai_4 _35824_ (.A1(_20690_),
    .A2(_05397_),
    .B1(_05399_),
    .Y(_01201_));
 sky130_fd_sc_hd__a41o_4 _35825_ (.A1(_02154_),
    .A2(_03165_),
    .A3(_02157_),
    .A4(_02160_),
    .B1(_05357_),
    .X(_05400_));
 sky130_fd_sc_hd__o21ai_4 _35826_ (.A1(_20738_),
    .A2(_05397_),
    .B1(_05400_),
    .Y(_01202_));
 sky130_fd_sc_hd__a41o_4 _35827_ (.A1(_02168_),
    .A2(_03167_),
    .A3(_02171_),
    .A4(_02174_),
    .B1(_05357_),
    .X(_05401_));
 sky130_fd_sc_hd__o21ai_4 _35828_ (.A1(_20780_),
    .A2(_05397_),
    .B1(_05401_),
    .Y(_01203_));
 sky130_fd_sc_hd__buf_1 _35829_ (.A(_05384_),
    .X(_05402_));
 sky130_fd_sc_hd__buf_1 _35830_ (.A(_05360_),
    .X(_05403_));
 sky130_fd_sc_hd__nand2_4 _35831_ (.A(_02372_),
    .B(_05403_),
    .Y(_05404_));
 sky130_fd_sc_hd__o21ai_4 _35832_ (.A1(_20813_),
    .A2(_05402_),
    .B1(_05404_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_4 _35833_ (.A(_02198_),
    .B(_05403_),
    .Y(_05405_));
 sky130_fd_sc_hd__o21ai_4 _35834_ (.A1(_20869_),
    .A2(_05402_),
    .B1(_05405_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_4 _35835_ (.A(_02378_),
    .B(_05403_),
    .Y(_05406_));
 sky130_fd_sc_hd__o21ai_4 _35836_ (.A1(_20918_),
    .A2(_05402_),
    .B1(_05406_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_4 _35837_ (.A(_02381_),
    .B(_05403_),
    .Y(_05407_));
 sky130_fd_sc_hd__o21ai_4 _35838_ (.A1(_20958_),
    .A2(_05402_),
    .B1(_05407_),
    .Y(_01208_));
 sky130_fd_sc_hd__nand2_4 _35839_ (.A(_02384_),
    .B(_05361_),
    .Y(_05408_));
 sky130_fd_sc_hd__o21ai_4 _35840_ (.A1(_21001_),
    .A2(_05363_),
    .B1(_05408_),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_4 _35841_ (.A(_21991_),
    .B(irq[2]),
    .Y(_05409_));
 sky130_fd_sc_hd__and4_4 _35842_ (.A(_18956_),
    .B(_18959_),
    .C(_18416_),
    .D(_18936_),
    .X(_05410_));
 sky130_fd_sc_hd__o32ai_4 _35843_ (.A1(_18315_),
    .A2(_18531_),
    .A3(_18303_),
    .B1(_05409_),
    .B2(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__a21o_4 _35844_ (.A1(_05411_),
    .A2(_19112_),
    .B1(_18392_),
    .X(_00350_));
 sky130_vsdinv _35845_ (.A(pcpi_rs1[31]),
    .Y(_05412_));
 sky130_fd_sc_hd__buf_1 _35846_ (.A(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__buf_1 _35847_ (.A(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__nor2_4 _35848_ (.A(_21833_),
    .B(_21325_),
    .Y(_05415_));
 sky130_fd_sc_hd__maj3_4 _35849_ (.A(_21854_),
    .B(_05415_),
    .C(_01506_),
    .X(_05416_));
 sky130_fd_sc_hd__nor2_4 _35850_ (.A(_01689_),
    .B(_18760_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_4 _35851_ (.A(_18727_),
    .B(_18733_),
    .Y(_05418_));
 sky130_fd_sc_hd__maj3_4 _35852_ (.A(_18764_),
    .B(_05418_),
    .C(_21309_),
    .X(_05419_));
 sky130_fd_sc_hd__maj3_4 _35853_ (.A(_18724_),
    .B(_05419_),
    .C(_21315_),
    .X(_05420_));
 sky130_fd_sc_hd__a21oi_4 _35854_ (.A1(_18763_),
    .A2(_18761_),
    .B1(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__o21a_4 _35855_ (.A1(_05417_),
    .A2(_05421_),
    .B1(_18756_),
    .X(_05422_));
 sky130_fd_sc_hd__o21a_4 _35856_ (.A1(_05416_),
    .A2(_05422_),
    .B1(_18745_),
    .X(_05423_));
 sky130_fd_sc_hd__nor2_4 _35857_ (.A(_18744_),
    .B(_18743_),
    .Y(_05424_));
 sky130_fd_sc_hd__nor3_4 _35858_ (.A(_21871_),
    .B(_21334_),
    .C(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__nor2_4 _35859_ (.A(_18709_),
    .B(_21262_),
    .Y(_05426_));
 sky130_fd_sc_hd__maj3_4 _35860_ (.A(_21670_),
    .B(_05426_),
    .C(_18716_),
    .X(_05427_));
 sky130_fd_sc_hd__maj3_4 _35861_ (.A(_18701_),
    .B(_05427_),
    .C(_18706_),
    .X(_05428_));
 sky130_fd_sc_hd__maj3_4 _35862_ (.A(_21707_),
    .B(_05428_),
    .C(_18696_),
    .X(_05429_));
 sky130_fd_sc_hd__and2_4 _35863_ (.A(_05429_),
    .B(_18692_),
    .X(_05430_));
 sky130_fd_sc_hd__nor2_4 _35864_ (.A(_01671_),
    .B(_21300_),
    .Y(_05431_));
 sky130_fd_sc_hd__nor2_4 _35865_ (.A(_18666_),
    .B(_21284_),
    .Y(_05432_));
 sky130_fd_sc_hd__maj3_4 _35866_ (.A(_21740_),
    .B(_05432_),
    .C(_18682_),
    .X(_05433_));
 sky130_fd_sc_hd__maj3_4 _35867_ (.A(_21751_),
    .B(_05433_),
    .C(_18677_),
    .X(_05434_));
 sky130_fd_sc_hd__o21a_4 _35868_ (.A1(_18687_),
    .A2(_18690_),
    .B1(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__nor2_4 _35869_ (.A(_18660_),
    .B(_21204_),
    .Y(_05436_));
 sky130_fd_sc_hd__maj3_4 _35870_ (.A(_21528_),
    .B(_05436_),
    .C(pcpi_rs2[9]),
    .X(_05437_));
 sky130_fd_sc_hd__maj3_4 _35871_ (.A(_21546_),
    .B(_05437_),
    .C(_21227_),
    .X(_05438_));
 sky130_fd_sc_hd__maj3_4 _35872_ (.A(_21564_),
    .B(_05438_),
    .C(_18658_),
    .X(_05439_));
 sky130_fd_sc_hd__o21ai_4 _35873_ (.A1(_18628_),
    .A2(_21343_),
    .B1(_18621_),
    .Y(_05440_));
 sky130_fd_sc_hd__nor3_4 _35874_ (.A(_18628_),
    .B(_18621_),
    .C(_21343_),
    .Y(_05441_));
 sky130_vsdinv _35875_ (.A(_18618_),
    .Y(_05442_));
 sky130_fd_sc_hd__a211o_4 _35876_ (.A1(_18301_),
    .A2(_05440_),
    .B1(_05441_),
    .C1(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__nand2_4 _35877_ (.A(_21389_),
    .B(_03446_),
    .Y(_05444_));
 sky130_fd_sc_hd__maj3_4 _35878_ (.A(_21408_),
    .B(_05444_),
    .C(_21152_),
    .X(_05445_));
 sky130_fd_sc_hd__nand2_4 _35879_ (.A(_18593_),
    .B(_18606_),
    .Y(_05446_));
 sky130_fd_sc_hd__a21oi_4 _35880_ (.A1(_05443_),
    .A2(_05445_),
    .B1(_05446_),
    .Y(_05447_));
 sky130_fd_sc_hd__nor2_4 _35881_ (.A(_18600_),
    .B(_21166_),
    .Y(_05448_));
 sky130_fd_sc_hd__maj3_4 _35882_ (.A(_21455_),
    .B(_05448_),
    .C(_18583_),
    .X(_05449_));
 sky130_fd_sc_hd__maj3_4 _35883_ (.A(_21471_),
    .B(_05449_),
    .C(_18595_),
    .X(_05450_));
 sky130_fd_sc_hd__o21a_4 _35884_ (.A1(_18591_),
    .A2(_18592_),
    .B1(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__a211o_4 _35885_ (.A1(_21486_),
    .A2(_18589_),
    .B1(_05447_),
    .C1(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__and2_4 _35886_ (.A(_05452_),
    .B(_18663_),
    .X(_05453_));
 sky130_fd_sc_hd__o21ai_4 _35887_ (.A1(_05439_),
    .A2(_05453_),
    .B1(_18649_),
    .Y(_05454_));
 sky130_fd_sc_hd__nand3_4 _35888_ (.A(_18641_),
    .B(_21579_),
    .C(_18647_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21a_4 _35889_ (.A1(_21601_),
    .A2(_21244_),
    .B1(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__maj3_4 _35890_ (.A(_01630_),
    .B(_05456_),
    .C(_21250_),
    .X(_05457_));
 sky130_fd_sc_hd__maj3_4 _35891_ (.A(_01636_),
    .B(_05457_),
    .C(_21257_),
    .X(_05458_));
 sky130_fd_sc_hd__a21boi_4 _35892_ (.A1(_05454_),
    .A2(_05458_),
    .B1_N(_18719_),
    .Y(_05459_));
 sky130_fd_sc_hd__o41a_4 _35893_ (.A1(_05430_),
    .A2(_05431_),
    .A3(_05435_),
    .A4(_05459_),
    .B1(_18772_),
    .X(_05460_));
 sky130_fd_sc_hd__a2111o_4 _35894_ (.A1(_05414_),
    .A2(_21339_),
    .B1(_05423_),
    .C1(_05425_),
    .D1(_05460_),
    .X(_05461_));
 sky130_vsdinv _35895_ (.A(_00000_),
    .Y(_05462_));
 sky130_fd_sc_hd__o41ai_4 _35896_ (.A1(_05424_),
    .A2(_05423_),
    .A3(_05425_),
    .A4(_05460_),
    .B1(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__a21oi_4 _35897_ (.A1(_05461_),
    .A2(_05424_),
    .B1(_05463_),
    .Y(_00001_));
 sky130_fd_sc_hd__and2_4 _35898_ (.A(_05461_),
    .B(_05462_),
    .X(_00002_));
 sky130_fd_sc_hd__and3_4 _35899_ (.A(_19054_),
    .B(_05112_),
    .C(_19060_),
    .X(_00492_));
 sky130_fd_sc_hd__nor4_4 _35900_ (.A(_19082_),
    .B(_23104_),
    .C(_22101_),
    .D(_19084_),
    .Y(_00213_));
 sky130_fd_sc_hd__buf_1 _35901_ (.A(_23678_),
    .X(_05464_));
 sky130_fd_sc_hd__a21oi_4 _35902_ (.A1(_18856_),
    .A2(_18868_),
    .B1(_05464_),
    .Y(_00003_));
 sky130_fd_sc_hd__nand2_4 _35903_ (.A(_05112_),
    .B(\cpu_state[0] ),
    .Y(_05465_));
 sky130_vsdinv _35904_ (.A(_05465_),
    .Y(_00658_));
 sky130_fd_sc_hd__nor2_4 _35905_ (.A(_22996_),
    .B(_18838_),
    .Y(_05466_));
 sky130_fd_sc_hd__o21ai_4 _35906_ (.A1(_05466_),
    .A2(_21392_),
    .B1(latched_is_lb),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_4 _35907_ (.A(_21391_),
    .B(_03874_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand3_4 _35908_ (.A(_21371_),
    .B(instr_lb),
    .C(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__a21oi_4 _35909_ (.A1(_05467_),
    .A2(_05469_),
    .B1(_05464_),
    .Y(_00375_));
 sky130_fd_sc_hd__nand3_4 _35910_ (.A(_21371_),
    .B(_18837_),
    .C(_24126_),
    .Y(_05470_));
 sky130_fd_sc_hd__o21ai_4 _35911_ (.A1(_21391_),
    .A2(_18848_),
    .B1(_04131_),
    .Y(_05471_));
 sky130_fd_sc_hd__nand3_4 _35912_ (.A(_05470_),
    .B(_05471_),
    .C(_18365_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand3_4 _35913_ (.A(_19092_),
    .B(_03874_),
    .C(latched_is_lh),
    .Y(_05473_));
 sky130_fd_sc_hd__a21oi_4 _35914_ (.A1(_05472_),
    .A2(_05473_),
    .B1(_05464_),
    .Y(_00376_));
 sky130_fd_sc_hd__nor2_4 _35915_ (.A(_19142_),
    .B(_23865_),
    .Y(_05474_));
 sky130_fd_sc_hd__nor2_4 _35916_ (.A(_18864_),
    .B(_19046_),
    .Y(_05475_));
 sky130_fd_sc_hd__o21a_4 _35917_ (.A1(_05474_),
    .A2(_05475_),
    .B1(_18522_),
    .X(_05476_));
 sky130_fd_sc_hd__a211o_4 _35918_ (.A1(_18857_),
    .A2(_21908_),
    .B1(_04002_),
    .C1(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__nand3_4 _35919_ (.A(_23030_),
    .B(_21950_),
    .C(_23113_),
    .Y(_05478_));
 sky130_fd_sc_hd__nor2_4 _35920_ (.A(_19070_),
    .B(\cpu_state[4] ),
    .Y(_05479_));
 sky130_fd_sc_hd__o21ai_4 _35921_ (.A1(_21583_),
    .A2(_05479_),
    .B1(_22875_),
    .Y(_05480_));
 sky130_fd_sc_hd__a41oi_4 _35922_ (.A1(_23463_),
    .A2(_05477_),
    .A3(_05478_),
    .A4(_05480_),
    .B1(_18286_),
    .Y(_00373_));
 sky130_fd_sc_hd__o21ai_4 _35923_ (.A1(_18866_),
    .A2(_18579_),
    .B1(_22845_),
    .Y(_05481_));
 sky130_fd_sc_hd__a21oi_4 _35924_ (.A1(_05481_),
    .A2(_18523_),
    .B1(_05464_),
    .Y(_00382_));
 sky130_fd_sc_hd__a41oi_4 _35925_ (.A1(_22009_),
    .A2(_21998_),
    .A3(_22020_),
    .A4(_22031_),
    .B1(_18557_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand4_4 _35926_ (.A(_22996_),
    .B(_19104_),
    .C(_19106_),
    .D(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__nand2_4 _35927_ (.A(_05475_),
    .B(_18522_),
    .Y(_05484_));
 sky130_fd_sc_hd__a21oi_4 _35928_ (.A1(_01761_),
    .A2(_18857_),
    .B1(_19037_),
    .Y(_05485_));
 sky130_fd_sc_hd__nor3_4 _35929_ (.A(_22814_),
    .B(_18322_),
    .C(_18515_),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_4 _35930_ (.A1(_21278_),
    .A2(_05486_),
    .B1(_18362_),
    .Y(_05487_));
 sky130_fd_sc_hd__a21oi_4 _35931_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand3_4 _35932_ (.A(_05479_),
    .B(_21226_),
    .C(_18270_),
    .Y(_05489_));
 sky130_vsdinv _35933_ (.A(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__a21o_4 _35934_ (.A1(_05483_),
    .A2(_05488_),
    .B1(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__nand4_4 _35935_ (.A(_18490_),
    .B(_18532_),
    .C(_18503_),
    .D(_18496_),
    .Y(_05492_));
 sky130_fd_sc_hd__a21o_4 _35936_ (.A1(_05492_),
    .A2(_18855_),
    .B1(_05490_),
    .X(_05493_));
 sky130_fd_sc_hd__nand2_4 _35937_ (.A(_05493_),
    .B(_22814_),
    .Y(_05494_));
 sky130_fd_sc_hd__buf_1 _35938_ (.A(_23678_),
    .X(_05495_));
 sky130_fd_sc_hd__a21oi_4 _35939_ (.A1(_05491_),
    .A2(_05494_),
    .B1(_05495_),
    .Y(_00383_));
 sky130_fd_sc_hd__or3_4 _35940_ (.A(_19100_),
    .B(\cpu_state[0] ),
    .C(_18477_),
    .X(_05496_));
 sky130_fd_sc_hd__o32ai_4 _35941_ (.A1(_03643_),
    .A2(_05496_),
    .A3(_21390_),
    .B1(_18834_),
    .B2(_18395_),
    .Y(_00419_));
 sky130_fd_sc_hd__a2bb2o_4 _35942_ (.A1_N(_18837_),
    .A2_N(_18395_),
    .B1(_18279_),
    .B2(_05468_),
    .X(_00417_));
 sky130_fd_sc_hd__nand3_4 _35943_ (.A(_05479_),
    .B(_21226_),
    .C(_18253_),
    .Y(_05497_));
 sky130_vsdinv _35944_ (.A(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_4 _35945_ (.A1(_19078_),
    .A2(_22705_),
    .B1(_22083_),
    .Y(_05499_));
 sky130_fd_sc_hd__o21ai_4 _35946_ (.A1(_18564_),
    .A2(_05482_),
    .B1(_18576_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_4 _35947_ (.A(_05499_),
    .B(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hd__nand2_4 _35948_ (.A(_18361_),
    .B(_18521_),
    .Y(_05502_));
 sky130_fd_sc_hd__o21a_4 _35949_ (.A1(_23710_),
    .A2(_18521_),
    .B1(_18399_),
    .X(_05503_));
 sky130_fd_sc_hd__and2_4 _35950_ (.A(_05479_),
    .B(_21225_),
    .X(_05504_));
 sky130_fd_sc_hd__nor2_4 _35951_ (.A(_19048_),
    .B(_23837_),
    .Y(_05505_));
 sky130_fd_sc_hd__a21oi_4 _35952_ (.A1(_05492_),
    .A2(_05505_),
    .B1(_18788_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21a_4 _35953_ (.A1(_23710_),
    .A2(_18802_),
    .B1(_18798_),
    .X(_05507_));
 sky130_fd_sc_hd__a2111o_4 _35954_ (.A1(_05502_),
    .A2(_05503_),
    .B1(_05504_),
    .C1(_05506_),
    .D1(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__a21oi_4 _35955_ (.A1(_05501_),
    .A2(_19122_),
    .B1(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__nand2_4 _35956_ (.A(_18273_),
    .B(_21226_),
    .Y(_05510_));
 sky130_fd_sc_hd__or3_4 _35957_ (.A(_05496_),
    .B(_05510_),
    .C(_19047_),
    .X(_05511_));
 sky130_fd_sc_hd__o41ai_4 _35958_ (.A1(_21031_),
    .A2(_23709_),
    .A3(_05498_),
    .A4(_05509_),
    .B1(_05511_),
    .Y(_00418_));
 sky130_fd_sc_hd__nor2_4 _35959_ (.A(_19101_),
    .B(_23462_),
    .Y(_05512_));
 sky130_fd_sc_hd__a211o_4 _35960_ (.A1(_18409_),
    .A2(_19130_),
    .B1(_18285_),
    .C1(_05512_),
    .X(_05513_));
 sky130_vsdinv _35961_ (.A(_05513_),
    .Y(_00294_));
 sky130_fd_sc_hd__a41o_4 _35962_ (.A1(_21948_),
    .A2(_22996_),
    .A3(_23159_),
    .A4(_21954_),
    .B1(_18463_),
    .X(_05514_));
 sky130_fd_sc_hd__nand4_4 _35963_ (.A(_18408_),
    .B(_19075_),
    .C(_23031_),
    .D(_23070_),
    .Y(_05515_));
 sky130_fd_sc_hd__a21oi_4 _35964_ (.A1(_05514_),
    .A2(_05515_),
    .B1(_05495_),
    .Y(_00295_));
 sky130_fd_sc_hd__o21a_4 _35965_ (.A1(pcpi_valid),
    .A2(_18535_),
    .B1(_23719_),
    .X(_05516_));
 sky130_fd_sc_hd__o21ai_4 _35966_ (.A1(_18537_),
    .A2(_18792_),
    .B1(_18535_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_4 _35967_ (.A(_05516_),
    .B(_05517_),
    .Y(_05518_));
 sky130_vsdinv _35968_ (.A(_05518_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand3_4 _35969_ (.A(_23706_),
    .B(_23789_),
    .C(_24128_),
    .Y(_05519_));
 sky130_fd_sc_hd__buf_1 _35970_ (.A(_24008_),
    .X(_05520_));
 sky130_fd_sc_hd__nand2_4 _35971_ (.A(_23691_),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__a21oi_4 _35972_ (.A1(_05519_),
    .A2(_05521_),
    .B1(_05495_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand3_4 _35973_ (.A(_18332_),
    .B(_18325_),
    .C(_18864_),
    .Y(_05522_));
 sky130_fd_sc_hd__and3_4 _35974_ (.A(_05522_),
    .B(_24000_),
    .C(_20932_),
    .X(_00365_));
 sky130_fd_sc_hd__buf_1 _35975_ (.A(_24078_),
    .X(_05523_));
 sky130_fd_sc_hd__buf_1 _35976_ (.A(_22708_),
    .X(_05524_));
 sky130_fd_sc_hd__o21a_4 _35977_ (.A1(_05523_),
    .A2(_05524_),
    .B1(instr_and),
    .X(_05525_));
 sky130_fd_sc_hd__nand3_4 _35978_ (.A(_24123_),
    .B(_23807_),
    .C(_24104_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand3_4 _35979_ (.A(_24058_),
    .B(_23784_),
    .C(_24102_),
    .Y(_05527_));
 sky130_fd_sc_hd__nor2_4 _35980_ (.A(_05526_),
    .B(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__o21a_4 _35981_ (.A1(_05525_),
    .A2(_05528_),
    .B1(_23379_),
    .X(_00248_));
 sky130_fd_sc_hd__o21a_4 _35982_ (.A1(_05523_),
    .A2(_05524_),
    .B1(instr_or),
    .X(_05529_));
 sky130_fd_sc_hd__nand3_4 _35983_ (.A(_23808_),
    .B(_23807_),
    .C(_24104_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_4 _35984_ (.A(_05530_),
    .B(_05527_),
    .Y(_05531_));
 sky130_fd_sc_hd__o21a_4 _35985_ (.A1(_05529_),
    .A2(_05531_),
    .B1(_23379_),
    .X(_00268_));
 sky130_fd_sc_hd__and4_4 _35986_ (.A(_18875_),
    .B(_23900_),
    .C(_24104_),
    .D(is_alu_reg_reg),
    .X(_05532_));
 sky130_fd_sc_hd__nand3_4 _35987_ (.A(_23822_),
    .B(_24170_),
    .C(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__buf_1 _35988_ (.A(_24053_),
    .X(_05534_));
 sky130_fd_sc_hd__buf_1 _35989_ (.A(_24054_),
    .X(_05535_));
 sky130_fd_sc_hd__o21ai_4 _35990_ (.A1(_05534_),
    .A2(_05535_),
    .B1(instr_sra),
    .Y(_05536_));
 sky130_fd_sc_hd__a21oi_4 _35991_ (.A1(_05533_),
    .A2(_05536_),
    .B1(_05495_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand3_4 _35992_ (.A(_24059_),
    .B(_24170_),
    .C(_05532_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_4 _35993_ (.A1(_05534_),
    .A2(_05535_),
    .B1(instr_srl),
    .Y(_05538_));
 sky130_fd_sc_hd__buf_1 _35994_ (.A(_23678_),
    .X(_05539_));
 sky130_fd_sc_hd__a21oi_4 _35995_ (.A1(_05537_),
    .A2(_05538_),
    .B1(_05539_),
    .Y(_00286_));
 sky130_fd_sc_hd__buf_1 _35996_ (.A(_24058_),
    .X(_05540_));
 sky130_fd_sc_hd__nand4_4 _35997_ (.A(_23785_),
    .B(_05540_),
    .C(_24107_),
    .D(_24124_),
    .Y(_05541_));
 sky130_fd_sc_hd__o21ai_4 _35998_ (.A1(_05534_),
    .A2(_05535_),
    .B1(_04643_),
    .Y(_05542_));
 sky130_fd_sc_hd__a21oi_4 _35999_ (.A1(_05541_),
    .A2(_05542_),
    .B1(_05539_),
    .Y(_00292_));
 sky130_fd_sc_hd__o21a_4 _36000_ (.A1(_24053_),
    .A2(_24054_),
    .B1(instr_sltu),
    .X(_05543_));
 sky130_fd_sc_hd__nand3_4 _36001_ (.A(_18878_),
    .B(_24123_),
    .C(_23831_),
    .Y(_05544_));
 sky130_fd_sc_hd__nor2_4 _36002_ (.A(_05544_),
    .B(_05527_),
    .Y(_05545_));
 sky130_fd_sc_hd__o21a_4 _36003_ (.A1(_05543_),
    .A2(_05545_),
    .B1(_23379_),
    .X(_00283_));
 sky130_fd_sc_hd__nand4_4 _36004_ (.A(_23785_),
    .B(_05540_),
    .C(_24107_),
    .D(_24081_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21ai_4 _36005_ (.A1(_05534_),
    .A2(_05535_),
    .B1(instr_slt),
    .Y(_05547_));
 sky130_fd_sc_hd__a21oi_4 _36006_ (.A1(_05546_),
    .A2(_05547_),
    .B1(_05539_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand4_4 _36007_ (.A(_23785_),
    .B(_05540_),
    .C(_24107_),
    .D(_24118_),
    .Y(_05548_));
 sky130_fd_sc_hd__buf_1 _36008_ (.A(_24053_),
    .X(_05549_));
 sky130_fd_sc_hd__buf_1 _36009_ (.A(_24054_),
    .X(_05550_));
 sky130_fd_sc_hd__o21ai_4 _36010_ (.A1(_05549_),
    .A2(_05550_),
    .B1(_04615_),
    .Y(_05551_));
 sky130_fd_sc_hd__a21oi_4 _36011_ (.A1(_05548_),
    .A2(_05551_),
    .B1(_05539_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand4_4 _36012_ (.A(_23784_),
    .B(_23822_),
    .C(_23815_),
    .D(_24062_),
    .Y(_05552_));
 sky130_fd_sc_hd__buf_1 _36013_ (.A(_18354_),
    .X(_05553_));
 sky130_fd_sc_hd__o21ai_4 _36014_ (.A1(_05549_),
    .A2(_05550_),
    .B1(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__buf_1 _36015_ (.A(_19426_),
    .X(_05555_));
 sky130_fd_sc_hd__a21oi_4 _36016_ (.A1(_05552_),
    .A2(_05554_),
    .B1(_05555_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand4_4 _36017_ (.A(_23784_),
    .B(_05540_),
    .C(_23815_),
    .D(_24062_),
    .Y(_05556_));
 sky130_fd_sc_hd__o21ai_4 _36018_ (.A1(_05549_),
    .A2(_05550_),
    .B1(instr_add),
    .Y(_05557_));
 sky130_fd_sc_hd__a21oi_4 _36019_ (.A1(_05556_),
    .A2(_05557_),
    .B1(_05555_),
    .Y(_00246_));
 sky130_fd_sc_hd__a2bb2o_4 _36020_ (.A1_N(_05526_),
    .A2_N(_23832_),
    .B1(instr_andi),
    .B2(_24115_),
    .X(_05558_));
 sky130_fd_sc_hd__and2_4 _36021_ (.A(_05558_),
    .B(_21335_),
    .X(_00249_));
 sky130_fd_sc_hd__a2bb2o_4 _36022_ (.A1_N(_05530_),
    .A2_N(_23832_),
    .B1(instr_ori),
    .B2(_24115_),
    .X(_05559_));
 sky130_fd_sc_hd__and2_4 _36023_ (.A(_05559_),
    .B(_23063_),
    .X(_00269_));
 sky130_fd_sc_hd__buf_1 _36024_ (.A(_24102_),
    .X(_05560_));
 sky130_fd_sc_hd__nand3_4 _36025_ (.A(_24124_),
    .B(_23793_),
    .C(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21ai_4 _36026_ (.A1(_05549_),
    .A2(_05550_),
    .B1(_04644_),
    .Y(_05562_));
 sky130_fd_sc_hd__a21oi_4 _36027_ (.A1(_05561_),
    .A2(_05562_),
    .B1(_05555_),
    .Y(_00293_));
 sky130_fd_sc_hd__a2bb2o_4 _36028_ (.A1_N(_05544_),
    .A2_N(_23832_),
    .B1(instr_sltiu),
    .B2(_24115_),
    .X(_05563_));
 sky130_fd_sc_hd__and2_4 _36029_ (.A(_05563_),
    .B(_23063_),
    .X(_00282_));
 sky130_fd_sc_hd__nand3_4 _36030_ (.A(_24081_),
    .B(_23793_),
    .C(_05560_),
    .Y(_05564_));
 sky130_fd_sc_hd__buf_1 _36031_ (.A(_24078_),
    .X(_05565_));
 sky130_fd_sc_hd__buf_1 _36032_ (.A(_21959_),
    .X(_05566_));
 sky130_fd_sc_hd__o21ai_4 _36033_ (.A1(_05565_),
    .A2(_05566_),
    .B1(instr_slti),
    .Y(_05567_));
 sky130_fd_sc_hd__a21oi_4 _36034_ (.A1(_05564_),
    .A2(_05567_),
    .B1(_05555_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand3_4 _36035_ (.A(_24120_),
    .B(_23793_),
    .C(_05560_),
    .Y(_05568_));
 sky130_fd_sc_hd__o21ai_4 _36036_ (.A1(_05565_),
    .A2(_05566_),
    .B1(instr_addi),
    .Y(_05569_));
 sky130_fd_sc_hd__buf_1 _36037_ (.A(_19426_),
    .X(_05570_));
 sky130_fd_sc_hd__a21oi_4 _36038_ (.A1(_05568_),
    .A2(_05569_),
    .B1(_05570_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_4 _36039_ (.A(_24005_),
    .B(_24008_),
    .Y(_05571_));
 sky130_fd_sc_hd__o22a_4 _36040_ (.A1(_18329_),
    .A2(_23853_),
    .B1(_05526_),
    .B2(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__nor2_4 _36041_ (.A(_19427_),
    .B(_05572_),
    .Y(_00253_));
 sky130_fd_sc_hd__a2bb2o_4 _36042_ (.A1_N(_05530_),
    .A2_N(_05571_),
    .B1(instr_bltu),
    .B2(_24100_),
    .X(_05573_));
 sky130_fd_sc_hd__and2_4 _36043_ (.A(_05573_),
    .B(_23063_),
    .X(_00255_));
 sky130_fd_sc_hd__nand4_4 _36044_ (.A(_05520_),
    .B(_24103_),
    .C(_23809_),
    .D(_23824_),
    .Y(_05574_));
 sky130_fd_sc_hd__o21ai_4 _36045_ (.A1(_05565_),
    .A2(_05566_),
    .B1(instr_bge),
    .Y(_05575_));
 sky130_fd_sc_hd__a21oi_4 _36046_ (.A1(_05574_),
    .A2(_05575_),
    .B1(_05570_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand3_4 _36047_ (.A(_24124_),
    .B(_05520_),
    .C(_05560_),
    .Y(_05576_));
 sky130_fd_sc_hd__o21ai_4 _36048_ (.A1(_05565_),
    .A2(_05566_),
    .B1(instr_blt),
    .Y(_05577_));
 sky130_fd_sc_hd__a21oi_4 _36049_ (.A1(_05576_),
    .A2(_05577_),
    .B1(_05570_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand3_4 _36050_ (.A(_24118_),
    .B(_05520_),
    .C(_24103_),
    .Y(_05578_));
 sky130_fd_sc_hd__o21ai_4 _36051_ (.A1(_05523_),
    .A2(_05524_),
    .B1(instr_bne),
    .Y(_05579_));
 sky130_fd_sc_hd__a21oi_4 _36052_ (.A1(_05578_),
    .A2(_05579_),
    .B1(_05570_),
    .Y(_00256_));
 sky130_fd_sc_hd__nand3_4 _36053_ (.A(_24120_),
    .B(_24008_),
    .C(_24103_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ai_4 _36054_ (.A1(_05523_),
    .A2(_05524_),
    .B1(instr_beq),
    .Y(_05581_));
 sky130_fd_sc_hd__a21oi_4 _36055_ (.A1(_05580_),
    .A2(_05581_),
    .B1(_18784_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_4 _36056_ (.A(_19126_),
    .B(\pcpi_mul.active[0] ),
    .Y(_05582_));
 sky130_vsdinv _36057_ (.A(_05582_),
    .Y(_00670_));
 sky130_fd_sc_hd__buf_1 _36058_ (.A(\pcpi_mul.rs1[0] ),
    .X(_05583_));
 sky130_fd_sc_hd__buf_1 _36059_ (.A(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__buf_1 _36060_ (.A(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__buf_1 _36061_ (.A(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_1 _36062_ (.A(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_1 _36063_ (.A(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__buf_1 _36064_ (.A(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__nand2_4 _36065_ (.A(_05589_),
    .B(_03422_),
    .Y(_05590_));
 sky130_vsdinv _36066_ (.A(_05590_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2_4 _36067_ (.A(instr_sub),
    .B(_18627_),
    .Y(_05591_));
 sky130_fd_sc_hd__xnor2_4 _36068_ (.A(mem_la_wdata[1]),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__xor2_4 _36069_ (.A(_21380_),
    .B(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__xor2_4 _36070_ (.A(_04546_),
    .B(_05593_),
    .X(_01388_));
 sky130_fd_sc_hd__nor2_4 _36071_ (.A(mem_la_wdata[0]),
    .B(mem_la_wdata[1]),
    .Y(_05594_));
 sky130_fd_sc_hd__buf_1 _36072_ (.A(_05594_),
    .X(_05595_));
 sky130_vsdinv _36073_ (.A(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__nand3_4 _36074_ (.A(_05596_),
    .B(instr_sub),
    .C(_18614_),
    .Y(_05597_));
 sky130_vsdinv _36075_ (.A(instr_sub),
    .Y(_05598_));
 sky130_fd_sc_hd__o21ai_4 _36076_ (.A1(_05598_),
    .A2(_05595_),
    .B1(_21140_),
    .Y(_05599_));
 sky130_fd_sc_hd__a21o_4 _36077_ (.A1(_05597_),
    .A2(_05599_),
    .B1(pcpi_rs1[2]),
    .X(_05600_));
 sky130_fd_sc_hd__nand3_4 _36078_ (.A(_05597_),
    .B(_05599_),
    .C(_18612_),
    .Y(_05601_));
 sky130_fd_sc_hd__nand2_4 _36079_ (.A(_05600_),
    .B(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__maj3_4 _36080_ (.A(pcpi_rs1[1]),
    .B(_05592_),
    .C(_18634_),
    .X(_05603_));
 sky130_fd_sc_hd__xnor2_4 _36081_ (.A(_05602_),
    .B(_05603_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor3_4 _36082_ (.A(_18627_),
    .B(_18621_),
    .C(mem_la_wdata[2]),
    .Y(_05604_));
 sky130_vsdinv _36083_ (.A(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand3_4 _36084_ (.A(_05605_),
    .B(_18347_),
    .C(mem_la_wdata[3]),
    .Y(_05606_));
 sky130_fd_sc_hd__buf_1 _36085_ (.A(_05598_),
    .X(_05607_));
 sky130_fd_sc_hd__o21ai_4 _36086_ (.A1(_05607_),
    .A2(_05604_),
    .B1(_21152_),
    .Y(_05608_));
 sky130_fd_sc_hd__a21o_4 _36087_ (.A1(_05606_),
    .A2(_05608_),
    .B1(_21421_),
    .X(_05609_));
 sky130_fd_sc_hd__nand3_4 _36088_ (.A(_05606_),
    .B(_05608_),
    .C(_18607_),
    .Y(_05610_));
 sky130_fd_sc_hd__and2_4 _36089_ (.A(_05609_),
    .B(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__a21boi_4 _36090_ (.A1(_05603_),
    .A2(_05600_),
    .B1_N(_05601_),
    .Y(_05612_));
 sky130_fd_sc_hd__xor2_4 _36091_ (.A(_05611_),
    .B(_05612_),
    .X(_05613_));
 sky130_vsdinv _36092_ (.A(_05613_),
    .Y(_01402_));
 sky130_fd_sc_hd__nand4_4 _36093_ (.A(_21108_),
    .B(_21122_),
    .C(_21151_),
    .D(_21139_),
    .Y(_05614_));
 sky130_fd_sc_hd__a21o_4 _36094_ (.A1(_05614_),
    .A2(_18346_),
    .B1(mem_la_wdata[4]),
    .X(_05615_));
 sky130_fd_sc_hd__buf_1 _36095_ (.A(_05614_),
    .X(_05616_));
 sky130_fd_sc_hd__nand3_4 _36096_ (.A(_05616_),
    .B(_18346_),
    .C(_18601_),
    .Y(_05617_));
 sky130_fd_sc_hd__a21oi_4 _36097_ (.A1(_05615_),
    .A2(_05617_),
    .B1(_18599_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand3_4 _36098_ (.A(_05615_),
    .B(pcpi_rs1[4]),
    .C(_05617_),
    .Y(_05619_));
 sky130_vsdinv _36099_ (.A(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__nor2_4 _36100_ (.A(_05618_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__a21oi_4 _36101_ (.A1(_05606_),
    .A2(_05608_),
    .B1(pcpi_rs1[3]),
    .Y(_05622_));
 sky130_fd_sc_hd__o21ai_4 _36102_ (.A1(_05622_),
    .A2(_05612_),
    .B1(_05610_),
    .Y(_05623_));
 sky130_fd_sc_hd__xor2_4 _36103_ (.A(_05621_),
    .B(_05623_),
    .X(_01403_));
 sky130_fd_sc_hd__buf_1 _36104_ (.A(_05598_),
    .X(_05624_));
 sky130_fd_sc_hd__buf_1 _36105_ (.A(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__and4_4 _36106_ (.A(_05594_),
    .B(_21151_),
    .C(_21139_),
    .D(_21165_),
    .X(_05626_));
 sky130_fd_sc_hd__or3_4 _36107_ (.A(_05625_),
    .B(_21178_),
    .C(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__o21ai_4 _36108_ (.A1(_05625_),
    .A2(_05626_),
    .B1(_21178_),
    .Y(_05628_));
 sky130_fd_sc_hd__a21o_4 _36109_ (.A1(_05627_),
    .A2(_05628_),
    .B1(_18581_),
    .X(_05629_));
 sky130_fd_sc_hd__nand3_4 _36110_ (.A(_05627_),
    .B(_05628_),
    .C(pcpi_rs1[5]),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_4 _36111_ (.A(_05629_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__a21oi_4 _36112_ (.A1(_05623_),
    .A2(_05621_),
    .B1(_05620_),
    .Y(_05632_));
 sky130_fd_sc_hd__xor2_4 _36113_ (.A(_05631_),
    .B(_05632_),
    .X(_01404_));
 sky130_fd_sc_hd__nand2_4 _36114_ (.A(_05623_),
    .B(_05621_),
    .Y(_05633_));
 sky130_fd_sc_hd__nand3_4 _36115_ (.A(_05633_),
    .B(_05619_),
    .C(_05630_),
    .Y(_05634_));
 sky130_fd_sc_hd__nor3_4 _36116_ (.A(mem_la_wdata[5]),
    .B(_18601_),
    .C(_05616_),
    .Y(_05635_));
 sky130_fd_sc_hd__o21ai_4 _36117_ (.A1(_05624_),
    .A2(_05635_),
    .B1(_21189_),
    .Y(_05636_));
 sky130_fd_sc_hd__a41oi_4 _36118_ (.A1(_21152_),
    .A2(_05604_),
    .A3(_21178_),
    .A4(_21165_),
    .B1(_05607_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_4 _36119_ (.A(_05637_),
    .B(mem_la_wdata[6]),
    .Y(_05638_));
 sky130_fd_sc_hd__and2_4 _36120_ (.A(_05636_),
    .B(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__xor2_4 _36121_ (.A(_21470_),
    .B(_05639_),
    .X(_05640_));
 sky130_vsdinv _36122_ (.A(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__a21o_4 _36123_ (.A1(_05634_),
    .A2(_05629_),
    .B1(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__nand3_4 _36124_ (.A(_05634_),
    .B(_05629_),
    .C(_05641_),
    .Y(_05643_));
 sky130_fd_sc_hd__and2_4 _36125_ (.A(_05642_),
    .B(_05643_),
    .X(_01405_));
 sky130_fd_sc_hd__nor4_4 _36126_ (.A(mem_la_wdata[6]),
    .B(mem_la_wdata[5]),
    .C(mem_la_wdata[4]),
    .D(_05614_),
    .Y(_05644_));
 sky130_fd_sc_hd__nor3_4 _36127_ (.A(_05624_),
    .B(_21197_),
    .C(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__o21a_4 _36128_ (.A1(_05607_),
    .A2(_05644_),
    .B1(_21197_),
    .X(_05646_));
 sky130_fd_sc_hd__nor2_4 _36129_ (.A(_05645_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__xor2_4 _36130_ (.A(_21486_),
    .B(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__nand3_4 _36131_ (.A(_05636_),
    .B(_05638_),
    .C(pcpi_rs1[6]),
    .Y(_05649_));
 sky130_fd_sc_hd__nand2_4 _36132_ (.A(_05643_),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__xnor2_4 _36133_ (.A(_05648_),
    .B(_05650_),
    .Y(_01406_));
 sky130_fd_sc_hd__a211o_4 _36134_ (.A1(_05644_),
    .A2(_21196_),
    .B1(_05624_),
    .C1(_18661_),
    .X(_05651_));
 sky130_fd_sc_hd__a41o_4 _36135_ (.A1(_05626_),
    .A2(_21196_),
    .A3(_21189_),
    .A4(_21177_),
    .B1(_05607_),
    .X(_05652_));
 sky130_fd_sc_hd__nand2_4 _36136_ (.A(_05652_),
    .B(_18661_),
    .Y(_05653_));
 sky130_fd_sc_hd__a21oi_4 _36137_ (.A1(_05651_),
    .A2(_05653_),
    .B1(_21505_),
    .Y(_05654_));
 sky130_vsdinv _36138_ (.A(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__nand3_4 _36139_ (.A(_05651_),
    .B(_21505_),
    .C(_05653_),
    .Y(_05656_));
 sky130_fd_sc_hd__and2_4 _36140_ (.A(_05655_),
    .B(_05656_),
    .X(_05657_));
 sky130_vsdinv _36141_ (.A(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__nor2_4 _36142_ (.A(_05640_),
    .B(_05648_),
    .Y(_05659_));
 sky130_fd_sc_hd__nand3_4 _36143_ (.A(_05634_),
    .B(_05659_),
    .C(_05629_),
    .Y(_05660_));
 sky130_fd_sc_hd__a21bo_4 _36144_ (.A1(_05647_),
    .A2(_18587_),
    .B1_N(_05649_),
    .X(_05661_));
 sky130_fd_sc_hd__o21ai_4 _36145_ (.A1(_18587_),
    .A2(_05647_),
    .B1(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__and2_4 _36146_ (.A(_05660_),
    .B(_05662_),
    .X(_05663_));
 sky130_fd_sc_hd__buf_1 _36147_ (.A(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__xor2_4 _36148_ (.A(_05658_),
    .B(_05664_),
    .X(_01407_));
 sky130_fd_sc_hd__nand2_4 _36149_ (.A(_18346_),
    .B(pcpi_rs2[8]),
    .Y(_05665_));
 sky130_fd_sc_hd__a21o_4 _36150_ (.A1(_05652_),
    .A2(_05665_),
    .B1(_21210_),
    .X(_05666_));
 sky130_fd_sc_hd__nand3_4 _36151_ (.A(_05652_),
    .B(_21211_),
    .C(_05665_),
    .Y(_05667_));
 sky130_fd_sc_hd__a21oi_4 _36152_ (.A1(_05666_),
    .A2(_05667_),
    .B1(pcpi_rs1[9]),
    .Y(_05668_));
 sky130_vsdinv _36153_ (.A(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand3_4 _36154_ (.A(_05666_),
    .B(_18650_),
    .C(_05667_),
    .Y(_05670_));
 sky130_fd_sc_hd__and2_4 _36155_ (.A(_05669_),
    .B(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__o21ai_4 _36156_ (.A1(_05658_),
    .A2(_05664_),
    .B1(_05655_),
    .Y(_05672_));
 sky130_fd_sc_hd__xor2_4 _36157_ (.A(_05671_),
    .B(_05672_),
    .X(_01408_));
 sky130_fd_sc_hd__nand4_4 _36158_ (.A(_21197_),
    .B(_05644_),
    .C(_21211_),
    .D(_21204_),
    .Y(_05673_));
 sky130_fd_sc_hd__buf_1 _36159_ (.A(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__a21o_4 _36160_ (.A1(_05674_),
    .A2(_18347_),
    .B1(pcpi_rs2[10]),
    .X(_05675_));
 sky130_fd_sc_hd__nand3_4 _36161_ (.A(_05674_),
    .B(_18347_),
    .C(pcpi_rs2[10]),
    .Y(_05676_));
 sky130_fd_sc_hd__nand3_4 _36162_ (.A(_05675_),
    .B(pcpi_rs1[10]),
    .C(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__a21o_4 _36163_ (.A1(_05675_),
    .A2(_05676_),
    .B1(pcpi_rs1[10]),
    .X(_05678_));
 sky130_fd_sc_hd__a21oi_4 _36164_ (.A1(_05655_),
    .A2(_05670_),
    .B1(_05668_),
    .Y(_05679_));
 sky130_fd_sc_hd__and4_4 _36165_ (.A(_05669_),
    .B(_05655_),
    .C(_05656_),
    .D(_05670_),
    .X(_05680_));
 sky130_vsdinv _36166_ (.A(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__a21oi_4 _36167_ (.A1(_05660_),
    .A2(_05662_),
    .B1(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__a211o_4 _36168_ (.A1(_05677_),
    .A2(_05678_),
    .B1(_05679_),
    .C1(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__and2_4 _36169_ (.A(_05678_),
    .B(_05677_),
    .X(_05684_));
 sky130_fd_sc_hd__o21ai_4 _36170_ (.A1(_05679_),
    .A2(_05682_),
    .B1(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__and2_4 _36171_ (.A(_05683_),
    .B(_05685_),
    .X(_01378_));
 sky130_fd_sc_hd__nor2_4 _36172_ (.A(pcpi_rs2[10]),
    .B(_05673_),
    .Y(_05686_));
 sky130_vsdinv _36173_ (.A(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__nand3_4 _36174_ (.A(_05687_),
    .B(_18348_),
    .C(_18658_),
    .Y(_05688_));
 sky130_fd_sc_hd__o21ai_4 _36175_ (.A1(_05625_),
    .A2(_05686_),
    .B1(_21230_),
    .Y(_05689_));
 sky130_fd_sc_hd__a21oi_4 _36176_ (.A1(_05688_),
    .A2(_05689_),
    .B1(_18656_),
    .Y(_05690_));
 sky130_fd_sc_hd__nand3_4 _36177_ (.A(_05688_),
    .B(_05689_),
    .C(pcpi_rs1[11]),
    .Y(_05691_));
 sky130_vsdinv _36178_ (.A(_05691_),
    .Y(_05692_));
 sky130_fd_sc_hd__nor2_4 _36179_ (.A(_05690_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand2_4 _36180_ (.A(_05685_),
    .B(_05677_),
    .Y(_05694_));
 sky130_fd_sc_hd__xor2_4 _36181_ (.A(_05693_),
    .B(_05694_),
    .X(_01379_));
 sky130_fd_sc_hd__buf_1 _36182_ (.A(_05625_),
    .X(_05695_));
 sky130_fd_sc_hd__nor3_4 _36183_ (.A(pcpi_rs2[11]),
    .B(_18654_),
    .C(_05674_),
    .Y(_05696_));
 sky130_fd_sc_hd__o21ai_4 _36184_ (.A1(_05695_),
    .A2(_05696_),
    .B1(_21236_),
    .Y(_05697_));
 sky130_vsdinv _36185_ (.A(_05696_),
    .Y(_05698_));
 sky130_fd_sc_hd__nand3_4 _36186_ (.A(_05698_),
    .B(_18348_),
    .C(_18647_),
    .Y(_05699_));
 sky130_fd_sc_hd__a21o_4 _36187_ (.A1(_05697_),
    .A2(_05699_),
    .B1(_18645_),
    .X(_05700_));
 sky130_fd_sc_hd__nand3_4 _36188_ (.A(_05699_),
    .B(_05697_),
    .C(pcpi_rs1[12]),
    .Y(_05701_));
 sky130_fd_sc_hd__and2_4 _36189_ (.A(_05700_),
    .B(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__a211o_4 _36190_ (.A1(_05694_),
    .A2(_05693_),
    .B1(_05692_),
    .C1(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__a21boi_4 _36191_ (.A1(_05685_),
    .A2(_05677_),
    .B1_N(_05693_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21ai_4 _36192_ (.A1(_05692_),
    .A2(_05704_),
    .B1(_05702_),
    .Y(_05705_));
 sky130_fd_sc_hd__and2_4 _36193_ (.A(_05703_),
    .B(_05705_),
    .X(_01380_));
 sky130_fd_sc_hd__nor4_4 _36194_ (.A(pcpi_rs2[12]),
    .B(pcpi_rs2[11]),
    .C(_18654_),
    .D(_05674_),
    .Y(_05706_));
 sky130_vsdinv _36195_ (.A(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand3_4 _36196_ (.A(_05707_),
    .B(_18348_),
    .C(pcpi_rs2[13]),
    .Y(_05708_));
 sky130_fd_sc_hd__o21ai_4 _36197_ (.A1(_05695_),
    .A2(_05706_),
    .B1(_21243_),
    .Y(_05709_));
 sky130_fd_sc_hd__a21oi_4 _36198_ (.A1(_05708_),
    .A2(_05709_),
    .B1(pcpi_rs1[13]),
    .Y(_05710_));
 sky130_fd_sc_hd__nand3_4 _36199_ (.A(_05708_),
    .B(_05709_),
    .C(pcpi_rs1[13]),
    .Y(_05711_));
 sky130_vsdinv _36200_ (.A(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__nor2_4 _36201_ (.A(_05710_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_4 _36202_ (.A(_05705_),
    .B(_05701_),
    .Y(_05714_));
 sky130_fd_sc_hd__xor2_4 _36203_ (.A(_05713_),
    .B(_05714_),
    .X(_01381_));
 sky130_fd_sc_hd__and4_4 _36204_ (.A(_05686_),
    .B(_21243_),
    .C(_21236_),
    .D(_21230_),
    .X(_05715_));
 sky130_vsdinv _36205_ (.A(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__nand3_4 _36206_ (.A(_05716_),
    .B(_18349_),
    .C(pcpi_rs2[14]),
    .Y(_05717_));
 sky130_fd_sc_hd__buf_1 _36207_ (.A(_05695_),
    .X(_05718_));
 sky130_fd_sc_hd__o21ai_4 _36208_ (.A1(_05718_),
    .A2(_05715_),
    .B1(_21250_),
    .Y(_05719_));
 sky130_fd_sc_hd__a21o_4 _36209_ (.A1(_05717_),
    .A2(_05719_),
    .B1(_18637_),
    .X(_05720_));
 sky130_fd_sc_hd__nand3_4 _36210_ (.A(_05717_),
    .B(_05719_),
    .C(pcpi_rs1[14]),
    .Y(_05721_));
 sky130_fd_sc_hd__and2_4 _36211_ (.A(_05720_),
    .B(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__a211o_4 _36212_ (.A1(_05714_),
    .A2(_05713_),
    .B1(_05712_),
    .C1(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__a21boi_4 _36213_ (.A1(_05705_),
    .A2(_05701_),
    .B1_N(_05713_),
    .Y(_05724_));
 sky130_fd_sc_hd__o21ai_4 _36214_ (.A1(_05712_),
    .A2(_05724_),
    .B1(_05722_),
    .Y(_05725_));
 sky130_fd_sc_hd__and2_4 _36215_ (.A(_05723_),
    .B(_05725_),
    .X(_01382_));
 sky130_fd_sc_hd__and4_4 _36216_ (.A(_05696_),
    .B(_21248_),
    .C(_21242_),
    .D(_21235_),
    .X(_05726_));
 sky130_vsdinv _36217_ (.A(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__a21o_4 _36218_ (.A1(_05727_),
    .A2(_18349_),
    .B1(_18643_),
    .X(_05728_));
 sky130_fd_sc_hd__nand3_4 _36219_ (.A(_05727_),
    .B(_18350_),
    .C(_18643_),
    .Y(_05729_));
 sky130_fd_sc_hd__a21oi_4 _36220_ (.A1(_05728_),
    .A2(_05729_),
    .B1(pcpi_rs1[15]),
    .Y(_05730_));
 sky130_fd_sc_hd__nand3_4 _36221_ (.A(_05728_),
    .B(pcpi_rs1[15]),
    .C(_05729_),
    .Y(_05731_));
 sky130_vsdinv _36222_ (.A(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__nor2_4 _36223_ (.A(_05730_),
    .B(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__nand2_4 _36224_ (.A(_05725_),
    .B(_05721_),
    .Y(_05734_));
 sky130_fd_sc_hd__xor2_4 _36225_ (.A(_05733_),
    .B(_05734_),
    .X(_01383_));
 sky130_fd_sc_hd__a41oi_4 _36226_ (.A1(_21256_),
    .A2(_05706_),
    .A3(_21249_),
    .A4(_21244_),
    .B1(_05695_),
    .Y(_05735_));
 sky130_fd_sc_hd__xor2_4 _36227_ (.A(_18711_),
    .B(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__xor2_4 _36228_ (.A(pcpi_rs1[16]),
    .B(_05736_),
    .X(_05737_));
 sky130_vsdinv _36229_ (.A(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__a21oi_4 _36230_ (.A1(_05734_),
    .A2(_05733_),
    .B1(_05732_),
    .Y(_05739_));
 sky130_fd_sc_hd__xor2_4 _36231_ (.A(_05738_),
    .B(_05739_),
    .X(_01384_));
 sky130_fd_sc_hd__and4_4 _36232_ (.A(_05706_),
    .B(_21256_),
    .C(_21249_),
    .D(_21243_),
    .X(_05740_));
 sky130_fd_sc_hd__a211o_4 _36233_ (.A1(_05740_),
    .A2(_21262_),
    .B1(_05718_),
    .C1(_21267_),
    .X(_05741_));
 sky130_fd_sc_hd__a211o_4 _36234_ (.A1(_18349_),
    .A2(_18711_),
    .B1(_18716_),
    .C1(_05735_),
    .X(_05742_));
 sky130_fd_sc_hd__nand2_4 _36235_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_4 _36236_ (.A(_05743_),
    .B(_21670_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand3_4 _36237_ (.A(_05741_),
    .B(_05742_),
    .C(pcpi_rs1[17]),
    .Y(_05745_));
 sky130_fd_sc_hd__and2_4 _36238_ (.A(_05744_),
    .B(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__nand2_4 _36239_ (.A(_05736_),
    .B(_18709_),
    .Y(_05747_));
 sky130_fd_sc_hd__o21ai_4 _36240_ (.A1(_05738_),
    .A2(_05739_),
    .B1(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__xor2_4 _36241_ (.A(_05746_),
    .B(_05748_),
    .X(_01385_));
 sky130_fd_sc_hd__nor2_4 _36242_ (.A(_18716_),
    .B(pcpi_rs2[16]),
    .Y(_05749_));
 sky130_fd_sc_hd__and4_4 _36243_ (.A(_05715_),
    .B(_21256_),
    .C(_21249_),
    .D(_05749_),
    .X(_05750_));
 sky130_vsdinv _36244_ (.A(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__nand3_4 _36245_ (.A(_05751_),
    .B(_18350_),
    .C(pcpi_rs2[18]),
    .Y(_05752_));
 sky130_fd_sc_hd__o21ai_4 _36246_ (.A1(_05718_),
    .A2(_05750_),
    .B1(_18702_),
    .Y(_05753_));
 sky130_fd_sc_hd__a21oi_4 _36247_ (.A1(_05752_),
    .A2(_05753_),
    .B1(pcpi_rs1[18]),
    .Y(_05754_));
 sky130_fd_sc_hd__nand3_4 _36248_ (.A(_05752_),
    .B(_05753_),
    .C(pcpi_rs1[18]),
    .Y(_05755_));
 sky130_vsdinv _36249_ (.A(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__nor2_4 _36250_ (.A(_05754_),
    .B(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__a21boi_4 _36251_ (.A1(_05725_),
    .A2(_05721_),
    .B1_N(_05733_),
    .Y(_05758_));
 sky130_fd_sc_hd__and2_4 _36252_ (.A(_05746_),
    .B(_05737_),
    .X(_05759_));
 sky130_fd_sc_hd__o21ai_4 _36253_ (.A1(_05732_),
    .A2(_05758_),
    .B1(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__a21bo_4 _36254_ (.A1(_05747_),
    .A2(_05745_),
    .B1_N(_05744_),
    .X(_05761_));
 sky130_fd_sc_hd__nand2_4 _36255_ (.A(_05760_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__xor2_4 _36256_ (.A(_05757_),
    .B(_05762_),
    .X(_01386_));
 sky130_fd_sc_hd__nand4_4 _36257_ (.A(_21257_),
    .B(_05726_),
    .C(_18703_),
    .D(_05749_),
    .Y(_05763_));
 sky130_fd_sc_hd__a21o_4 _36258_ (.A1(_05763_),
    .A2(_18350_),
    .B1(_18695_),
    .X(_05764_));
 sky130_fd_sc_hd__nand3_4 _36259_ (.A(_05763_),
    .B(_18351_),
    .C(_18695_),
    .Y(_05765_));
 sky130_fd_sc_hd__a21o_4 _36260_ (.A1(_05764_),
    .A2(_05765_),
    .B1(pcpi_rs1[19]),
    .X(_05766_));
 sky130_fd_sc_hd__nand3_4 _36261_ (.A(_05764_),
    .B(pcpi_rs1[19]),
    .C(_05765_),
    .Y(_05767_));
 sky130_fd_sc_hd__and2_4 _36262_ (.A(_05766_),
    .B(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__a211o_4 _36263_ (.A1(_05762_),
    .A2(_05757_),
    .B1(_05756_),
    .C1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__a21boi_4 _36264_ (.A1(_05760_),
    .A2(_05761_),
    .B1_N(_05757_),
    .Y(_05770_));
 sky130_fd_sc_hd__o21ai_4 _36265_ (.A1(_05756_),
    .A2(_05770_),
    .B1(_05768_),
    .Y(_05771_));
 sky130_fd_sc_hd__and2_4 _36266_ (.A(_05769_),
    .B(_05771_),
    .X(_01387_));
 sky130_fd_sc_hd__nand4_4 _36267_ (.A(_21277_),
    .B(_05740_),
    .C(_18703_),
    .D(_05749_),
    .Y(_05772_));
 sky130_fd_sc_hd__a21o_4 _36268_ (.A1(_05772_),
    .A2(_18351_),
    .B1(pcpi_rs2[20]),
    .X(_05773_));
 sky130_fd_sc_hd__buf_1 _36269_ (.A(_05772_),
    .X(_05774_));
 sky130_fd_sc_hd__nand3_4 _36270_ (.A(_05774_),
    .B(_18351_),
    .C(pcpi_rs2[20]),
    .Y(_05775_));
 sky130_fd_sc_hd__a21oi_4 _36271_ (.A1(_05773_),
    .A2(_05775_),
    .B1(_18665_),
    .Y(_05776_));
 sky130_fd_sc_hd__nand3_4 _36272_ (.A(_05773_),
    .B(pcpi_rs1[20]),
    .C(_05775_),
    .Y(_05777_));
 sky130_vsdinv _36273_ (.A(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__nor2_4 _36274_ (.A(_05776_),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_4 _36275_ (.A(_05771_),
    .B(_05767_),
    .Y(_05780_));
 sky130_fd_sc_hd__xor2_4 _36276_ (.A(_05779_),
    .B(_05780_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2_4 _36277_ (.A(_18667_),
    .B(_05774_),
    .Y(_05781_));
 sky130_vsdinv _36278_ (.A(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__nand3_4 _36279_ (.A(_05782_),
    .B(_18352_),
    .C(_18681_),
    .Y(_05783_));
 sky130_fd_sc_hd__buf_1 _36280_ (.A(_05718_),
    .X(_05784_));
 sky130_fd_sc_hd__o21ai_4 _36281_ (.A1(_05784_),
    .A2(_05781_),
    .B1(_21289_),
    .Y(_05785_));
 sky130_fd_sc_hd__a21oi_4 _36282_ (.A1(_05783_),
    .A2(_05785_),
    .B1(_18680_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand3_4 _36283_ (.A(_05783_),
    .B(_05785_),
    .C(_18680_),
    .Y(_05787_));
 sky130_vsdinv _36284_ (.A(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__nor2_4 _36285_ (.A(_05786_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__a21oi_4 _36286_ (.A1(_05780_),
    .A2(_05779_),
    .B1(_05778_),
    .Y(_05790_));
 sky130_fd_sc_hd__xnor2_4 _36287_ (.A(_05789_),
    .B(_05790_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor3_4 _36288_ (.A(pcpi_rs2[21]),
    .B(pcpi_rs2[20]),
    .C(_05774_),
    .Y(_05791_));
 sky130_vsdinv _36289_ (.A(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__nand3_4 _36290_ (.A(_05792_),
    .B(_18352_),
    .C(pcpi_rs2[22]),
    .Y(_05793_));
 sky130_fd_sc_hd__o21ai_4 _36291_ (.A1(_05784_),
    .A2(_05791_),
    .B1(_18674_),
    .Y(_05794_));
 sky130_fd_sc_hd__a21oi_4 _36292_ (.A1(_05793_),
    .A2(_05794_),
    .B1(_18672_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand3_4 _36293_ (.A(_05793_),
    .B(_05794_),
    .C(pcpi_rs1[22]),
    .Y(_05796_));
 sky130_vsdinv _36294_ (.A(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__nor2_4 _36295_ (.A(_05795_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__o21ai_4 _36296_ (.A1(_05786_),
    .A2(_05790_),
    .B1(_05787_),
    .Y(_05799_));
 sky130_fd_sc_hd__xor2_4 _36297_ (.A(_05798_),
    .B(_05799_),
    .X(_01391_));
 sky130_fd_sc_hd__nor4_4 _36298_ (.A(pcpi_rs2[22]),
    .B(_18681_),
    .C(_18667_),
    .D(_05774_),
    .Y(_05800_));
 sky130_vsdinv _36299_ (.A(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__nand3_4 _36300_ (.A(_05801_),
    .B(_18353_),
    .C(_18689_),
    .Y(_05802_));
 sky130_fd_sc_hd__buf_1 _36301_ (.A(_05784_),
    .X(_05803_));
 sky130_fd_sc_hd__o21ai_4 _36302_ (.A1(_05803_),
    .A2(_05800_),
    .B1(_21300_),
    .Y(_05804_));
 sky130_fd_sc_hd__a21oi_4 _36303_ (.A1(_05802_),
    .A2(_05804_),
    .B1(_18688_),
    .Y(_05805_));
 sky130_fd_sc_hd__nand3_4 _36304_ (.A(_05802_),
    .B(_05804_),
    .C(_01671_),
    .Y(_05806_));
 sky130_vsdinv _36305_ (.A(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__nor2_4 _36306_ (.A(_05805_),
    .B(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__a21oi_4 _36307_ (.A1(_05799_),
    .A2(_05798_),
    .B1(_05797_),
    .Y(_05809_));
 sky130_fd_sc_hd__xnor2_4 _36308_ (.A(_05808_),
    .B(_05809_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand4_4 _36309_ (.A(_21299_),
    .B(_05781_),
    .C(_18674_),
    .D(_21289_),
    .Y(_05810_));
 sky130_fd_sc_hd__a21o_4 _36310_ (.A1(_05810_),
    .A2(_18352_),
    .B1(_18733_),
    .X(_05811_));
 sky130_fd_sc_hd__nand3_4 _36311_ (.A(_05810_),
    .B(_18353_),
    .C(_18734_),
    .Y(_05812_));
 sky130_fd_sc_hd__a21o_4 _36312_ (.A1(_05811_),
    .A2(_05812_),
    .B1(_18731_),
    .X(_05813_));
 sky130_fd_sc_hd__nand3_4 _36313_ (.A(_05811_),
    .B(_18731_),
    .C(_05812_),
    .Y(_05814_));
 sky130_fd_sc_hd__and2_4 _36314_ (.A(_05813_),
    .B(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__o21ai_4 _36315_ (.A1(_05805_),
    .A2(_05809_),
    .B1(_05806_),
    .Y(_05816_));
 sky130_fd_sc_hd__xor2_4 _36316_ (.A(_05815_),
    .B(_05816_),
    .X(_01393_));
 sky130_fd_sc_hd__nor2_4 _36317_ (.A(pcpi_rs2[24]),
    .B(_05810_),
    .Y(_05817_));
 sky130_vsdinv _36318_ (.A(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand3_4 _36319_ (.A(_05818_),
    .B(_18353_),
    .C(pcpi_rs2[25]),
    .Y(_05819_));
 sky130_fd_sc_hd__o21ai_4 _36320_ (.A1(_05784_),
    .A2(_05817_),
    .B1(_21309_),
    .Y(_05820_));
 sky130_fd_sc_hd__a21o_4 _36321_ (.A1(_05819_),
    .A2(_05820_),
    .B1(_18765_),
    .X(_05821_));
 sky130_fd_sc_hd__nand3_4 _36322_ (.A(_05819_),
    .B(_05820_),
    .C(_18765_),
    .Y(_05822_));
 sky130_fd_sc_hd__nand2_4 _36323_ (.A(_05821_),
    .B(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__a21boi_4 _36324_ (.A1(_05816_),
    .A2(_05813_),
    .B1_N(_05814_),
    .Y(_05824_));
 sky130_fd_sc_hd__xor2_4 _36325_ (.A(_05823_),
    .B(_05824_),
    .X(_01394_));
 sky130_fd_sc_hd__and4_4 _36326_ (.A(_05800_),
    .B(_21308_),
    .C(_18729_),
    .D(_21300_),
    .X(_05825_));
 sky130_vsdinv _36327_ (.A(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__nand3_4 _36328_ (.A(_05826_),
    .B(_18354_),
    .C(pcpi_rs2[26]),
    .Y(_05827_));
 sky130_fd_sc_hd__o21ai_4 _36329_ (.A1(_05803_),
    .A2(_05825_),
    .B1(_21315_),
    .Y(_05828_));
 sky130_fd_sc_hd__a21oi_4 _36330_ (.A1(_05827_),
    .A2(_05828_),
    .B1(_18721_),
    .Y(_05829_));
 sky130_fd_sc_hd__nand3_4 _36331_ (.A(_05827_),
    .B(_05828_),
    .C(_18724_),
    .Y(_05830_));
 sky130_vsdinv _36332_ (.A(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__nor2_4 _36333_ (.A(_05829_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__and4_4 _36334_ (.A(_05821_),
    .B(_05814_),
    .C(_05813_),
    .D(_05822_),
    .X(_05833_));
 sky130_fd_sc_hd__a21boi_4 _36335_ (.A1(_05814_),
    .A2(_05822_),
    .B1_N(_05821_),
    .Y(_05834_));
 sky130_fd_sc_hd__a21oi_4 _36336_ (.A1(_05816_),
    .A2(_05833_),
    .B1(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__xnor2_4 _36337_ (.A(_05832_),
    .B(_05835_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor4_4 _36338_ (.A(pcpi_rs2[26]),
    .B(pcpi_rs2[25]),
    .C(_18733_),
    .D(_05810_),
    .Y(_05836_));
 sky130_vsdinv _36339_ (.A(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__buf_1 _36340_ (.A(_18354_),
    .X(_05838_));
 sky130_fd_sc_hd__nand3_4 _36341_ (.A(_05837_),
    .B(_05838_),
    .C(_18762_),
    .Y(_05839_));
 sky130_fd_sc_hd__o21ai_4 _36342_ (.A1(_05803_),
    .A2(_05836_),
    .B1(_18760_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_4 _36343_ (.A(_05839_),
    .B(_05840_),
    .Y(_05841_));
 sky130_fd_sc_hd__nand2_4 _36344_ (.A(_05841_),
    .B(_21822_),
    .Y(_05842_));
 sky130_fd_sc_hd__nand3_4 _36345_ (.A(_05839_),
    .B(_05840_),
    .C(_01689_),
    .Y(_05843_));
 sky130_fd_sc_hd__and2_4 _36346_ (.A(_05842_),
    .B(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__o21ai_4 _36347_ (.A1(_05829_),
    .A2(_05835_),
    .B1(_05830_),
    .Y(_05845_));
 sky130_fd_sc_hd__xor2_4 _36348_ (.A(_05844_),
    .B(_05845_),
    .X(_01396_));
 sky130_fd_sc_hd__and4_4 _36349_ (.A(_05817_),
    .B(_18759_),
    .C(_21314_),
    .D(_21309_),
    .X(_05846_));
 sky130_vsdinv _36350_ (.A(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__nand3_4 _36351_ (.A(_05847_),
    .B(_05553_),
    .C(_18747_),
    .Y(_05848_));
 sky130_fd_sc_hd__o21ai_4 _36352_ (.A1(_05803_),
    .A2(_05846_),
    .B1(_21325_),
    .Y(_05849_));
 sky130_fd_sc_hd__a21o_4 _36353_ (.A1(_05848_),
    .A2(_05849_),
    .B1(_01694_),
    .X(_05850_));
 sky130_fd_sc_hd__nand3_4 _36354_ (.A(_05848_),
    .B(_05849_),
    .C(_01694_),
    .Y(_05851_));
 sky130_fd_sc_hd__and2_4 _36355_ (.A(_05850_),
    .B(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__nand3_4 _36356_ (.A(_05832_),
    .B(_05843_),
    .C(_05842_),
    .Y(_05853_));
 sky130_fd_sc_hd__maj3_4 _36357_ (.A(_21822_),
    .B(_05841_),
    .C(_05830_),
    .X(_05854_));
 sky130_fd_sc_hd__o21ai_4 _36358_ (.A1(_05853_),
    .A2(_05835_),
    .B1(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__xor2_4 _36359_ (.A(_05852_),
    .B(_05855_),
    .X(_01397_));
 sky130_fd_sc_hd__nand4_4 _36360_ (.A(_21325_),
    .B(_05825_),
    .C(_18759_),
    .D(_21315_),
    .Y(_05856_));
 sky130_fd_sc_hd__a21o_4 _36361_ (.A1(_05856_),
    .A2(_05838_),
    .B1(_18752_),
    .X(_05857_));
 sky130_fd_sc_hd__nand3_4 _36362_ (.A(_05856_),
    .B(_05553_),
    .C(_01506_),
    .Y(_05858_));
 sky130_fd_sc_hd__a21o_4 _36363_ (.A1(_05857_),
    .A2(_05858_),
    .B1(_21855_),
    .X(_05859_));
 sky130_fd_sc_hd__nand3_4 _36364_ (.A(_05857_),
    .B(_21879_),
    .C(_05858_),
    .Y(_05860_));
 sky130_fd_sc_hd__nand2_4 _36365_ (.A(_05859_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__a21boi_4 _36366_ (.A1(_05855_),
    .A2(_05850_),
    .B1_N(_05851_),
    .Y(_05862_));
 sky130_fd_sc_hd__xor2_4 _36367_ (.A(_05861_),
    .B(_05862_),
    .X(_01398_));
 sky130_fd_sc_hd__nand4_4 _36368_ (.A(_21329_),
    .B(_05836_),
    .C(_21324_),
    .D(_18759_),
    .Y(_05863_));
 sky130_fd_sc_hd__a21o_4 _36369_ (.A1(_05863_),
    .A2(_05838_),
    .B1(_21334_),
    .X(_05864_));
 sky130_fd_sc_hd__nand3_4 _36370_ (.A(_05863_),
    .B(_05838_),
    .C(_21334_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21o_4 _36371_ (.A1(_05864_),
    .A2(_05865_),
    .B1(_21870_),
    .X(_05866_));
 sky130_fd_sc_hd__nand3_4 _36372_ (.A(_05864_),
    .B(_21870_),
    .C(_05865_),
    .Y(_05867_));
 sky130_fd_sc_hd__and2_4 _36373_ (.A(_05866_),
    .B(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__buf_1 _36374_ (.A(_05868_),
    .X(_05869_));
 sky130_vsdinv _36375_ (.A(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__and4_4 _36376_ (.A(_05859_),
    .B(_05850_),
    .C(_05851_),
    .D(_05860_),
    .X(_05871_));
 sky130_fd_sc_hd__a21boi_4 _36377_ (.A1(_05851_),
    .A2(_05860_),
    .B1_N(_05859_),
    .Y(_05872_));
 sky130_fd_sc_hd__a21oi_4 _36378_ (.A1(_05855_),
    .A2(_05871_),
    .B1(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__xor2_4 _36379_ (.A(_05870_),
    .B(_05873_),
    .X(_01400_));
 sky130_fd_sc_hd__o21ai_4 _36380_ (.A1(_05870_),
    .A2(_05873_),
    .B1(_05866_),
    .Y(_05874_));
 sky130_fd_sc_hd__o21a_4 _36381_ (.A1(_18737_),
    .A2(_05863_),
    .B1(_05553_),
    .X(_05875_));
 sky130_fd_sc_hd__xor2_4 _36382_ (.A(_05424_),
    .B(_05875_),
    .X(_05876_));
 sky130_vsdinv _36383_ (.A(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__nand2_4 _36384_ (.A(_05874_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__a21o_4 _36385_ (.A1(_05855_),
    .A2(_05871_),
    .B1(_05872_),
    .X(_05879_));
 sky130_fd_sc_hd__nand2_4 _36386_ (.A(_05879_),
    .B(_05869_),
    .Y(_05880_));
 sky130_fd_sc_hd__nand3_4 _36387_ (.A(_05880_),
    .B(_05866_),
    .C(_05876_),
    .Y(_05881_));
 sky130_fd_sc_hd__nand2_4 _36388_ (.A(_05878_),
    .B(_05881_),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_4 _36389_ (.A(_18632_),
    .B(_04546_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_4 _36390_ (.A(_05587_),
    .B(_03437_),
    .Y(_05882_));
 sky130_fd_sc_hd__buf_1 _36391_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05883_));
 sky130_fd_sc_hd__buf_1 _36392_ (.A(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__buf_1 _36393_ (.A(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__buf_1 _36394_ (.A(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__buf_1 _36395_ (.A(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__nand2_4 _36396_ (.A(_05887_),
    .B(_03422_),
    .Y(_05888_));
 sky130_fd_sc_hd__xnor2_4 _36397_ (.A(_05882_),
    .B(_05888_),
    .Y(_05889_));
 sky130_vsdinv _36398_ (.A(_05889_),
    .Y(_01410_));
 sky130_fd_sc_hd__nor2_4 _36399_ (.A(_05882_),
    .B(_05888_),
    .Y(_05890_));
 sky130_vsdinv _36400_ (.A(\pcpi_mul.rs2[1] ),
    .Y(_05891_));
 sky130_fd_sc_hd__buf_1 _36401_ (.A(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_1 _36402_ (.A(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__a2bb2o_4 _36403_ (.A1_N(_03250_),
    .A2_N(_05893_),
    .B1(_05587_),
    .B2(_03445_),
    .X(_05894_));
 sky130_fd_sc_hd__buf_1 _36404_ (.A(_03228_),
    .X(_05895_));
 sky130_fd_sc_hd__buf_1 _36405_ (.A(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__buf_1 _36406_ (.A(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__nand4_4 _36407_ (.A(_05897_),
    .B(_05887_),
    .C(_03437_),
    .D(_03445_),
    .Y(_05898_));
 sky130_fd_sc_hd__buf_1 _36408_ (.A(\pcpi_mul.rs1[2] ),
    .X(_05899_));
 sky130_fd_sc_hd__buf_1 _36409_ (.A(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__buf_1 _36410_ (.A(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_1 _36411_ (.A(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__nand2_4 _36412_ (.A(_05902_),
    .B(_03422_),
    .Y(_05903_));
 sky130_vsdinv _36413_ (.A(_05903_),
    .Y(_05904_));
 sky130_fd_sc_hd__a21o_4 _36414_ (.A1(_05894_),
    .A2(_05898_),
    .B1(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__nand3_4 _36415_ (.A(_05894_),
    .B(_05898_),
    .C(_05904_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand2_4 _36416_ (.A(_05905_),
    .B(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__xnor2_4 _36417_ (.A(_05890_),
    .B(_05907_),
    .Y(_01411_));
 sky130_fd_sc_hd__nand3_4 _36418_ (.A(_05905_),
    .B(_05890_),
    .C(_05906_),
    .Y(_05908_));
 sky130_fd_sc_hd__buf_1 _36419_ (.A(\pcpi_mul.rs2[2] ),
    .X(_05909_));
 sky130_fd_sc_hd__buf_1 _36420_ (.A(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__buf_1 _36421_ (.A(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__a2bb2o_4 _36422_ (.A1_N(_03254_),
    .A2_N(_05893_),
    .B1(_05886_),
    .B2(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__nand4_4 _36423_ (.A(_05887_),
    .B(_05902_),
    .C(_03437_),
    .D(_03445_),
    .Y(_05913_));
 sky130_fd_sc_hd__buf_1 _36424_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05914_));
 sky130_fd_sc_hd__buf_1 _36425_ (.A(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__buf_1 _36426_ (.A(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__buf_1 _36427_ (.A(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__nand2_4 _36428_ (.A(_05917_),
    .B(_03421_),
    .Y(_05918_));
 sky130_vsdinv _36429_ (.A(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__a21o_4 _36430_ (.A1(_05912_),
    .A2(_05913_),
    .B1(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__nand3_4 _36431_ (.A(_05912_),
    .B(_05913_),
    .C(_05919_),
    .Y(_05921_));
 sky130_fd_sc_hd__nand2_4 _36432_ (.A(_05897_),
    .B(_03455_),
    .Y(_05922_));
 sky130_vsdinv _36433_ (.A(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__a21o_4 _36434_ (.A1(_05920_),
    .A2(_05921_),
    .B1(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__nand3_4 _36435_ (.A(_05920_),
    .B(_05923_),
    .C(_05921_),
    .Y(_05925_));
 sky130_fd_sc_hd__buf_1 _36436_ (.A(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__a21boi_4 _36437_ (.A1(_05894_),
    .A2(_05904_),
    .B1_N(_05898_),
    .Y(_05927_));
 sky130_vsdinv _36438_ (.A(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__a21o_4 _36439_ (.A1(_05924_),
    .A2(_05926_),
    .B1(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__nand3_4 _36440_ (.A(_05924_),
    .B(_05926_),
    .C(_05928_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand2_4 _36441_ (.A(_05929_),
    .B(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__xor2_4 _36442_ (.A(_05908_),
    .B(_05931_),
    .X(_01412_));
 sky130_vsdinv _36443_ (.A(_05908_),
    .Y(_05932_));
 sky130_vsdinv _36444_ (.A(_05930_),
    .Y(_05933_));
 sky130_fd_sc_hd__a21oi_4 _36445_ (.A1(_05929_),
    .A2(_05932_),
    .B1(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__buf_1 _36446_ (.A(_03252_),
    .X(_05935_));
 sky130_fd_sc_hd__buf_1 _36447_ (.A(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__buf_1 _36448_ (.A(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__buf_1 _36449_ (.A(\pcpi_mul.rs2[2] ),
    .X(_05938_));
 sky130_fd_sc_hd__buf_1 _36450_ (.A(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__buf_1 _36451_ (.A(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__nand2_4 _36452_ (.A(_05937_),
    .B(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__buf_1 _36453_ (.A(_05914_),
    .X(_05942_));
 sky130_fd_sc_hd__buf_1 _36454_ (.A(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__buf_1 _36455_ (.A(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__nand2_4 _36456_ (.A(_05944_),
    .B(_03436_),
    .Y(_05945_));
 sky130_fd_sc_hd__nand2_4 _36457_ (.A(_05941_),
    .B(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__buf_1 _36458_ (.A(_03434_),
    .X(_05947_));
 sky130_fd_sc_hd__buf_1 _36459_ (.A(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__nand4_4 _36460_ (.A(_05937_),
    .B(_05917_),
    .C(_05948_),
    .D(_05911_),
    .Y(_05949_));
 sky130_fd_sc_hd__buf_1 _36461_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05950_));
 sky130_fd_sc_hd__buf_1 _36462_ (.A(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__buf_1 _36463_ (.A(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__buf_1 _36464_ (.A(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__buf_1 _36465_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05954_));
 sky130_fd_sc_hd__buf_1 _36466_ (.A(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__buf_1 _36467_ (.A(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__nand2_4 _36468_ (.A(_05953_),
    .B(_05956_),
    .Y(_05957_));
 sky130_vsdinv _36469_ (.A(_05957_),
    .Y(_05958_));
 sky130_fd_sc_hd__a21o_4 _36470_ (.A1(_05946_),
    .A2(_05949_),
    .B1(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__nand3_4 _36471_ (.A(_05946_),
    .B(_05949_),
    .C(_05958_),
    .Y(_05960_));
 sky130_fd_sc_hd__buf_1 _36472_ (.A(_05583_),
    .X(_05961_));
 sky130_fd_sc_hd__buf_1 _36473_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05962_));
 sky130_fd_sc_hd__buf_1 _36474_ (.A(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__nand2_4 _36475_ (.A(_05961_),
    .B(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__buf_1 _36476_ (.A(_05883_),
    .X(_05965_));
 sky130_fd_sc_hd__buf_1 _36477_ (.A(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__buf_1 _36478_ (.A(_03452_),
    .X(_05967_));
 sky130_fd_sc_hd__nand2_4 _36479_ (.A(_05966_),
    .B(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__nor2_4 _36480_ (.A(_05964_),
    .B(_05968_),
    .Y(_05969_));
 sky130_vsdinv _36481_ (.A(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand2_4 _36482_ (.A(_05964_),
    .B(_05968_),
    .Y(_05971_));
 sky130_fd_sc_hd__nand2_4 _36483_ (.A(_05970_),
    .B(_05971_),
    .Y(_05972_));
 sky130_vsdinv _36484_ (.A(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__a21o_4 _36485_ (.A1(_05959_),
    .A2(_05960_),
    .B1(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__nand3_4 _36486_ (.A(_05973_),
    .B(_05959_),
    .C(_05960_),
    .Y(_05975_));
 sky130_fd_sc_hd__nand2_4 _36487_ (.A(_05974_),
    .B(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__or2_4 _36488_ (.A(_05925_),
    .B(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__nand2_4 _36489_ (.A(_05976_),
    .B(_05926_),
    .Y(_05978_));
 sky130_fd_sc_hd__a21boi_4 _36490_ (.A1(_05912_),
    .A2(_05919_),
    .B1_N(_05913_),
    .Y(_05979_));
 sky130_vsdinv _36491_ (.A(_05979_),
    .Y(_05980_));
 sky130_fd_sc_hd__a21o_4 _36492_ (.A1(_05977_),
    .A2(_05978_),
    .B1(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__nand3_4 _36493_ (.A(_05977_),
    .B(_05978_),
    .C(_05980_),
    .Y(_05982_));
 sky130_fd_sc_hd__nand2_4 _36494_ (.A(_05981_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__xor2_4 _36495_ (.A(_05934_),
    .B(_05983_),
    .X(_01413_));
 sky130_fd_sc_hd__nand3_4 _36496_ (.A(_05929_),
    .B(_05932_),
    .C(_05930_),
    .Y(_05984_));
 sky130_fd_sc_hd__or2_4 _36497_ (.A(_05984_),
    .B(_05983_),
    .X(_05985_));
 sky130_vsdinv _36498_ (.A(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__buf_1 _36499_ (.A(_05965_),
    .X(_05987_));
 sky130_fd_sc_hd__nand2_4 _36500_ (.A(_05987_),
    .B(_05963_),
    .Y(_05988_));
 sky130_fd_sc_hd__buf_1 _36501_ (.A(_03471_),
    .X(_05989_));
 sky130_fd_sc_hd__nand2_4 _36502_ (.A(_05961_),
    .B(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2_4 _36503_ (.A(_05988_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__buf_1 _36504_ (.A(_03464_),
    .X(_05992_));
 sky130_fd_sc_hd__nand4_4 _36505_ (.A(_05584_),
    .B(_05966_),
    .C(_05992_),
    .D(_03472_),
    .Y(_05993_));
 sky130_fd_sc_hd__nand2_4 _36506_ (.A(_05991_),
    .B(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__buf_1 _36507_ (.A(_03452_),
    .X(_05995_));
 sky130_fd_sc_hd__nand2_4 _36508_ (.A(_03253_),
    .B(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__nand2_4 _36509_ (.A(_05994_),
    .B(_05996_),
    .Y(_05997_));
 sky130_vsdinv _36510_ (.A(_05996_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand3_4 _36511_ (.A(_05991_),
    .B(_05993_),
    .C(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__nand2_4 _36512_ (.A(_05997_),
    .B(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2_4 _36513_ (.A(_06000_),
    .B(_05970_),
    .Y(_06001_));
 sky130_fd_sc_hd__nand3_4 _36514_ (.A(_05997_),
    .B(_05969_),
    .C(_05999_),
    .Y(_06002_));
 sky130_fd_sc_hd__buf_1 _36515_ (.A(_05909_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2_4 _36516_ (.A(_05916_),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2_4 _36517_ (.A(_05952_),
    .B(_05947_),
    .Y(_06005_));
 sky130_fd_sc_hd__nand2_4 _36518_ (.A(_06004_),
    .B(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__buf_4 _36519_ (.A(_05914_),
    .X(_06007_));
 sky130_fd_sc_hd__buf_4 _36520_ (.A(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__buf_4 _36521_ (.A(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__buf_1 _36522_ (.A(_03261_),
    .X(_06010_));
 sky130_fd_sc_hd__buf_1 _36523_ (.A(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__buf_1 _36524_ (.A(\pcpi_mul.rs2[1] ),
    .X(_06012_));
 sky130_fd_sc_hd__buf_1 _36525_ (.A(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__buf_1 _36526_ (.A(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__buf_1 _36527_ (.A(_03442_),
    .X(_06015_));
 sky130_fd_sc_hd__buf_1 _36528_ (.A(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__nand4_4 _36529_ (.A(_06009_),
    .B(_06011_),
    .C(_06014_),
    .D(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__buf_1 _36530_ (.A(\pcpi_mul.rs1[5] ),
    .X(_06018_));
 sky130_fd_sc_hd__buf_1 _36531_ (.A(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__buf_1 _36532_ (.A(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__buf_1 _36533_ (.A(_05954_),
    .X(_06021_));
 sky130_fd_sc_hd__nand2_4 _36534_ (.A(_06020_),
    .B(_06021_),
    .Y(_06022_));
 sky130_vsdinv _36535_ (.A(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__a21o_4 _36536_ (.A1(_06006_),
    .A2(_06017_),
    .B1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__nand3_4 _36537_ (.A(_06006_),
    .B(_06017_),
    .C(_06023_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2_4 _36538_ (.A(_06024_),
    .B(_06025_),
    .Y(_06026_));
 sky130_vsdinv _36539_ (.A(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__a21o_4 _36540_ (.A1(_06001_),
    .A2(_06002_),
    .B1(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__nand3_4 _36541_ (.A(_06027_),
    .B(_06001_),
    .C(_06002_),
    .Y(_06029_));
 sky130_fd_sc_hd__nand2_4 _36542_ (.A(_06028_),
    .B(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand2_4 _36543_ (.A(_06030_),
    .B(_05975_),
    .Y(_06031_));
 sky130_vsdinv _36544_ (.A(_05975_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand3_4 _36545_ (.A(_06028_),
    .B(_06032_),
    .C(_06029_),
    .Y(_06033_));
 sky130_fd_sc_hd__nand2_4 _36546_ (.A(_06031_),
    .B(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__a21boi_4 _36547_ (.A1(_05946_),
    .A2(_05958_),
    .B1_N(_05949_),
    .Y(_06035_));
 sky130_fd_sc_hd__nand2_4 _36548_ (.A(_06034_),
    .B(_06035_),
    .Y(_06036_));
 sky130_vsdinv _36549_ (.A(_06035_),
    .Y(_06037_));
 sky130_fd_sc_hd__nand3_4 _36550_ (.A(_06031_),
    .B(_06037_),
    .C(_06033_),
    .Y(_06038_));
 sky130_fd_sc_hd__nand2_4 _36551_ (.A(_06036_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__maj3_4 _36552_ (.A(_05926_),
    .B(_05976_),
    .C(_05979_),
    .X(_06040_));
 sky130_fd_sc_hd__nand2_4 _36553_ (.A(_06039_),
    .B(_06040_),
    .Y(_06041_));
 sky130_vsdinv _36554_ (.A(_06040_),
    .Y(_06042_));
 sky130_fd_sc_hd__nand3_4 _36555_ (.A(_06036_),
    .B(_06042_),
    .C(_06038_),
    .Y(_06043_));
 sky130_fd_sc_hd__nand2_4 _36556_ (.A(_06041_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__nand3_4 _36557_ (.A(_05981_),
    .B(_05933_),
    .C(_05982_),
    .Y(_06045_));
 sky130_fd_sc_hd__nand2_4 _36558_ (.A(_06044_),
    .B(_06045_),
    .Y(_06046_));
 sky130_vsdinv _36559_ (.A(_06045_),
    .Y(_06047_));
 sky130_fd_sc_hd__nand3_4 _36560_ (.A(_06047_),
    .B(_06041_),
    .C(_06043_),
    .Y(_06048_));
 sky130_fd_sc_hd__nand3_4 _36561_ (.A(_05986_),
    .B(_06046_),
    .C(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__buf_1 _36562_ (.A(_03248_),
    .X(_06050_));
 sky130_fd_sc_hd__buf_1 _36563_ (.A(\pcpi_mul.rs2[5] ),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _36564_ (.A(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__nand2_4 _36565_ (.A(_06050_),
    .B(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__buf_1 _36566_ (.A(\pcpi_mul.rs1[2] ),
    .X(_06054_));
 sky130_fd_sc_hd__buf_1 _36567_ (.A(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__buf_1 _36568_ (.A(_05962_),
    .X(_06056_));
 sky130_fd_sc_hd__nand2_4 _36569_ (.A(_06055_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__nand2_4 _36570_ (.A(_06053_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__buf_1 _36571_ (.A(_05962_),
    .X(_06059_));
 sky130_fd_sc_hd__nand4_4 _36572_ (.A(_05987_),
    .B(_05900_),
    .C(_06059_),
    .D(_05989_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_4 _36573_ (.A(_06058_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__nand2_4 _36574_ (.A(_05915_),
    .B(_05995_),
    .Y(_06062_));
 sky130_fd_sc_hd__nand2_4 _36575_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_vsdinv _36576_ (.A(_06062_),
    .Y(_06064_));
 sky130_fd_sc_hd__nand3_4 _36577_ (.A(_06058_),
    .B(_06060_),
    .C(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_4 _36578_ (.A(_06063_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__a21boi_4 _36579_ (.A1(_05991_),
    .A2(_05998_),
    .B1_N(_05993_),
    .Y(_06067_));
 sky130_fd_sc_hd__nand2_4 _36580_ (.A(_06066_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__nand2_4 _36581_ (.A(_05999_),
    .B(_05993_),
    .Y(_06069_));
 sky130_fd_sc_hd__nand3_4 _36582_ (.A(_06069_),
    .B(_06063_),
    .C(_06065_),
    .Y(_06070_));
 sky130_fd_sc_hd__nand2_4 _36583_ (.A(_06068_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__buf_1 _36584_ (.A(_05951_),
    .X(_06072_));
 sky130_fd_sc_hd__buf_1 _36585_ (.A(_05938_),
    .X(_06073_));
 sky130_fd_sc_hd__nand2_4 _36586_ (.A(_06072_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__buf_1 _36587_ (.A(_03267_),
    .X(_06075_));
 sky130_fd_sc_hd__buf_1 _36588_ (.A(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__nand2_4 _36589_ (.A(_06076_),
    .B(_03435_),
    .Y(_06077_));
 sky130_fd_sc_hd__nand2_4 _36590_ (.A(_06074_),
    .B(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__buf_1 _36591_ (.A(_03434_),
    .X(_06079_));
 sky130_fd_sc_hd__buf_1 _36592_ (.A(\pcpi_mul.rs2[2] ),
    .X(_06080_));
 sky130_fd_sc_hd__buf_1 _36593_ (.A(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__nand4_4 _36594_ (.A(_05952_),
    .B(_06020_),
    .C(_06079_),
    .D(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__buf_1 _36595_ (.A(\pcpi_mul.rs1[6] ),
    .X(_06083_));
 sky130_fd_sc_hd__buf_1 _36596_ (.A(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__buf_1 _36597_ (.A(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__buf_1 _36598_ (.A(_05954_),
    .X(_06086_));
 sky130_fd_sc_hd__nand2_4 _36599_ (.A(_06085_),
    .B(_06086_),
    .Y(_06087_));
 sky130_vsdinv _36600_ (.A(_06087_),
    .Y(_06088_));
 sky130_fd_sc_hd__a21o_4 _36601_ (.A1(_06078_),
    .A2(_06082_),
    .B1(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__nand3_4 _36602_ (.A(_06078_),
    .B(_06082_),
    .C(_06088_),
    .Y(_06090_));
 sky130_fd_sc_hd__nand2_4 _36603_ (.A(_06089_),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__nand2_4 _36604_ (.A(_06071_),
    .B(_06091_),
    .Y(_06092_));
 sky130_vsdinv _36605_ (.A(_06091_),
    .Y(_06093_));
 sky130_fd_sc_hd__nand3_4 _36606_ (.A(_06093_),
    .B(_06068_),
    .C(_06070_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_4 _36607_ (.A(_06092_),
    .B(_06094_),
    .Y(_06095_));
 sky130_vsdinv _36608_ (.A(_06002_),
    .Y(_06096_));
 sky130_fd_sc_hd__a21oi_4 _36609_ (.A1(_06027_),
    .A2(_06001_),
    .B1(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__nand2_4 _36610_ (.A(_06095_),
    .B(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__a21o_4 _36611_ (.A1(_06027_),
    .A2(_06001_),
    .B1(_06096_),
    .X(_06099_));
 sky130_fd_sc_hd__nand3_4 _36612_ (.A(_06099_),
    .B(_06092_),
    .C(_06094_),
    .Y(_06100_));
 sky130_fd_sc_hd__nand2_4 _36613_ (.A(_06098_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__a21boi_4 _36614_ (.A1(_06006_),
    .A2(_06023_),
    .B1_N(_06017_),
    .Y(_06102_));
 sky130_fd_sc_hd__nand2_4 _36615_ (.A(_06101_),
    .B(_06102_),
    .Y(_06103_));
 sky130_vsdinv _36616_ (.A(_06102_),
    .Y(_06104_));
 sky130_fd_sc_hd__nand3_4 _36617_ (.A(_06098_),
    .B(_06100_),
    .C(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__nand2_4 _36618_ (.A(_06103_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__nand2_4 _36619_ (.A(_05588_),
    .B(_03478_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand2_4 _36620_ (.A(_06106_),
    .B(_06107_),
    .Y(_06108_));
 sky130_vsdinv _36621_ (.A(_06107_),
    .Y(_06109_));
 sky130_fd_sc_hd__nand3_4 _36622_ (.A(_06103_),
    .B(_06109_),
    .C(_06105_),
    .Y(_06110_));
 sky130_fd_sc_hd__nand2_4 _36623_ (.A(_06108_),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__a21boi_4 _36624_ (.A1(_06031_),
    .A2(_06037_),
    .B1_N(_06033_),
    .Y(_06112_));
 sky130_fd_sc_hd__nand2_4 _36625_ (.A(_06111_),
    .B(_06112_),
    .Y(_06113_));
 sky130_vsdinv _36626_ (.A(_06112_),
    .Y(_06114_));
 sky130_fd_sc_hd__nand3_4 _36627_ (.A(_06108_),
    .B(_06110_),
    .C(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__nand2_4 _36628_ (.A(_06113_),
    .B(_06115_),
    .Y(_06116_));
 sky130_vsdinv _36629_ (.A(_06043_),
    .Y(_06117_));
 sky130_fd_sc_hd__a21o_4 _36630_ (.A1(_06047_),
    .A2(_06041_),
    .B1(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__nand2_4 _36631_ (.A(_06116_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__nand4_4 _36632_ (.A(_06043_),
    .B(_06113_),
    .C(_06048_),
    .D(_06115_),
    .Y(_06120_));
 sky130_fd_sc_hd__nand2_4 _36633_ (.A(_06119_),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__xnor2_4 _36634_ (.A(_06049_),
    .B(_06121_),
    .Y(_01469_));
 sky130_vsdinv _36635_ (.A(_06049_),
    .Y(_06122_));
 sky130_fd_sc_hd__nand2_4 _36636_ (.A(_06121_),
    .B(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__or2_4 _36637_ (.A(_06048_),
    .B(_06116_),
    .X(_06124_));
 sky130_fd_sc_hd__nand2_4 _36638_ (.A(_06123_),
    .B(_06124_),
    .Y(_06125_));
 sky130_fd_sc_hd__buf_1 _36639_ (.A(_03252_),
    .X(_06126_));
 sky130_fd_sc_hd__buf_1 _36640_ (.A(_06126_),
    .X(_06127_));
 sky130_fd_sc_hd__buf_1 _36641_ (.A(_03471_),
    .X(_06128_));
 sky130_fd_sc_hd__nand2_4 _36642_ (.A(_06127_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__buf_1 _36643_ (.A(_03464_),
    .X(_06130_));
 sky130_fd_sc_hd__nand2_4 _36644_ (.A(_06008_),
    .B(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__nand2_4 _36645_ (.A(_06129_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__buf_1 _36646_ (.A(_05935_),
    .X(_06133_));
 sky130_fd_sc_hd__buf_1 _36647_ (.A(\pcpi_mul.rs2[4] ),
    .X(_06134_));
 sky130_fd_sc_hd__buf_1 _36648_ (.A(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__buf_1 _36649_ (.A(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__buf_1 _36650_ (.A(_03470_),
    .X(_06137_));
 sky130_fd_sc_hd__buf_1 _36651_ (.A(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__nand4_4 _36652_ (.A(_06133_),
    .B(_05943_),
    .C(_06136_),
    .D(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__nand2_4 _36653_ (.A(_06132_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__buf_1 _36654_ (.A(_05950_),
    .X(_06141_));
 sky130_fd_sc_hd__buf_1 _36655_ (.A(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__buf_1 _36656_ (.A(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__buf_1 _36657_ (.A(_05967_),
    .X(_06144_));
 sky130_fd_sc_hd__nand2_4 _36658_ (.A(_06143_),
    .B(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__nand2_4 _36659_ (.A(_06140_),
    .B(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__nand4_4 _36660_ (.A(_05953_),
    .B(_06132_),
    .C(_06139_),
    .D(_06144_),
    .Y(_06147_));
 sky130_fd_sc_hd__nand2_4 _36661_ (.A(_06146_),
    .B(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__a21boi_4 _36662_ (.A1(_06058_),
    .A2(_06064_),
    .B1_N(_06060_),
    .Y(_06149_));
 sky130_fd_sc_hd__nand2_4 _36663_ (.A(_06148_),
    .B(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__nand2_4 _36664_ (.A(_06065_),
    .B(_06060_),
    .Y(_06151_));
 sky130_fd_sc_hd__nand3_4 _36665_ (.A(_06151_),
    .B(_06146_),
    .C(_06147_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2_4 _36666_ (.A(_06150_),
    .B(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__buf_1 _36667_ (.A(\pcpi_mul.rs1[7] ),
    .X(_06154_));
 sky130_fd_sc_hd__buf_1 _36668_ (.A(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__buf_1 _36669_ (.A(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__nand2_4 _36670_ (.A(_06156_),
    .B(_05956_),
    .Y(_06157_));
 sky130_vsdinv _36671_ (.A(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__buf_1 _36672_ (.A(_03267_),
    .X(_06159_));
 sky130_fd_sc_hd__buf_1 _36673_ (.A(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__buf_1 _36674_ (.A(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__nand2_4 _36675_ (.A(_06161_),
    .B(_06016_),
    .Y(_06162_));
 sky130_fd_sc_hd__buf_1 _36676_ (.A(_03271_),
    .X(_06163_));
 sky130_fd_sc_hd__buf_1 _36677_ (.A(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__buf_1 _36678_ (.A(_06013_),
    .X(_06165_));
 sky130_fd_sc_hd__nand2_4 _36679_ (.A(_06164_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__nand2_4 _36680_ (.A(_06162_),
    .B(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__buf_1 _36681_ (.A(_06076_),
    .X(_06168_));
 sky130_fd_sc_hd__buf_1 _36682_ (.A(_06083_),
    .X(_06169_));
 sky130_fd_sc_hd__buf_1 _36683_ (.A(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__buf_1 _36684_ (.A(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__nand4_4 _36685_ (.A(_06168_),
    .B(_06171_),
    .C(_05948_),
    .D(_05940_),
    .Y(_06172_));
 sky130_fd_sc_hd__nand2_4 _36686_ (.A(_06167_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__xor2_4 _36687_ (.A(_06158_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__nand2_4 _36688_ (.A(_06153_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__xor2_4 _36689_ (.A(_06157_),
    .B(_06173_),
    .X(_06176_));
 sky130_fd_sc_hd__nand3_4 _36690_ (.A(_06176_),
    .B(_06150_),
    .C(_06152_),
    .Y(_06177_));
 sky130_fd_sc_hd__nand2_4 _36691_ (.A(_06175_),
    .B(_06177_),
    .Y(_06178_));
 sky130_vsdinv _36692_ (.A(_06070_),
    .Y(_06179_));
 sky130_fd_sc_hd__a21oi_4 _36693_ (.A1(_06093_),
    .A2(_06068_),
    .B1(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__nand2_4 _36694_ (.A(_06178_),
    .B(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__a21o_4 _36695_ (.A1(_06093_),
    .A2(_06068_),
    .B1(_06179_),
    .X(_06182_));
 sky130_fd_sc_hd__nand3_4 _36696_ (.A(_06182_),
    .B(_06175_),
    .C(_06177_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand2_4 _36697_ (.A(_06181_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__a21boi_4 _36698_ (.A1(_06078_),
    .A2(_06088_),
    .B1_N(_06082_),
    .Y(_06185_));
 sky130_fd_sc_hd__nand2_4 _36699_ (.A(_06184_),
    .B(_06185_),
    .Y(_06186_));
 sky130_vsdinv _36700_ (.A(_06185_),
    .Y(_06187_));
 sky130_fd_sc_hd__nand3_4 _36701_ (.A(_06181_),
    .B(_06183_),
    .C(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__nand2_4 _36702_ (.A(_06186_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_4 _36703_ (.A(_05897_),
    .B(_03483_),
    .Y(_06190_));
 sky130_fd_sc_hd__nand2_4 _36704_ (.A(_05887_),
    .B(_03478_),
    .Y(_06191_));
 sky130_fd_sc_hd__nor2_4 _36705_ (.A(_06190_),
    .B(_06191_),
    .Y(_06192_));
 sky130_vsdinv _36706_ (.A(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__nand2_4 _36707_ (.A(_06190_),
    .B(_06191_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_4 _36708_ (.A(_06193_),
    .B(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__nand2_4 _36709_ (.A(_06189_),
    .B(_06195_),
    .Y(_06196_));
 sky130_vsdinv _36710_ (.A(_06195_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand3_4 _36711_ (.A(_06186_),
    .B(_06197_),
    .C(_06188_),
    .Y(_06198_));
 sky130_fd_sc_hd__nand2_4 _36712_ (.A(_06196_),
    .B(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__nand2_4 _36713_ (.A(_06199_),
    .B(_06110_),
    .Y(_06200_));
 sky130_vsdinv _36714_ (.A(_06110_),
    .Y(_06201_));
 sky130_fd_sc_hd__nand3_4 _36715_ (.A(_06201_),
    .B(_06196_),
    .C(_06198_),
    .Y(_06202_));
 sky130_fd_sc_hd__nand2_4 _36716_ (.A(_06200_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__a21boi_4 _36717_ (.A1(_06098_),
    .A2(_06104_),
    .B1_N(_06100_),
    .Y(_06204_));
 sky130_fd_sc_hd__nand2_4 _36718_ (.A(_06203_),
    .B(_06204_),
    .Y(_06205_));
 sky130_vsdinv _36719_ (.A(_06204_),
    .Y(_06206_));
 sky130_fd_sc_hd__nand3_4 _36720_ (.A(_06200_),
    .B(_06202_),
    .C(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__buf_1 _36721_ (.A(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__nand2_4 _36722_ (.A(_06205_),
    .B(_06208_),
    .Y(_06209_));
 sky130_vsdinv _36723_ (.A(_06115_),
    .Y(_06210_));
 sky130_fd_sc_hd__a21oi_4 _36724_ (.A1(_06113_),
    .A2(_06117_),
    .B1(_06210_),
    .Y(_06211_));
 sky130_vsdinv _36725_ (.A(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_4 _36726_ (.A(_06209_),
    .B(_06212_),
    .Y(_06213_));
 sky130_fd_sc_hd__nand3_4 _36727_ (.A(_06205_),
    .B(_06211_),
    .C(_06208_),
    .Y(_06214_));
 sky130_fd_sc_hd__nand2_4 _36728_ (.A(_06213_),
    .B(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__xnor2_4 _36729_ (.A(_06125_),
    .B(_06215_),
    .Y(_06216_));
 sky130_vsdinv _36730_ (.A(_06216_),
    .Y(_01470_));
 sky130_vsdinv _36731_ (.A(_06207_),
    .Y(_06217_));
 sky130_fd_sc_hd__a21oi_4 _36732_ (.A1(_06205_),
    .A2(_06210_),
    .B1(_06217_),
    .Y(_06218_));
 sky130_vsdinv _36733_ (.A(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__buf_1 _36734_ (.A(_03471_),
    .X(_06220_));
 sky130_fd_sc_hd__nand2_4 _36735_ (.A(_05943_),
    .B(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__buf_1 _36736_ (.A(_05950_),
    .X(_06222_));
 sky130_fd_sc_hd__buf_1 _36737_ (.A(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__nand2_4 _36738_ (.A(_06223_),
    .B(_05992_),
    .Y(_06224_));
 sky130_fd_sc_hd__nand2_4 _36739_ (.A(_06221_),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__buf_1 _36740_ (.A(_05914_),
    .X(_06226_));
 sky130_fd_sc_hd__buf_1 _36741_ (.A(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__buf_1 _36742_ (.A(_06135_),
    .X(_06228_));
 sky130_fd_sc_hd__buf_1 _36743_ (.A(_06137_),
    .X(_06229_));
 sky130_fd_sc_hd__nand4_4 _36744_ (.A(_06227_),
    .B(_06223_),
    .C(_06228_),
    .D(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__buf_1 _36745_ (.A(\pcpi_mul.rs2[3] ),
    .X(_06231_));
 sky130_fd_sc_hd__buf_1 _36746_ (.A(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__nand2_4 _36747_ (.A(_06076_),
    .B(_06232_),
    .Y(_06233_));
 sky130_vsdinv _36748_ (.A(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__a21o_4 _36749_ (.A1(_06225_),
    .A2(_06230_),
    .B1(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__nand3_4 _36750_ (.A(_06225_),
    .B(_06230_),
    .C(_06234_),
    .Y(_06236_));
 sky130_fd_sc_hd__nand2_4 _36751_ (.A(_06235_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__maj3_4 _36752_ (.A(_06129_),
    .B(_06131_),
    .C(_06145_),
    .X(_06238_));
 sky130_fd_sc_hd__nand2_4 _36753_ (.A(_06237_),
    .B(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__nand2_4 _36754_ (.A(_06147_),
    .B(_06139_),
    .Y(_06240_));
 sky130_fd_sc_hd__nand3_4 _36755_ (.A(_06240_),
    .B(_06236_),
    .C(_06235_),
    .Y(_06241_));
 sky130_fd_sc_hd__nand2_4 _36756_ (.A(_06239_),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__buf_1 _36757_ (.A(\pcpi_mul.rs1[6] ),
    .X(_06243_));
 sky130_fd_sc_hd__buf_1 _36758_ (.A(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__buf_1 _36759_ (.A(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__nand2_4 _36760_ (.A(_06245_),
    .B(_06081_),
    .Y(_06246_));
 sky130_fd_sc_hd__buf_1 _36761_ (.A(_03274_),
    .X(_06247_));
 sky130_fd_sc_hd__buf_1 _36762_ (.A(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__nand2_4 _36763_ (.A(_06248_),
    .B(_06079_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand2_4 _36764_ (.A(_06246_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__buf_1 _36765_ (.A(_06154_),
    .X(_06251_));
 sky130_fd_sc_hd__buf_1 _36766_ (.A(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__nand4_4 _36767_ (.A(_06164_),
    .B(_06252_),
    .C(_06014_),
    .D(_06016_),
    .Y(_06253_));
 sky130_fd_sc_hd__buf_1 _36768_ (.A(\pcpi_mul.rs1[8] ),
    .X(_06254_));
 sky130_fd_sc_hd__buf_1 _36769_ (.A(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__buf_1 _36770_ (.A(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__nand2_4 _36771_ (.A(_06256_),
    .B(_06021_),
    .Y(_06257_));
 sky130_vsdinv _36772_ (.A(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__a21o_4 _36773_ (.A1(_06250_),
    .A2(_06253_),
    .B1(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__nand3_4 _36774_ (.A(_06250_),
    .B(_06253_),
    .C(_06258_),
    .Y(_06260_));
 sky130_fd_sc_hd__and2_4 _36775_ (.A(_06259_),
    .B(_06260_),
    .X(_06261_));
 sky130_vsdinv _36776_ (.A(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__nand2_4 _36777_ (.A(_06242_),
    .B(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__nand3_4 _36778_ (.A(_06239_),
    .B(_06241_),
    .C(_06261_),
    .Y(_06264_));
 sky130_fd_sc_hd__nand2_4 _36779_ (.A(_06263_),
    .B(_06264_),
    .Y(_06265_));
 sky130_vsdinv _36780_ (.A(_06152_),
    .Y(_06266_));
 sky130_fd_sc_hd__a21oi_4 _36781_ (.A1(_06176_),
    .A2(_06150_),
    .B1(_06266_),
    .Y(_06267_));
 sky130_fd_sc_hd__nand2_4 _36782_ (.A(_06265_),
    .B(_06267_),
    .Y(_06268_));
 sky130_vsdinv _36783_ (.A(_06267_),
    .Y(_06269_));
 sky130_fd_sc_hd__nand3_4 _36784_ (.A(_06269_),
    .B(_06264_),
    .C(_06263_),
    .Y(_06270_));
 sky130_fd_sc_hd__nand2_4 _36785_ (.A(_06268_),
    .B(_06270_),
    .Y(_06271_));
 sky130_fd_sc_hd__a21boi_4 _36786_ (.A1(_06167_),
    .A2(_06158_),
    .B1_N(_06172_),
    .Y(_06272_));
 sky130_fd_sc_hd__nand2_4 _36787_ (.A(_06271_),
    .B(_06272_),
    .Y(_06273_));
 sky130_vsdinv _36788_ (.A(_06272_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand3_4 _36789_ (.A(_06268_),
    .B(_06270_),
    .C(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__buf_1 _36790_ (.A(_05987_),
    .X(_06276_));
 sky130_fd_sc_hd__buf_8 _36791_ (.A(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__nand2_4 _36792_ (.A(_06277_),
    .B(_03483_),
    .Y(_06278_));
 sky130_fd_sc_hd__nand2_4 _36793_ (.A(_05896_),
    .B(_03493_),
    .Y(_06279_));
 sky130_fd_sc_hd__nand2_4 _36794_ (.A(_06278_),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__nand4_4 _36795_ (.A(_05896_),
    .B(_06277_),
    .C(_03483_),
    .D(_03493_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_4 _36796_ (.A(_05902_),
    .B(_03478_),
    .Y(_06282_));
 sky130_vsdinv _36797_ (.A(_06282_),
    .Y(_06283_));
 sky130_fd_sc_hd__a21o_4 _36798_ (.A1(_06280_),
    .A2(_06281_),
    .B1(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__nand3_4 _36799_ (.A(_06280_),
    .B(_06281_),
    .C(_06283_),
    .Y(_06285_));
 sky130_fd_sc_hd__nand2_4 _36800_ (.A(_06284_),
    .B(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__xor2_4 _36801_ (.A(_06193_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__a21o_4 _36802_ (.A1(_06273_),
    .A2(_06275_),
    .B1(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__nand3_4 _36803_ (.A(_06273_),
    .B(_06287_),
    .C(_06275_),
    .Y(_06289_));
 sky130_vsdinv _36804_ (.A(_06198_),
    .Y(_06290_));
 sky130_fd_sc_hd__a21o_4 _36805_ (.A1(_06288_),
    .A2(_06289_),
    .B1(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__nand3_4 _36806_ (.A(_06288_),
    .B(_06290_),
    .C(_06289_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_4 _36807_ (.A(_06291_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__a21boi_4 _36808_ (.A1(_06181_),
    .A2(_06187_),
    .B1_N(_06183_),
    .Y(_06294_));
 sky130_fd_sc_hd__nand2_4 _36809_ (.A(_06202_),
    .B(_06294_),
    .Y(_06295_));
 sky130_vsdinv _36810_ (.A(_06294_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand4_4 _36811_ (.A(_06201_),
    .B(_06196_),
    .C(_06198_),
    .D(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__nand2_4 _36812_ (.A(_06295_),
    .B(_06297_),
    .Y(_06298_));
 sky130_fd_sc_hd__nand2_4 _36813_ (.A(_06293_),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand4_4 _36814_ (.A(_06291_),
    .B(_06295_),
    .C(_06292_),
    .D(_06297_),
    .Y(_06300_));
 sky130_fd_sc_hd__nand2_4 _36815_ (.A(_06299_),
    .B(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__nand2_4 _36816_ (.A(_06219_),
    .B(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__nand3_4 _36817_ (.A(_06205_),
    .B(_06210_),
    .C(_06208_),
    .Y(_06303_));
 sky130_fd_sc_hd__nand4_4 _36818_ (.A(_06208_),
    .B(_06303_),
    .C(_06300_),
    .D(_06299_),
    .Y(_06304_));
 sky130_fd_sc_hd__nand2_4 _36819_ (.A(_06302_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__nand2_4 _36820_ (.A(_06125_),
    .B(_06215_),
    .Y(_06306_));
 sky130_fd_sc_hd__nand3_4 _36821_ (.A(_06113_),
    .B(_06117_),
    .C(_06115_),
    .Y(_06307_));
 sky130_fd_sc_hd__or2_4 _36822_ (.A(_06307_),
    .B(_06209_),
    .X(_06308_));
 sky130_fd_sc_hd__nand2_4 _36823_ (.A(_06306_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__xor2_4 _36824_ (.A(_06305_),
    .B(_06309_),
    .X(_01471_));
 sky130_fd_sc_hd__nor2_4 _36825_ (.A(_06303_),
    .B(_06301_),
    .Y(_06310_));
 sky130_fd_sc_hd__a21oi_4 _36826_ (.A1(_06309_),
    .A2(_06305_),
    .B1(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__a21boi_4 _36827_ (.A1(_06239_),
    .A2(_06261_),
    .B1_N(_06241_),
    .Y(_06312_));
 sky130_vsdinv _36828_ (.A(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__buf_1 _36829_ (.A(_03470_),
    .X(_06314_));
 sky130_fd_sc_hd__buf_1 _36830_ (.A(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__nand2_4 _36831_ (.A(_05952_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__buf_1 _36832_ (.A(_06075_),
    .X(_06317_));
 sky130_fd_sc_hd__buf_1 _36833_ (.A(_06135_),
    .X(_06318_));
 sky130_fd_sc_hd__nand2_4 _36834_ (.A(_06317_),
    .B(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__nand2_4 _36835_ (.A(_06316_),
    .B(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__buf_1 _36836_ (.A(_06056_),
    .X(_06321_));
 sky130_fd_sc_hd__buf_1 _36837_ (.A(_06051_),
    .X(_06322_));
 sky130_fd_sc_hd__buf_1 _36838_ (.A(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__nand4_4 _36839_ (.A(_06011_),
    .B(_06020_),
    .C(_06321_),
    .D(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__buf_1 _36840_ (.A(_06083_),
    .X(_06325_));
 sky130_fd_sc_hd__buf_1 _36841_ (.A(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__buf_1 _36842_ (.A(_03452_),
    .X(_06327_));
 sky130_fd_sc_hd__buf_1 _36843_ (.A(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__nand2_4 _36844_ (.A(_06326_),
    .B(_06328_),
    .Y(_06329_));
 sky130_vsdinv _36845_ (.A(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__a21o_4 _36846_ (.A1(_06320_),
    .A2(_06324_),
    .B1(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__nand3_4 _36847_ (.A(_06320_),
    .B(_06324_),
    .C(_06330_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_4 _36848_ (.A(_06331_),
    .B(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__a21boi_4 _36849_ (.A1(_06225_),
    .A2(_06234_),
    .B1_N(_06230_),
    .Y(_06334_));
 sky130_fd_sc_hd__nand2_4 _36850_ (.A(_06333_),
    .B(_06334_),
    .Y(_06335_));
 sky130_vsdinv _36851_ (.A(_06334_),
    .Y(_06336_));
 sky130_fd_sc_hd__nand3_4 _36852_ (.A(_06336_),
    .B(_06331_),
    .C(_06332_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_4 _36853_ (.A(_06335_),
    .B(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__buf_1 _36854_ (.A(_03274_),
    .X(_06339_));
 sky130_fd_sc_hd__buf_1 _36855_ (.A(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__nand2_4 _36856_ (.A(_06340_),
    .B(_06073_),
    .Y(_06341_));
 sky130_fd_sc_hd__buf_1 _36857_ (.A(_03279_),
    .X(_06342_));
 sky130_fd_sc_hd__buf_1 _36858_ (.A(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__nand2_4 _36859_ (.A(_06343_),
    .B(_03435_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand2_4 _36860_ (.A(_06341_),
    .B(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__buf_1 _36861_ (.A(_06254_),
    .X(_06346_));
 sky130_fd_sc_hd__buf_1 _36862_ (.A(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__nand4_4 _36863_ (.A(_06248_),
    .B(_06347_),
    .C(_06079_),
    .D(_06081_),
    .Y(_06348_));
 sky130_fd_sc_hd__buf_1 _36864_ (.A(_03289_),
    .X(_06349_));
 sky130_fd_sc_hd__buf_1 _36865_ (.A(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__nand2_4 _36866_ (.A(_06350_),
    .B(_06086_),
    .Y(_06351_));
 sky130_vsdinv _36867_ (.A(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__a21o_4 _36868_ (.A1(_06345_),
    .A2(_06348_),
    .B1(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__nand3_4 _36869_ (.A(_06345_),
    .B(_06348_),
    .C(_06352_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand2_4 _36870_ (.A(_06353_),
    .B(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__nand2_4 _36871_ (.A(_06338_),
    .B(_06355_),
    .Y(_06356_));
 sky130_vsdinv _36872_ (.A(_06355_),
    .Y(_06357_));
 sky130_fd_sc_hd__nand3_4 _36873_ (.A(_06335_),
    .B(_06337_),
    .C(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand3_4 _36874_ (.A(_06313_),
    .B(_06356_),
    .C(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand2_4 _36875_ (.A(_06356_),
    .B(_06358_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2_4 _36876_ (.A(_06360_),
    .B(_06312_),
    .Y(_06361_));
 sky130_fd_sc_hd__nand2_4 _36877_ (.A(_06359_),
    .B(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__a21boi_4 _36878_ (.A1(_06250_),
    .A2(_06258_),
    .B1_N(_06253_),
    .Y(_06363_));
 sky130_fd_sc_hd__nand2_4 _36879_ (.A(_06362_),
    .B(_06363_),
    .Y(_06364_));
 sky130_vsdinv _36880_ (.A(_06363_),
    .Y(_06365_));
 sky130_fd_sc_hd__nand3_4 _36881_ (.A(_06359_),
    .B(_06361_),
    .C(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__nand2_4 _36882_ (.A(_06364_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__nand3_4 _36883_ (.A(_06284_),
    .B(_06192_),
    .C(_06285_),
    .Y(_06368_));
 sky130_vsdinv _36884_ (.A(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__buf_1 _36885_ (.A(_05883_),
    .X(_06370_));
 sky130_fd_sc_hd__buf_1 _36886_ (.A(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__buf_1 _36887_ (.A(_03490_),
    .X(_06372_));
 sky130_fd_sc_hd__buf_1 _36888_ (.A(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__nand2_4 _36889_ (.A(_06371_),
    .B(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__buf_1 _36890_ (.A(\pcpi_mul.rs2[7] ),
    .X(_06375_));
 sky130_fd_sc_hd__buf_1 _36891_ (.A(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__buf_1 _36892_ (.A(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__nand2_4 _36893_ (.A(_05901_),
    .B(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_4 _36894_ (.A(_06374_),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__buf_1 _36895_ (.A(_03252_),
    .X(_06380_));
 sky130_fd_sc_hd__buf_1 _36896_ (.A(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__nand4_4 _36897_ (.A(_06276_),
    .B(_06381_),
    .C(_06377_),
    .D(_06373_),
    .Y(_06382_));
 sky130_fd_sc_hd__buf_1 _36898_ (.A(\pcpi_mul.rs1[3] ),
    .X(_06383_));
 sky130_fd_sc_hd__buf_1 _36899_ (.A(_06383_),
    .X(_06384_));
 sky130_fd_sc_hd__buf_1 _36900_ (.A(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__nand2_4 _36901_ (.A(_06385_),
    .B(_03477_),
    .Y(_06386_));
 sky130_vsdinv _36902_ (.A(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__a21o_4 _36903_ (.A1(_06379_),
    .A2(_06382_),
    .B1(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__nand3_4 _36904_ (.A(_06379_),
    .B(_06382_),
    .C(_06387_),
    .Y(_06389_));
 sky130_fd_sc_hd__a21boi_4 _36905_ (.A1(_06280_),
    .A2(_06283_),
    .B1_N(_06281_),
    .Y(_06390_));
 sky130_fd_sc_hd__a21boi_4 _36906_ (.A1(_06388_),
    .A2(_06389_),
    .B1_N(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__nand2_4 _36907_ (.A(_06388_),
    .B(_06389_),
    .Y(_06392_));
 sky130_fd_sc_hd__nor2_4 _36908_ (.A(_06390_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__nor2_4 _36909_ (.A(_06391_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__xor2_4 _36910_ (.A(_06369_),
    .B(_06394_),
    .X(_06395_));
 sky130_vsdinv _36911_ (.A(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__nand2_4 _36912_ (.A(_06367_),
    .B(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__nand3_4 _36913_ (.A(_06364_),
    .B(_06395_),
    .C(_06366_),
    .Y(_06398_));
 sky130_fd_sc_hd__buf_1 _36914_ (.A(_06398_),
    .X(_06399_));
 sky130_vsdinv _36915_ (.A(_06289_),
    .Y(_06400_));
 sky130_fd_sc_hd__a21o_4 _36916_ (.A1(_06397_),
    .A2(_06399_),
    .B1(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__nand3_4 _36917_ (.A(_06397_),
    .B(_06400_),
    .C(_06399_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand2_4 _36918_ (.A(_06401_),
    .B(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2_4 _36919_ (.A(_05589_),
    .B(_03497_),
    .Y(_06404_));
 sky130_fd_sc_hd__nand2_4 _36920_ (.A(_06403_),
    .B(_06404_),
    .Y(_06405_));
 sky130_vsdinv _36921_ (.A(_06404_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand3_4 _36922_ (.A(_06401_),
    .B(_06406_),
    .C(_06402_),
    .Y(_06407_));
 sky130_fd_sc_hd__nand2_4 _36923_ (.A(_06405_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__a21o_4 _36924_ (.A1(_06270_),
    .A2(_06275_),
    .B1(_06292_),
    .X(_06409_));
 sky130_fd_sc_hd__nand3_4 _36925_ (.A(_06292_),
    .B(_06270_),
    .C(_06275_),
    .Y(_06410_));
 sky130_fd_sc_hd__nand2_4 _36926_ (.A(_06409_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_4 _36927_ (.A(_06408_),
    .B(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__nand4_4 _36928_ (.A(_06407_),
    .B(_06405_),
    .C(_06409_),
    .D(_06410_),
    .Y(_06413_));
 sky130_fd_sc_hd__nand2_4 _36929_ (.A(_06412_),
    .B(_06413_),
    .Y(_06414_));
 sky130_fd_sc_hd__nand2_4 _36930_ (.A(_06300_),
    .B(_06297_),
    .Y(_06415_));
 sky130_vsdinv _36931_ (.A(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__nand2_4 _36932_ (.A(_06414_),
    .B(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__nand3_4 _36933_ (.A(_06412_),
    .B(_06413_),
    .C(_06415_),
    .Y(_06418_));
 sky130_fd_sc_hd__nand3_4 _36934_ (.A(_06299_),
    .B(_06217_),
    .C(_06300_),
    .Y(_06419_));
 sky130_vsdinv _36935_ (.A(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__a21oi_4 _36936_ (.A1(_06417_),
    .A2(_06418_),
    .B1(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__nand3_4 _36937_ (.A(_06417_),
    .B(_06420_),
    .C(_06418_),
    .Y(_06422_));
 sky130_vsdinv _36938_ (.A(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__nor2_4 _36939_ (.A(_06421_),
    .B(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__xnor2_4 _36940_ (.A(_06311_),
    .B(_06424_),
    .Y(_01472_));
 sky130_fd_sc_hd__o21ai_4 _36941_ (.A1(_06421_),
    .A2(_06311_),
    .B1(_06422_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_4 _36942_ (.A(_06020_),
    .B(_06323_),
    .Y(_06426_));
 sky130_fd_sc_hd__buf_1 _36943_ (.A(_06056_),
    .X(_06427_));
 sky130_fd_sc_hd__nand2_4 _36944_ (.A(_06245_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__nand2_4 _36945_ (.A(_06426_),
    .B(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__buf_1 _36946_ (.A(_06059_),
    .X(_06430_));
 sky130_fd_sc_hd__buf_1 _36947_ (.A(_06051_),
    .X(_06431_));
 sky130_fd_sc_hd__buf_1 _36948_ (.A(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__nand4_4 _36949_ (.A(_06161_),
    .B(_06164_),
    .C(_06430_),
    .D(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__nand2_4 _36950_ (.A(_06156_),
    .B(_03454_),
    .Y(_06434_));
 sky130_vsdinv _36951_ (.A(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__a21o_4 _36952_ (.A1(_06429_),
    .A2(_06433_),
    .B1(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__nand3_4 _36953_ (.A(_06429_),
    .B(_06433_),
    .C(_06435_),
    .Y(_06437_));
 sky130_fd_sc_hd__nand2_4 _36954_ (.A(_06436_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__a21boi_4 _36955_ (.A1(_06320_),
    .A2(_06330_),
    .B1_N(_06324_),
    .Y(_06439_));
 sky130_fd_sc_hd__nand2_4 _36956_ (.A(_06438_),
    .B(_06439_),
    .Y(_06440_));
 sky130_vsdinv _36957_ (.A(_06439_),
    .Y(_06441_));
 sky130_fd_sc_hd__nand3_4 _36958_ (.A(_06441_),
    .B(_06437_),
    .C(_06436_),
    .Y(_06442_));
 sky130_fd_sc_hd__nand2_4 _36959_ (.A(_06440_),
    .B(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__buf_1 _36960_ (.A(_06346_),
    .X(_06444_));
 sky130_fd_sc_hd__nand2_4 _36961_ (.A(_06444_),
    .B(_06081_),
    .Y(_06445_));
 sky130_fd_sc_hd__buf_1 _36962_ (.A(_03289_),
    .X(_06446_));
 sky130_fd_sc_hd__buf_1 _36963_ (.A(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__nand2_4 _36964_ (.A(_06447_),
    .B(_06079_),
    .Y(_06448_));
 sky130_fd_sc_hd__nand2_4 _36965_ (.A(_06445_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__buf_1 _36966_ (.A(\pcpi_mul.rs1[9] ),
    .X(_06450_));
 sky130_fd_sc_hd__buf_1 _36967_ (.A(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__buf_1 _36968_ (.A(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__nand4_4 _36969_ (.A(_06256_),
    .B(_06452_),
    .C(_06014_),
    .D(_03444_),
    .Y(_06453_));
 sky130_fd_sc_hd__buf_1 _36970_ (.A(\pcpi_mul.rs1[10] ),
    .X(_06454_));
 sky130_fd_sc_hd__buf_1 _36971_ (.A(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__buf_1 _36972_ (.A(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__nand2_4 _36973_ (.A(_06456_),
    .B(_03420_),
    .Y(_06457_));
 sky130_vsdinv _36974_ (.A(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__a21o_4 _36975_ (.A1(_06449_),
    .A2(_06453_),
    .B1(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__nand3_4 _36976_ (.A(_06449_),
    .B(_06453_),
    .C(_06458_),
    .Y(_06460_));
 sky130_fd_sc_hd__and2_4 _36977_ (.A(_06459_),
    .B(_06460_),
    .X(_06461_));
 sky130_vsdinv _36978_ (.A(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_4 _36979_ (.A(_06443_),
    .B(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__nand3_4 _36980_ (.A(_06440_),
    .B(_06442_),
    .C(_06461_),
    .Y(_06464_));
 sky130_fd_sc_hd__nand2_4 _36981_ (.A(_06463_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__a21boi_4 _36982_ (.A1(_06335_),
    .A2(_06357_),
    .B1_N(_06337_),
    .Y(_06466_));
 sky130_fd_sc_hd__nand2_4 _36983_ (.A(_06465_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__nand2_4 _36984_ (.A(_06358_),
    .B(_06337_),
    .Y(_06468_));
 sky130_fd_sc_hd__nand3_4 _36985_ (.A(_06468_),
    .B(_06464_),
    .C(_06463_),
    .Y(_06469_));
 sky130_fd_sc_hd__nand2_4 _36986_ (.A(_06467_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__a21boi_4 _36987_ (.A1(_06345_),
    .A2(_06352_),
    .B1_N(_06348_),
    .Y(_06471_));
 sky130_fd_sc_hd__nand2_4 _36988_ (.A(_06470_),
    .B(_06471_),
    .Y(_06472_));
 sky130_vsdinv _36989_ (.A(_06471_),
    .Y(_06473_));
 sky130_fd_sc_hd__nand3_4 _36990_ (.A(_06467_),
    .B(_06473_),
    .C(_06469_),
    .Y(_06474_));
 sky130_fd_sc_hd__nand2_4 _36991_ (.A(_06472_),
    .B(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__nand2_4 _36992_ (.A(_05901_),
    .B(_06373_),
    .Y(_06476_));
 sky130_fd_sc_hd__buf_1 _36993_ (.A(_06375_),
    .X(_06477_));
 sky130_fd_sc_hd__buf_1 _36994_ (.A(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__nand2_4 _36995_ (.A(_06385_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__nand2_4 _36996_ (.A(_06476_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__buf_1 _36997_ (.A(\pcpi_mul.rs2[8] ),
    .X(_06481_));
 sky130_fd_sc_hd__buf_1 _36998_ (.A(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__buf_1 _36999_ (.A(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__nand4_4 _37000_ (.A(_05937_),
    .B(_06009_),
    .C(_03482_),
    .D(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__nand2_4 _37001_ (.A(_06143_),
    .B(_03477_),
    .Y(_06485_));
 sky130_vsdinv _37002_ (.A(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__a21o_4 _37003_ (.A1(_06480_),
    .A2(_06484_),
    .B1(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__nand3_4 _37004_ (.A(_06480_),
    .B(_06484_),
    .C(_06486_),
    .Y(_06488_));
 sky130_fd_sc_hd__a21boi_4 _37005_ (.A1(_06379_),
    .A2(_06387_),
    .B1_N(_06382_),
    .Y(_06489_));
 sky130_fd_sc_hd__a21boi_4 _37006_ (.A1(_06487_),
    .A2(_06488_),
    .B1_N(_06489_),
    .Y(_06490_));
 sky130_vsdinv _37007_ (.A(_06489_),
    .Y(_06491_));
 sky130_fd_sc_hd__and3_4 _37008_ (.A(_06491_),
    .B(_06488_),
    .C(_06487_),
    .X(_06492_));
 sky130_fd_sc_hd__buf_1 _37009_ (.A(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__nor2_4 _37010_ (.A(_06490_),
    .B(_06493_),
    .Y(_06494_));
 sky130_vsdinv _37011_ (.A(_06393_),
    .Y(_06495_));
 sky130_fd_sc_hd__o21ai_4 _37012_ (.A1(_06368_),
    .A2(_06391_),
    .B1(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__xor2_4 _37013_ (.A(_06494_),
    .B(_06496_),
    .X(_06497_));
 sky130_vsdinv _37014_ (.A(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_4 _37015_ (.A(_06475_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__nand3_4 _37016_ (.A(_06472_),
    .B(_06497_),
    .C(_06474_),
    .Y(_06500_));
 sky130_fd_sc_hd__nand2_4 _37017_ (.A(_06499_),
    .B(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__nand2_4 _37018_ (.A(_06501_),
    .B(_06399_),
    .Y(_06502_));
 sky130_vsdinv _37019_ (.A(_06398_),
    .Y(_06503_));
 sky130_fd_sc_hd__nand3_4 _37020_ (.A(_06503_),
    .B(_06499_),
    .C(_06500_),
    .Y(_06504_));
 sky130_fd_sc_hd__buf_1 _37021_ (.A(_03499_),
    .X(_06505_));
 sky130_fd_sc_hd__buf_1 _37022_ (.A(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__buf_1 _37023_ (.A(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__nand2_4 _37024_ (.A(_05586_),
    .B(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__nand2_4 _37025_ (.A(_06277_),
    .B(_03497_),
    .Y(_06509_));
 sky130_fd_sc_hd__nor2_4 _37026_ (.A(_06508_),
    .B(_06509_),
    .Y(_06510_));
 sky130_vsdinv _37027_ (.A(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__nand2_4 _37028_ (.A(_06508_),
    .B(_06509_),
    .Y(_06512_));
 sky130_fd_sc_hd__nand2_4 _37029_ (.A(_06511_),
    .B(_06512_),
    .Y(_06513_));
 sky130_vsdinv _37030_ (.A(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__a21oi_4 _37031_ (.A1(_06502_),
    .A2(_06504_),
    .B1(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__nand3_4 _37032_ (.A(_06502_),
    .B(_06514_),
    .C(_06504_),
    .Y(_06516_));
 sky130_vsdinv _37033_ (.A(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__o21ai_4 _37034_ (.A1(_06515_),
    .A2(_06517_),
    .B1(_06407_),
    .Y(_06518_));
 sky130_vsdinv _37035_ (.A(_06407_),
    .Y(_06519_));
 sky130_fd_sc_hd__a21o_4 _37036_ (.A1(_06502_),
    .A2(_06504_),
    .B1(_06514_),
    .X(_06520_));
 sky130_fd_sc_hd__nand3_4 _37037_ (.A(_06519_),
    .B(_06520_),
    .C(_06516_),
    .Y(_06521_));
 sky130_fd_sc_hd__nand2_4 _37038_ (.A(_06518_),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__nand2_4 _37039_ (.A(_06366_),
    .B(_06359_),
    .Y(_06523_));
 sky130_fd_sc_hd__xor2_4 _37040_ (.A(_06523_),
    .B(_06402_),
    .X(_06524_));
 sky130_fd_sc_hd__nand2_4 _37041_ (.A(_06522_),
    .B(_06524_),
    .Y(_06525_));
 sky130_vsdinv _37042_ (.A(_06524_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand3_4 _37043_ (.A(_06518_),
    .B(_06521_),
    .C(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__nand2_4 _37044_ (.A(_06413_),
    .B(_06409_),
    .Y(_06528_));
 sky130_fd_sc_hd__a21oi_4 _37045_ (.A1(_06525_),
    .A2(_06527_),
    .B1(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__nand3_4 _37046_ (.A(_06525_),
    .B(_06527_),
    .C(_06528_),
    .Y(_06530_));
 sky130_vsdinv _37047_ (.A(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__o21ai_4 _37048_ (.A1(_06529_),
    .A2(_06531_),
    .B1(_06418_),
    .Y(_06532_));
 sky130_fd_sc_hd__nand2_4 _37049_ (.A(_06525_),
    .B(_06527_),
    .Y(_06533_));
 sky130_vsdinv _37050_ (.A(_06528_),
    .Y(_06534_));
 sky130_fd_sc_hd__nand2_4 _37051_ (.A(_06533_),
    .B(_06534_),
    .Y(_06535_));
 sky130_vsdinv _37052_ (.A(_06418_),
    .Y(_06536_));
 sky130_fd_sc_hd__nand3_4 _37053_ (.A(_06535_),
    .B(_06536_),
    .C(_06530_),
    .Y(_06537_));
 sky130_fd_sc_hd__nand2_4 _37054_ (.A(_06532_),
    .B(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__xnor2_4 _37055_ (.A(_06425_),
    .B(_06538_),
    .Y(_01415_));
 sky130_vsdinv _37056_ (.A(_06537_),
    .Y(_06539_));
 sky130_fd_sc_hd__a21oi_4 _37057_ (.A1(_06425_),
    .A2(_06532_),
    .B1(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__a21boi_4 _37058_ (.A1(_06440_),
    .A2(_06461_),
    .B1_N(_06442_),
    .Y(_06541_));
 sky130_vsdinv _37059_ (.A(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__nand2_4 _37060_ (.A(_06085_),
    .B(_06220_),
    .Y(_06543_));
 sky130_fd_sc_hd__buf_1 _37061_ (.A(\pcpi_mul.rs1[7] ),
    .X(_06544_));
 sky130_fd_sc_hd__buf_1 _37062_ (.A(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__nand2_4 _37063_ (.A(_06545_),
    .B(_03465_),
    .Y(_06546_));
 sky130_fd_sc_hd__nand2_4 _37064_ (.A(_06543_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand4_4 _37065_ (.A(_06326_),
    .B(_06340_),
    .C(_06136_),
    .D(_06315_),
    .Y(_06548_));
 sky130_fd_sc_hd__buf_1 _37066_ (.A(_03279_),
    .X(_06549_));
 sky130_fd_sc_hd__buf_1 _37067_ (.A(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__buf_1 _37068_ (.A(_06231_),
    .X(_06551_));
 sky130_fd_sc_hd__nand2_4 _37069_ (.A(_06550_),
    .B(_06551_),
    .Y(_06552_));
 sky130_vsdinv _37070_ (.A(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__a21o_4 _37071_ (.A1(_06547_),
    .A2(_06548_),
    .B1(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__nand3_4 _37072_ (.A(_06547_),
    .B(_06548_),
    .C(_06553_),
    .Y(_06555_));
 sky130_fd_sc_hd__nand2_4 _37073_ (.A(_06554_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__a21boi_4 _37074_ (.A1(_06429_),
    .A2(_06435_),
    .B1_N(_06433_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_4 _37075_ (.A(_06556_),
    .B(_06557_),
    .Y(_06558_));
 sky130_vsdinv _37076_ (.A(_06557_),
    .Y(_06559_));
 sky130_fd_sc_hd__nand3_4 _37077_ (.A(_06559_),
    .B(_06555_),
    .C(_06554_),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_4 _37078_ (.A(_06452_),
    .B(_06016_),
    .Y(_06561_));
 sky130_fd_sc_hd__nand2_4 _37079_ (.A(_06456_),
    .B(_06165_),
    .Y(_06562_));
 sky130_fd_sc_hd__nand2_4 _37080_ (.A(_06561_),
    .B(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__buf_1 _37081_ (.A(_03290_),
    .X(_06564_));
 sky130_fd_sc_hd__buf_1 _37082_ (.A(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__buf_1 _37083_ (.A(\pcpi_mul.rs1[10] ),
    .X(_06566_));
 sky130_fd_sc_hd__buf_1 _37084_ (.A(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__buf_1 _37085_ (.A(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__nand4_4 _37086_ (.A(_06565_),
    .B(_06568_),
    .C(_03436_),
    .D(_05940_),
    .Y(_06569_));
 sky130_fd_sc_hd__buf_1 _37087_ (.A(_03297_),
    .X(_06570_));
 sky130_fd_sc_hd__buf_1 _37088_ (.A(_06570_),
    .X(_06571_));
 sky130_fd_sc_hd__buf_1 _37089_ (.A(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__nand2_4 _37090_ (.A(_06572_),
    .B(_03420_),
    .Y(_06573_));
 sky130_vsdinv _37091_ (.A(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__a21o_4 _37092_ (.A1(_06563_),
    .A2(_06569_),
    .B1(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__nand3_4 _37093_ (.A(_06563_),
    .B(_06569_),
    .C(_06574_),
    .Y(_06576_));
 sky130_fd_sc_hd__and2_4 _37094_ (.A(_06575_),
    .B(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__nand3_4 _37095_ (.A(_06558_),
    .B(_06560_),
    .C(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__nand2_4 _37096_ (.A(_06558_),
    .B(_06560_),
    .Y(_06579_));
 sky130_vsdinv _37097_ (.A(_06577_),
    .Y(_06580_));
 sky130_fd_sc_hd__nand2_4 _37098_ (.A(_06579_),
    .B(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__nand3_4 _37099_ (.A(_06542_),
    .B(_06578_),
    .C(_06581_),
    .Y(_06582_));
 sky130_fd_sc_hd__nand2_4 _37100_ (.A(_06581_),
    .B(_06578_),
    .Y(_06583_));
 sky130_fd_sc_hd__nand2_4 _37101_ (.A(_06583_),
    .B(_06541_),
    .Y(_06584_));
 sky130_fd_sc_hd__a21boi_4 _37102_ (.A1(_06449_),
    .A2(_06458_),
    .B1_N(_06453_),
    .Y(_06585_));
 sky130_vsdinv _37103_ (.A(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__a21o_4 _37104_ (.A1(_06582_),
    .A2(_06584_),
    .B1(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__nand3_4 _37105_ (.A(_06582_),
    .B(_06584_),
    .C(_06586_),
    .Y(_06588_));
 sky130_fd_sc_hd__nand2_4 _37106_ (.A(_06587_),
    .B(_06588_),
    .Y(_06589_));
 sky130_vsdinv _37107_ (.A(_06490_),
    .Y(_06590_));
 sky130_fd_sc_hd__a21oi_4 _37108_ (.A1(_06590_),
    .A2(_06393_),
    .B1(_06493_),
    .Y(_06591_));
 sky130_fd_sc_hd__buf_1 _37109_ (.A(\pcpi_mul.rs2[8] ),
    .X(_06592_));
 sky130_fd_sc_hd__buf_1 _37110_ (.A(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__buf_1 _37111_ (.A(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__buf_1 _37112_ (.A(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__nand2_4 _37113_ (.A(_05944_),
    .B(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__buf_1 _37114_ (.A(_06223_),
    .X(_06597_));
 sky130_fd_sc_hd__buf_1 _37115_ (.A(\pcpi_mul.rs2[7] ),
    .X(_06598_));
 sky130_fd_sc_hd__buf_1 _37116_ (.A(_06598_),
    .X(_06599_));
 sky130_fd_sc_hd__buf_1 _37117_ (.A(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__buf_1 _37118_ (.A(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__nand2_4 _37119_ (.A(_06597_),
    .B(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__nand2_4 _37120_ (.A(_06596_),
    .B(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__nand4_4 _37121_ (.A(_05917_),
    .B(_05953_),
    .C(_06601_),
    .D(_03493_),
    .Y(_06604_));
 sky130_fd_sc_hd__buf_1 _37122_ (.A(\pcpi_mul.rs2[6] ),
    .X(_06605_));
 sky130_fd_sc_hd__buf_1 _37123_ (.A(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__buf_1 _37124_ (.A(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__nand2_4 _37125_ (.A(_06168_),
    .B(_06607_),
    .Y(_06608_));
 sky130_vsdinv _37126_ (.A(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__a21o_4 _37127_ (.A1(_06603_),
    .A2(_06604_),
    .B1(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__nand3_4 _37128_ (.A(_06603_),
    .B(_06604_),
    .C(_06609_),
    .Y(_06611_));
 sky130_fd_sc_hd__a21o_4 _37129_ (.A1(_06610_),
    .A2(_06611_),
    .B1(_06510_),
    .X(_06612_));
 sky130_fd_sc_hd__nand3_4 _37130_ (.A(_06610_),
    .B(_06510_),
    .C(_06611_),
    .Y(_06613_));
 sky130_fd_sc_hd__a21boi_4 _37131_ (.A1(_06480_),
    .A2(_06486_),
    .B1_N(_06484_),
    .Y(_06614_));
 sky130_vsdinv _37132_ (.A(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__a21o_4 _37133_ (.A1(_06612_),
    .A2(_06613_),
    .B1(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__nand3_4 _37134_ (.A(_06612_),
    .B(_06615_),
    .C(_06613_),
    .Y(_06617_));
 sky130_fd_sc_hd__nand2_4 _37135_ (.A(_06616_),
    .B(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__xnor2_4 _37136_ (.A(_06591_),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__nand2_4 _37137_ (.A(_06589_),
    .B(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__xor2_4 _37138_ (.A(_06591_),
    .B(_06618_),
    .X(_06621_));
 sky130_fd_sc_hd__nand3_4 _37139_ (.A(_06621_),
    .B(_06588_),
    .C(_06587_),
    .Y(_06622_));
 sky130_fd_sc_hd__nand2_4 _37140_ (.A(_06620_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand3_4 _37141_ (.A(_06494_),
    .B(_06369_),
    .C(_06394_),
    .Y(_06624_));
 sky130_fd_sc_hd__nand2_4 _37142_ (.A(_06500_),
    .B(_06624_),
    .Y(_06625_));
 sky130_vsdinv _37143_ (.A(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__nand2_4 _37144_ (.A(_06623_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__buf_1 _37145_ (.A(_06622_),
    .X(_06628_));
 sky130_fd_sc_hd__nand3_4 _37146_ (.A(_06620_),
    .B(_06625_),
    .C(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__nand2_4 _37147_ (.A(_06627_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__nand2_4 _37148_ (.A(_06381_),
    .B(_03496_),
    .Y(_06631_));
 sky130_fd_sc_hd__buf_1 _37149_ (.A(_06505_),
    .X(_06632_));
 sky130_fd_sc_hd__nand2_4 _37150_ (.A(_06371_),
    .B(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__buf_1 _37151_ (.A(_05583_),
    .X(_06634_));
 sky130_fd_sc_hd__buf_1 _37152_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06635_));
 sky130_fd_sc_hd__buf_1 _37153_ (.A(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__buf_1 _37154_ (.A(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__nand2_4 _37155_ (.A(_06634_),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__xnor2_4 _37156_ (.A(_06633_),
    .B(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__xor2_4 _37157_ (.A(_06631_),
    .B(_06639_),
    .X(_06640_));
 sky130_vsdinv _37158_ (.A(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_4 _37159_ (.A(_06630_),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__nand3_4 _37160_ (.A(_06627_),
    .B(_06640_),
    .C(_06629_),
    .Y(_06643_));
 sky130_fd_sc_hd__nand2_4 _37161_ (.A(_06642_),
    .B(_06643_),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_4 _37162_ (.A(_06644_),
    .B(_06516_),
    .Y(_06645_));
 sky130_fd_sc_hd__nand3_4 _37163_ (.A(_06642_),
    .B(_06517_),
    .C(_06643_),
    .Y(_06646_));
 sky130_fd_sc_hd__nand2_4 _37164_ (.A(_06645_),
    .B(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__nand2_4 _37165_ (.A(_06474_),
    .B(_06469_),
    .Y(_06648_));
 sky130_fd_sc_hd__xor2_4 _37166_ (.A(_06648_),
    .B(_06504_),
    .X(_06649_));
 sky130_fd_sc_hd__nand2_4 _37167_ (.A(_06647_),
    .B(_06649_),
    .Y(_06650_));
 sky130_vsdinv _37168_ (.A(_06649_),
    .Y(_06651_));
 sky130_fd_sc_hd__nand3_4 _37169_ (.A(_06645_),
    .B(_06651_),
    .C(_06646_),
    .Y(_06652_));
 sky130_fd_sc_hd__nand2_4 _37170_ (.A(_06650_),
    .B(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__a21boi_4 _37171_ (.A1(_06518_),
    .A2(_06526_),
    .B1_N(_06521_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_4 _37172_ (.A(_06653_),
    .B(_06654_),
    .Y(_06655_));
 sky130_vsdinv _37173_ (.A(_06654_),
    .Y(_06656_));
 sky130_fd_sc_hd__nand3_4 _37174_ (.A(_06656_),
    .B(_06650_),
    .C(_06652_),
    .Y(_06657_));
 sky130_fd_sc_hd__nand2_4 _37175_ (.A(_06655_),
    .B(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__nand4_4 _37176_ (.A(_06400_),
    .B(_06397_),
    .C(_06399_),
    .D(_06523_),
    .Y(_06659_));
 sky130_fd_sc_hd__nand2_4 _37177_ (.A(_06658_),
    .B(_06659_),
    .Y(_06660_));
 sky130_vsdinv _37178_ (.A(_06659_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand3_4 _37179_ (.A(_06655_),
    .B(_06657_),
    .C(_06661_),
    .Y(_06662_));
 sky130_fd_sc_hd__a21oi_4 _37180_ (.A1(_06660_),
    .A2(_06662_),
    .B1(_06531_),
    .Y(_06663_));
 sky130_fd_sc_hd__nand3_4 _37181_ (.A(_06660_),
    .B(_06531_),
    .C(_06662_),
    .Y(_06664_));
 sky130_vsdinv _37182_ (.A(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__nor2_4 _37183_ (.A(_06663_),
    .B(_06665_),
    .Y(_06666_));
 sky130_fd_sc_hd__xnor2_4 _37184_ (.A(_06540_),
    .B(_06666_),
    .Y(_01416_));
 sky130_fd_sc_hd__o21ai_4 _37185_ (.A1(_06663_),
    .A2(_06540_),
    .B1(_06664_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand2_4 _37186_ (.A(_06597_),
    .B(_06483_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_4 _37187_ (.A(_06161_),
    .B(_03482_),
    .Y(_06669_));
 sky130_fd_sc_hd__nand2_4 _37188_ (.A(_06668_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand4_4 _37189_ (.A(_06597_),
    .B(_06168_),
    .C(_06601_),
    .D(_06595_),
    .Y(_06671_));
 sky130_fd_sc_hd__nand2_4 _37190_ (.A(_06171_),
    .B(_06607_),
    .Y(_06672_));
 sky130_vsdinv _37191_ (.A(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nand3_4 _37192_ (.A(_06670_),
    .B(_06671_),
    .C(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__a21o_4 _37193_ (.A1(_06670_),
    .A2(_06671_),
    .B1(_06673_),
    .X(_06675_));
 sky130_fd_sc_hd__maj3_4 _37194_ (.A(_06631_),
    .B(_06633_),
    .C(_06638_),
    .X(_06676_));
 sky130_vsdinv _37195_ (.A(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__a21o_4 _37196_ (.A1(_06674_),
    .A2(_06675_),
    .B1(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__nand3_4 _37197_ (.A(_06677_),
    .B(_06674_),
    .C(_06675_),
    .Y(_06679_));
 sky130_fd_sc_hd__a21boi_4 _37198_ (.A1(_06603_),
    .A2(_06609_),
    .B1_N(_06604_),
    .Y(_06680_));
 sky130_vsdinv _37199_ (.A(_06680_),
    .Y(_06681_));
 sky130_fd_sc_hd__a21o_4 _37200_ (.A1(_06678_),
    .A2(_06679_),
    .B1(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__nand3_4 _37201_ (.A(_06678_),
    .B(_06681_),
    .C(_06679_),
    .Y(_06683_));
 sky130_fd_sc_hd__a21boi_4 _37202_ (.A1(_06612_),
    .A2(_06615_),
    .B1_N(_06613_),
    .Y(_06684_));
 sky130_vsdinv _37203_ (.A(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__a21o_4 _37204_ (.A1(_06682_),
    .A2(_06683_),
    .B1(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__nand3_4 _37205_ (.A(_06682_),
    .B(_06683_),
    .C(_06685_),
    .Y(_06687_));
 sky130_fd_sc_hd__nand3_4 _37206_ (.A(_06616_),
    .B(_06493_),
    .C(_06617_),
    .Y(_06688_));
 sky130_vsdinv _37207_ (.A(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__a21o_4 _37208_ (.A1(_06686_),
    .A2(_06687_),
    .B1(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__nand3_4 _37209_ (.A(_06686_),
    .B(_06689_),
    .C(_06687_),
    .Y(_06691_));
 sky130_fd_sc_hd__nand2_4 _37210_ (.A(_06690_),
    .B(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__nand2_4 _37211_ (.A(_06340_),
    .B(_06138_),
    .Y(_06693_));
 sky130_fd_sc_hd__nand2_4 _37212_ (.A(_06343_),
    .B(_03465_),
    .Y(_06694_));
 sky130_fd_sc_hd__nand2_4 _37213_ (.A(_06693_),
    .B(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__buf_1 _37214_ (.A(_06052_),
    .X(_06696_));
 sky130_fd_sc_hd__nand4_4 _37215_ (.A(_06252_),
    .B(_06444_),
    .C(_06321_),
    .D(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__nand2_4 _37216_ (.A(_06565_),
    .B(_06144_),
    .Y(_06698_));
 sky130_fd_sc_hd__a21bo_4 _37217_ (.A1(_06695_),
    .A2(_06697_),
    .B1_N(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__nand4_4 _37218_ (.A(_06565_),
    .B(_06695_),
    .C(_06697_),
    .D(_06144_),
    .Y(_06700_));
 sky130_fd_sc_hd__a21boi_4 _37219_ (.A1(_06547_),
    .A2(_06553_),
    .B1_N(_06548_),
    .Y(_06701_));
 sky130_fd_sc_hd__a21boi_4 _37220_ (.A1(_06699_),
    .A2(_06700_),
    .B1_N(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__nand2_4 _37221_ (.A(_06699_),
    .B(_06700_),
    .Y(_06703_));
 sky130_fd_sc_hd__nor2_4 _37222_ (.A(_06701_),
    .B(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__buf_1 _37223_ (.A(_03442_),
    .X(_06705_));
 sky130_fd_sc_hd__buf_1 _37224_ (.A(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__nand2_4 _37225_ (.A(_06568_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__o21ai_4 _37226_ (.A1(_03299_),
    .A2(_05893_),
    .B1(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__nand4_4 _37227_ (.A(_06568_),
    .B(_06572_),
    .C(_05948_),
    .D(_05911_),
    .Y(_06709_));
 sky130_fd_sc_hd__buf_1 _37228_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06710_));
 sky130_fd_sc_hd__buf_1 _37229_ (.A(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__buf_1 _37230_ (.A(_06711_),
    .X(_06712_));
 sky130_fd_sc_hd__buf_1 _37231_ (.A(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__nand2_4 _37232_ (.A(_06713_),
    .B(_05956_),
    .Y(_06714_));
 sky130_vsdinv _37233_ (.A(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__a21o_4 _37234_ (.A1(_06708_),
    .A2(_06709_),
    .B1(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__nand3_4 _37235_ (.A(_06708_),
    .B(_06709_),
    .C(_06715_),
    .Y(_06717_));
 sky130_fd_sc_hd__and2_4 _37236_ (.A(_06716_),
    .B(_06717_),
    .X(_06718_));
 sky130_vsdinv _37237_ (.A(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__o21ai_4 _37238_ (.A1(_06702_),
    .A2(_06704_),
    .B1(_06719_),
    .Y(_06720_));
 sky130_vsdinv _37239_ (.A(_06704_),
    .Y(_06721_));
 sky130_vsdinv _37240_ (.A(_06702_),
    .Y(_06722_));
 sky130_fd_sc_hd__nand3_4 _37241_ (.A(_06721_),
    .B(_06718_),
    .C(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__a21boi_4 _37242_ (.A1(_06558_),
    .A2(_06577_),
    .B1_N(_06560_),
    .Y(_06724_));
 sky130_vsdinv _37243_ (.A(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__a21o_4 _37244_ (.A1(_06720_),
    .A2(_06723_),
    .B1(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__nand3_4 _37245_ (.A(_06725_),
    .B(_06723_),
    .C(_06720_),
    .Y(_06727_));
 sky130_fd_sc_hd__a21boi_4 _37246_ (.A1(_06563_),
    .A2(_06574_),
    .B1_N(_06569_),
    .Y(_06728_));
 sky130_vsdinv _37247_ (.A(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__a21o_4 _37248_ (.A1(_06726_),
    .A2(_06727_),
    .B1(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__nand3_4 _37249_ (.A(_06726_),
    .B(_06729_),
    .C(_06727_),
    .Y(_06731_));
 sky130_fd_sc_hd__nand2_4 _37250_ (.A(_06730_),
    .B(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__nand2_4 _37251_ (.A(_06692_),
    .B(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand4_4 _37252_ (.A(_06731_),
    .B(_06690_),
    .C(_06730_),
    .D(_06691_),
    .Y(_06734_));
 sky130_fd_sc_hd__nand2_4 _37253_ (.A(_06733_),
    .B(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__nand4_4 _37254_ (.A(_06393_),
    .B(_06616_),
    .C(_06494_),
    .D(_06617_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand3_4 _37255_ (.A(_06735_),
    .B(_06628_),
    .C(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand2_4 _37256_ (.A(_06628_),
    .B(_06736_),
    .Y(_06738_));
 sky130_fd_sc_hd__nand3_4 _37257_ (.A(_06733_),
    .B(_06734_),
    .C(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__nand2_4 _37258_ (.A(_06737_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__nand2_4 _37259_ (.A(_05586_),
    .B(_03514_),
    .Y(_06741_));
 sky130_fd_sc_hd__buf_1 _37260_ (.A(_03499_),
    .X(_06742_));
 sky130_fd_sc_hd__buf_1 _37261_ (.A(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__nand2_4 _37262_ (.A(_05936_),
    .B(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__o21ai_4 _37263_ (.A1(_03250_),
    .A2(_03506_),
    .B1(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__buf_1 _37264_ (.A(_05884_),
    .X(_06746_));
 sky130_fd_sc_hd__buf_1 _37265_ (.A(_03504_),
    .X(_06747_));
 sky130_fd_sc_hd__buf_1 _37266_ (.A(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__nand4_4 _37267_ (.A(_06746_),
    .B(_05936_),
    .C(_06743_),
    .D(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__buf_1 _37268_ (.A(\pcpi_mul.rs2[9] ),
    .X(_06750_));
 sky130_fd_sc_hd__buf_1 _37269_ (.A(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__nand2_4 _37270_ (.A(_05943_),
    .B(_06751_),
    .Y(_06752_));
 sky130_vsdinv _37271_ (.A(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__a21o_4 _37272_ (.A1(_06745_),
    .A2(_06749_),
    .B1(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__nand3_4 _37273_ (.A(_06745_),
    .B(_06753_),
    .C(_06749_),
    .Y(_06755_));
 sky130_fd_sc_hd__nand2_4 _37274_ (.A(_06754_),
    .B(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__xor2_4 _37275_ (.A(_06741_),
    .B(_06756_),
    .X(_06757_));
 sky130_vsdinv _37276_ (.A(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__nand2_4 _37277_ (.A(_06740_),
    .B(_06758_),
    .Y(_06759_));
 sky130_fd_sc_hd__nand3_4 _37278_ (.A(_06737_),
    .B(_06757_),
    .C(_06739_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_4 _37279_ (.A(_06759_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_4 _37280_ (.A(_06761_),
    .B(_06643_),
    .Y(_06762_));
 sky130_vsdinv _37281_ (.A(_06643_),
    .Y(_06763_));
 sky130_fd_sc_hd__nand3_4 _37282_ (.A(_06759_),
    .B(_06763_),
    .C(_06760_),
    .Y(_06764_));
 sky130_fd_sc_hd__nand2_4 _37283_ (.A(_06762_),
    .B(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__nand2_4 _37284_ (.A(_06588_),
    .B(_06582_),
    .Y(_06766_));
 sky130_fd_sc_hd__xor2_4 _37285_ (.A(_06766_),
    .B(_06629_),
    .X(_06767_));
 sky130_fd_sc_hd__nand2_4 _37286_ (.A(_06765_),
    .B(_06767_),
    .Y(_06768_));
 sky130_vsdinv _37287_ (.A(_06767_),
    .Y(_06769_));
 sky130_fd_sc_hd__nand3_4 _37288_ (.A(_06762_),
    .B(_06764_),
    .C(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__nand2_4 _37289_ (.A(_06768_),
    .B(_06770_),
    .Y(_06771_));
 sky130_fd_sc_hd__a21boi_4 _37290_ (.A1(_06645_),
    .A2(_06651_),
    .B1_N(_06646_),
    .Y(_06772_));
 sky130_fd_sc_hd__nand2_4 _37291_ (.A(_06771_),
    .B(_06772_),
    .Y(_06773_));
 sky130_vsdinv _37292_ (.A(_06772_),
    .Y(_06774_));
 sky130_fd_sc_hd__nand3_4 _37293_ (.A(_06768_),
    .B(_06770_),
    .C(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__nand2_4 _37294_ (.A(_06773_),
    .B(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__nand4_4 _37295_ (.A(_06503_),
    .B(_06499_),
    .C(_06500_),
    .D(_06648_),
    .Y(_06777_));
 sky130_fd_sc_hd__nand2_4 _37296_ (.A(_06776_),
    .B(_06777_),
    .Y(_06778_));
 sky130_vsdinv _37297_ (.A(_06777_),
    .Y(_06779_));
 sky130_fd_sc_hd__nand3_4 _37298_ (.A(_06773_),
    .B(_06775_),
    .C(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__nand2_4 _37299_ (.A(_06778_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__a21boi_4 _37300_ (.A1(_06655_),
    .A2(_06661_),
    .B1_N(_06657_),
    .Y(_06782_));
 sky130_fd_sc_hd__nand2_4 _37301_ (.A(_06781_),
    .B(_06782_),
    .Y(_06783_));
 sky130_vsdinv _37302_ (.A(_06782_),
    .Y(_06784_));
 sky130_fd_sc_hd__nand3_4 _37303_ (.A(_06778_),
    .B(_06780_),
    .C(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__and2_4 _37304_ (.A(_06783_),
    .B(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__xnor2_4 _37305_ (.A(_06667_),
    .B(_06786_),
    .Y(_06787_));
 sky130_vsdinv _37306_ (.A(_06787_),
    .Y(_01417_));
 sky130_fd_sc_hd__buf_1 _37307_ (.A(_06592_),
    .X(_06788_));
 sky130_fd_sc_hd__buf_1 _37308_ (.A(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__nand2_4 _37309_ (.A(_06317_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__buf_1 _37310_ (.A(_06599_),
    .X(_06791_));
 sky130_fd_sc_hd__nand2_4 _37311_ (.A(_06326_),
    .B(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__nand2_4 _37312_ (.A(_06790_),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__buf_1 _37313_ (.A(_06372_),
    .X(_06794_));
 sky130_fd_sc_hd__nand4_4 _37314_ (.A(_06161_),
    .B(_06164_),
    .C(_06377_),
    .D(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__buf_1 _37315_ (.A(\pcpi_mul.rs2[6] ),
    .X(_06796_));
 sky130_fd_sc_hd__buf_1 _37316_ (.A(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__nand2_4 _37317_ (.A(_06252_),
    .B(_06797_),
    .Y(_06798_));
 sky130_vsdinv _37318_ (.A(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__nand3_4 _37319_ (.A(_06793_),
    .B(_06795_),
    .C(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__a21o_4 _37320_ (.A1(_06793_),
    .A2(_06795_),
    .B1(_06799_),
    .X(_06801_));
 sky130_fd_sc_hd__a21boi_4 _37321_ (.A1(_06745_),
    .A2(_06753_),
    .B1_N(_06749_),
    .Y(_06802_));
 sky130_vsdinv _37322_ (.A(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__a21o_4 _37323_ (.A1(_06800_),
    .A2(_06801_),
    .B1(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__nand3_4 _37324_ (.A(_06803_),
    .B(_06800_),
    .C(_06801_),
    .Y(_06805_));
 sky130_fd_sc_hd__nand2_4 _37325_ (.A(_06804_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__a21boi_4 _37326_ (.A1(_06670_),
    .A2(_06673_),
    .B1_N(_06671_),
    .Y(_06807_));
 sky130_fd_sc_hd__nand2_4 _37327_ (.A(_06806_),
    .B(_06807_),
    .Y(_06808_));
 sky130_vsdinv _37328_ (.A(_06807_),
    .Y(_06809_));
 sky130_fd_sc_hd__nand3_4 _37329_ (.A(_06804_),
    .B(_06809_),
    .C(_06805_),
    .Y(_06810_));
 sky130_fd_sc_hd__nand2_4 _37330_ (.A(_06808_),
    .B(_06810_),
    .Y(_06811_));
 sky130_vsdinv _37331_ (.A(_06741_),
    .Y(_06812_));
 sky130_fd_sc_hd__nand3_4 _37332_ (.A(_06754_),
    .B(_06812_),
    .C(_06755_),
    .Y(_06813_));
 sky130_fd_sc_hd__nand2_4 _37333_ (.A(_06811_),
    .B(_06813_),
    .Y(_06814_));
 sky130_vsdinv _37334_ (.A(_06813_),
    .Y(_06815_));
 sky130_fd_sc_hd__nand3_4 _37335_ (.A(_06808_),
    .B(_06815_),
    .C(_06810_),
    .Y(_06816_));
 sky130_fd_sc_hd__nand2_4 _37336_ (.A(_06814_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__a21boi_4 _37337_ (.A1(_06678_),
    .A2(_06681_),
    .B1_N(_06679_),
    .Y(_06818_));
 sky130_fd_sc_hd__nand2_4 _37338_ (.A(_06817_),
    .B(_06818_),
    .Y(_06819_));
 sky130_vsdinv _37339_ (.A(_06818_),
    .Y(_06820_));
 sky130_fd_sc_hd__nand3_4 _37340_ (.A(_06814_),
    .B(_06820_),
    .C(_06816_),
    .Y(_06821_));
 sky130_fd_sc_hd__nand2_4 _37341_ (.A(_06819_),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__nand2_4 _37342_ (.A(_06822_),
    .B(_06687_),
    .Y(_06823_));
 sky130_vsdinv _37343_ (.A(_06687_),
    .Y(_06824_));
 sky130_fd_sc_hd__nand3_4 _37344_ (.A(_06819_),
    .B(_06824_),
    .C(_06821_),
    .Y(_06825_));
 sky130_fd_sc_hd__nand2_4 _37345_ (.A(_06823_),
    .B(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__maj3_4 _37346_ (.A(_06698_),
    .B(_06693_),
    .C(_06694_),
    .X(_06827_));
 sky130_fd_sc_hd__nand2_4 _37347_ (.A(_06343_),
    .B(_03472_),
    .Y(_06828_));
 sky130_fd_sc_hd__nand2_4 _37348_ (.A(_06564_),
    .B(_05992_),
    .Y(_06829_));
 sky130_fd_sc_hd__nand2_4 _37349_ (.A(_06828_),
    .B(_06829_),
    .Y(_06830_));
 sky130_fd_sc_hd__nand4_4 _37350_ (.A(_06347_),
    .B(_06350_),
    .C(_06136_),
    .D(_06315_),
    .Y(_06831_));
 sky130_fd_sc_hd__buf_1 _37351_ (.A(_03293_),
    .X(_06832_));
 sky130_fd_sc_hd__buf_1 _37352_ (.A(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__nand2_4 _37353_ (.A(_06833_),
    .B(_06551_),
    .Y(_06834_));
 sky130_vsdinv _37354_ (.A(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__a21o_4 _37355_ (.A1(_06830_),
    .A2(_06831_),
    .B1(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__nand3_4 _37356_ (.A(_06830_),
    .B(_06831_),
    .C(_06835_),
    .Y(_06837_));
 sky130_fd_sc_hd__nand2_4 _37357_ (.A(_06836_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_4 _37358_ (.A(_06827_),
    .B(_06838_),
    .Y(_06839_));
 sky130_vsdinv _37359_ (.A(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__nand2_4 _37360_ (.A(_06838_),
    .B(_06827_),
    .Y(_06841_));
 sky130_fd_sc_hd__buf_1 _37361_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06842_));
 sky130_fd_sc_hd__buf_1 _37362_ (.A(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__nand2_4 _37363_ (.A(_06843_),
    .B(_06080_),
    .Y(_06844_));
 sky130_fd_sc_hd__o21ai_4 _37364_ (.A1(_03304_),
    .A2(_05892_),
    .B1(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__buf_1 _37365_ (.A(_03297_),
    .X(_06846_));
 sky130_fd_sc_hd__buf_1 _37366_ (.A(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__buf_1 _37367_ (.A(_06710_),
    .X(_06848_));
 sky130_fd_sc_hd__buf_1 _37368_ (.A(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__nand4_4 _37369_ (.A(_06847_),
    .B(_06849_),
    .C(_06013_),
    .D(_06015_),
    .Y(_06850_));
 sky130_fd_sc_hd__buf_1 _37370_ (.A(_03309_),
    .X(_06851_));
 sky130_fd_sc_hd__buf_1 _37371_ (.A(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__buf_1 _37372_ (.A(\pcpi_mul.rs2[0] ),
    .X(_06853_));
 sky130_fd_sc_hd__nand2_4 _37373_ (.A(_06852_),
    .B(_06853_),
    .Y(_06854_));
 sky130_vsdinv _37374_ (.A(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__a21o_4 _37375_ (.A1(_06845_),
    .A2(_06850_),
    .B1(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__nand3_4 _37376_ (.A(_06845_),
    .B(_06850_),
    .C(_06855_),
    .Y(_06857_));
 sky130_fd_sc_hd__and2_4 _37377_ (.A(_06856_),
    .B(_06857_),
    .X(_06858_));
 sky130_fd_sc_hd__buf_1 _37378_ (.A(_06858_),
    .X(_06859_));
 sky130_fd_sc_hd__a21o_4 _37379_ (.A1(_06840_),
    .A2(_06841_),
    .B1(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__nand3_4 _37380_ (.A(_06840_),
    .B(_06859_),
    .C(_06841_),
    .Y(_06861_));
 sky130_fd_sc_hd__a21oi_4 _37381_ (.A1(_06722_),
    .A2(_06718_),
    .B1(_06704_),
    .Y(_06862_));
 sky130_vsdinv _37382_ (.A(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__a21o_4 _37383_ (.A1(_06860_),
    .A2(_06861_),
    .B1(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__nand3_4 _37384_ (.A(_06863_),
    .B(_06860_),
    .C(_06861_),
    .Y(_06865_));
 sky130_fd_sc_hd__nand2_4 _37385_ (.A(_06864_),
    .B(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__a21boi_4 _37386_ (.A1(_06708_),
    .A2(_06715_),
    .B1_N(_06709_),
    .Y(_06867_));
 sky130_fd_sc_hd__nand2_4 _37387_ (.A(_06866_),
    .B(_06867_),
    .Y(_06868_));
 sky130_vsdinv _37388_ (.A(_06867_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand3_4 _37389_ (.A(_06864_),
    .B(_06865_),
    .C(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__and2_4 _37390_ (.A(_06868_),
    .B(_06870_),
    .X(_06871_));
 sky130_vsdinv _37391_ (.A(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__nand2_4 _37392_ (.A(_06826_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand3_4 _37393_ (.A(_06871_),
    .B(_06823_),
    .C(_06825_),
    .Y(_06874_));
 sky130_fd_sc_hd__nand2_4 _37394_ (.A(_06873_),
    .B(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__nand2_4 _37395_ (.A(_06734_),
    .B(_06691_),
    .Y(_06876_));
 sky130_vsdinv _37396_ (.A(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__nand2_4 _37397_ (.A(_06875_),
    .B(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__nand3_4 _37398_ (.A(_06873_),
    .B(_06876_),
    .C(_06874_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_4 _37399_ (.A(_06878_),
    .B(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__buf_1 _37400_ (.A(_03512_),
    .X(_06881_));
 sky130_vsdinv _37401_ (.A(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__a2bb2o_4 _37402_ (.A1_N(_03250_),
    .A2_N(_06882_),
    .B1(_05897_),
    .B2(_03519_),
    .X(_06883_));
 sky130_fd_sc_hd__nand4_4 _37403_ (.A(_05586_),
    .B(_06277_),
    .C(_03514_),
    .D(_03519_),
    .Y(_06884_));
 sky130_fd_sc_hd__buf_1 _37404_ (.A(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__nand2_4 _37405_ (.A(_06883_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__buf_1 _37406_ (.A(_06742_),
    .X(_06887_));
 sky130_fd_sc_hd__buf_1 _37407_ (.A(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__nand2_4 _37408_ (.A(_06385_),
    .B(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__o21ai_4 _37409_ (.A1(_03254_),
    .A2(_03506_),
    .B1(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__buf_1 _37410_ (.A(_06742_),
    .X(_06891_));
 sky130_fd_sc_hd__buf_1 _37411_ (.A(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__buf_1 _37412_ (.A(_06635_),
    .X(_06893_));
 sky130_fd_sc_hd__buf_1 _37413_ (.A(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__nand4_4 _37414_ (.A(_05937_),
    .B(_06009_),
    .C(_06892_),
    .D(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__buf_1 _37415_ (.A(_06751_),
    .X(_06896_));
 sky130_fd_sc_hd__nand2_4 _37416_ (.A(_06143_),
    .B(_06896_),
    .Y(_06897_));
 sky130_vsdinv _37417_ (.A(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__a21o_4 _37418_ (.A1(_06890_),
    .A2(_06895_),
    .B1(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__nand3_4 _37419_ (.A(_06890_),
    .B(_06895_),
    .C(_06898_),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_4 _37420_ (.A(_06899_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__xor2_4 _37421_ (.A(_06886_),
    .B(_06901_),
    .X(_06902_));
 sky130_vsdinv _37422_ (.A(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand2_4 _37423_ (.A(_06880_),
    .B(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__nand3_4 _37424_ (.A(_06878_),
    .B(_06902_),
    .C(_06879_),
    .Y(_06905_));
 sky130_fd_sc_hd__nand2_4 _37425_ (.A(_06904_),
    .B(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__nand2_4 _37426_ (.A(_06906_),
    .B(_06760_),
    .Y(_06907_));
 sky130_vsdinv _37427_ (.A(_06760_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand3_4 _37428_ (.A(_06904_),
    .B(_06908_),
    .C(_06905_),
    .Y(_06909_));
 sky130_fd_sc_hd__nand2_4 _37429_ (.A(_06907_),
    .B(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__nand2_4 _37430_ (.A(_06731_),
    .B(_06727_),
    .Y(_06911_));
 sky130_fd_sc_hd__xor2_4 _37431_ (.A(_06911_),
    .B(_06739_),
    .X(_06912_));
 sky130_fd_sc_hd__nand2_4 _37432_ (.A(_06910_),
    .B(_06912_),
    .Y(_06913_));
 sky130_vsdinv _37433_ (.A(_06912_),
    .Y(_06914_));
 sky130_fd_sc_hd__nand3_4 _37434_ (.A(_06907_),
    .B(_06909_),
    .C(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__nand2_4 _37435_ (.A(_06913_),
    .B(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__a21boi_4 _37436_ (.A1(_06762_),
    .A2(_06769_),
    .B1_N(_06764_),
    .Y(_06917_));
 sky130_fd_sc_hd__nand2_4 _37437_ (.A(_06916_),
    .B(_06917_),
    .Y(_06918_));
 sky130_vsdinv _37438_ (.A(_06917_),
    .Y(_06919_));
 sky130_fd_sc_hd__nand3_4 _37439_ (.A(_06913_),
    .B(_06919_),
    .C(_06915_),
    .Y(_06920_));
 sky130_fd_sc_hd__nand2_4 _37440_ (.A(_06918_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__and4_4 _37441_ (.A(_06620_),
    .B(_06625_),
    .C(_06628_),
    .D(_06766_),
    .X(_06922_));
 sky130_vsdinv _37442_ (.A(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__nand2_4 _37443_ (.A(_06921_),
    .B(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__nand3_4 _37444_ (.A(_06918_),
    .B(_06922_),
    .C(_06920_),
    .Y(_06925_));
 sky130_fd_sc_hd__nand2_4 _37445_ (.A(_06924_),
    .B(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__a21boi_4 _37446_ (.A1(_06773_),
    .A2(_06779_),
    .B1_N(_06775_),
    .Y(_06927_));
 sky130_fd_sc_hd__nand2_4 _37447_ (.A(_06926_),
    .B(_06927_),
    .Y(_06928_));
 sky130_vsdinv _37448_ (.A(_06927_),
    .Y(_06929_));
 sky130_fd_sc_hd__nand3_4 _37449_ (.A(_06924_),
    .B(_06929_),
    .C(_06925_),
    .Y(_06930_));
 sky130_fd_sc_hd__nand2_4 _37450_ (.A(_06928_),
    .B(_06930_),
    .Y(_06931_));
 sky130_vsdinv _37451_ (.A(_06785_),
    .Y(_06932_));
 sky130_fd_sc_hd__a21oi_4 _37452_ (.A1(_06667_),
    .A2(_06783_),
    .B1(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__xor2_4 _37453_ (.A(_06931_),
    .B(_06933_),
    .X(_01418_));
 sky130_fd_sc_hd__nand2_4 _37454_ (.A(_06870_),
    .B(_06865_),
    .Y(_06934_));
 sky130_fd_sc_hd__xor2_4 _37455_ (.A(_06934_),
    .B(_06879_),
    .X(_06935_));
 sky130_fd_sc_hd__a21boi_4 _37456_ (.A1(_06890_),
    .A2(_06898_),
    .B1_N(_06895_),
    .Y(_06936_));
 sky130_fd_sc_hd__buf_1 _37457_ (.A(\pcpi_mul.rs1[6] ),
    .X(_06937_));
 sky130_fd_sc_hd__buf_1 _37458_ (.A(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__buf_1 _37459_ (.A(_06481_),
    .X(_06939_));
 sky130_fd_sc_hd__nand2_4 _37460_ (.A(_06938_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__buf_1 _37461_ (.A(\pcpi_mul.rs1[7] ),
    .X(_06941_));
 sky130_fd_sc_hd__buf_1 _37462_ (.A(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__nand2_4 _37463_ (.A(_06942_),
    .B(_03481_),
    .Y(_06943_));
 sky130_fd_sc_hd__nand2_4 _37464_ (.A(_06940_),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__buf_1 _37465_ (.A(_06247_),
    .X(_06945_));
 sky130_fd_sc_hd__buf_1 _37466_ (.A(_06598_),
    .X(_06946_));
 sky130_fd_sc_hd__buf_1 _37467_ (.A(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__nand4_4 _37468_ (.A(_06326_),
    .B(_06945_),
    .C(_06947_),
    .D(_06789_),
    .Y(_06948_));
 sky130_fd_sc_hd__buf_1 _37469_ (.A(_06605_),
    .X(_06949_));
 sky130_fd_sc_hd__nand2_4 _37470_ (.A(_06550_),
    .B(_06949_),
    .Y(_06950_));
 sky130_vsdinv _37471_ (.A(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__a21o_4 _37472_ (.A1(_06944_),
    .A2(_06948_),
    .B1(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__nand3_4 _37473_ (.A(_06944_),
    .B(_06948_),
    .C(_06951_),
    .Y(_06953_));
 sky130_fd_sc_hd__nand2_4 _37474_ (.A(_06952_),
    .B(_06953_),
    .Y(_06954_));
 sky130_fd_sc_hd__nor2_4 _37475_ (.A(_06936_),
    .B(_06954_),
    .Y(_06955_));
 sky130_vsdinv _37476_ (.A(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__nand2_4 _37477_ (.A(_06954_),
    .B(_06936_),
    .Y(_06957_));
 sky130_fd_sc_hd__a21boi_4 _37478_ (.A1(_06793_),
    .A2(_06799_),
    .B1_N(_06795_),
    .Y(_06958_));
 sky130_vsdinv _37479_ (.A(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__a21o_4 _37480_ (.A1(_06956_),
    .A2(_06957_),
    .B1(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__nand3_4 _37481_ (.A(_06956_),
    .B(_06959_),
    .C(_06957_),
    .Y(_06961_));
 sky130_fd_sc_hd__nand4_4 _37482_ (.A(_06883_),
    .B(_06899_),
    .C(_06885_),
    .D(_06900_),
    .Y(_06962_));
 sky130_vsdinv _37483_ (.A(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__a21o_4 _37484_ (.A1(_06960_),
    .A2(_06961_),
    .B1(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__nand3_4 _37485_ (.A(_06960_),
    .B(_06963_),
    .C(_06961_),
    .Y(_06965_));
 sky130_fd_sc_hd__a21boi_4 _37486_ (.A1(_06804_),
    .A2(_06809_),
    .B1_N(_06805_),
    .Y(_06966_));
 sky130_vsdinv _37487_ (.A(_06966_),
    .Y(_06967_));
 sky130_fd_sc_hd__a21o_4 _37488_ (.A1(_06964_),
    .A2(_06965_),
    .B1(_06967_),
    .X(_06968_));
 sky130_fd_sc_hd__nand3_4 _37489_ (.A(_06964_),
    .B(_06967_),
    .C(_06965_),
    .Y(_06969_));
 sky130_fd_sc_hd__a21boi_4 _37490_ (.A1(_06814_),
    .A2(_06820_),
    .B1_N(_06816_),
    .Y(_06970_));
 sky130_vsdinv _37491_ (.A(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__a21oi_4 _37492_ (.A1(_06968_),
    .A2(_06969_),
    .B1(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand3_4 _37493_ (.A(_06968_),
    .B(_06971_),
    .C(_06969_),
    .Y(_06973_));
 sky130_vsdinv _37494_ (.A(_06973_),
    .Y(_06974_));
 sky130_fd_sc_hd__a21boi_4 _37495_ (.A1(_06830_),
    .A2(_06835_),
    .B1_N(_06831_),
    .Y(_06975_));
 sky130_fd_sc_hd__nand2_4 _37496_ (.A(_06350_),
    .B(_06138_),
    .Y(_06976_));
 sky130_fd_sc_hd__buf_1 _37497_ (.A(_06832_),
    .X(_06977_));
 sky130_fd_sc_hd__nand2_4 _37498_ (.A(_06977_),
    .B(_06318_),
    .Y(_06978_));
 sky130_fd_sc_hd__nand2_4 _37499_ (.A(_06976_),
    .B(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__buf_1 _37500_ (.A(_06446_),
    .X(_06980_));
 sky130_fd_sc_hd__buf_1 _37501_ (.A(_03294_),
    .X(_06981_));
 sky130_fd_sc_hd__nand4_4 _37502_ (.A(_06980_),
    .B(_06981_),
    .C(_06321_),
    .D(_06323_),
    .Y(_06982_));
 sky130_fd_sc_hd__buf_1 _37503_ (.A(_06843_),
    .X(_06983_));
 sky130_fd_sc_hd__nand2_4 _37504_ (.A(_06983_),
    .B(_06328_),
    .Y(_06984_));
 sky130_vsdinv _37505_ (.A(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__a21o_4 _37506_ (.A1(_06979_),
    .A2(_06982_),
    .B1(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__nand3_4 _37507_ (.A(_06979_),
    .B(_06982_),
    .C(_06985_),
    .Y(_06987_));
 sky130_fd_sc_hd__nand2_4 _37508_ (.A(_06986_),
    .B(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__nor2_4 _37509_ (.A(_06975_),
    .B(_06988_),
    .Y(_06989_));
 sky130_vsdinv _37510_ (.A(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__buf_1 _37511_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06991_));
 sky130_fd_sc_hd__buf_1 _37512_ (.A(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__buf_1 _37513_ (.A(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__nand2_4 _37514_ (.A(_06993_),
    .B(_03421_),
    .Y(_06994_));
 sky130_fd_sc_hd__buf_1 _37515_ (.A(_06848_),
    .X(_06995_));
 sky130_fd_sc_hd__buf_1 _37516_ (.A(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__nand2_4 _37517_ (.A(_06996_),
    .B(_06706_),
    .Y(_06997_));
 sky130_fd_sc_hd__buf_1 _37518_ (.A(_03309_),
    .X(_06998_));
 sky130_fd_sc_hd__buf_1 _37519_ (.A(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__buf_1 _37520_ (.A(_06999_),
    .X(_07000_));
 sky130_fd_sc_hd__buf_1 _37521_ (.A(_06012_),
    .X(_07001_));
 sky130_fd_sc_hd__buf_1 _37522_ (.A(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__nand2_4 _37523_ (.A(_07000_),
    .B(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__nand2_4 _37524_ (.A(_06997_),
    .B(_07003_),
    .Y(_07004_));
 sky130_fd_sc_hd__buf_1 _37525_ (.A(_03310_),
    .X(_07005_));
 sky130_fd_sc_hd__buf_1 _37526_ (.A(_07005_),
    .X(_07006_));
 sky130_fd_sc_hd__nand4_4 _37527_ (.A(_06713_),
    .B(_07006_),
    .C(_06014_),
    .D(_03444_),
    .Y(_07007_));
 sky130_fd_sc_hd__nand2_4 _37528_ (.A(_07004_),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__xor2_4 _37529_ (.A(_06994_),
    .B(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__a21boi_4 _37530_ (.A1(_06986_),
    .A2(_06987_),
    .B1_N(_06975_),
    .Y(_07010_));
 sky130_vsdinv _37531_ (.A(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__nand3_4 _37532_ (.A(_06990_),
    .B(_07009_),
    .C(_07011_),
    .Y(_07012_));
 sky130_vsdinv _37533_ (.A(_07009_),
    .Y(_07013_));
 sky130_fd_sc_hd__o21ai_4 _37534_ (.A1(_07010_),
    .A2(_06989_),
    .B1(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__a21oi_4 _37535_ (.A1(_06859_),
    .A2(_06841_),
    .B1(_06839_),
    .Y(_07015_));
 sky130_vsdinv _37536_ (.A(_07015_),
    .Y(_07016_));
 sky130_fd_sc_hd__a21o_4 _37537_ (.A1(_07012_),
    .A2(_07014_),
    .B1(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__nand3_4 _37538_ (.A(_07016_),
    .B(_07012_),
    .C(_07014_),
    .Y(_07018_));
 sky130_fd_sc_hd__a21boi_4 _37539_ (.A1(_06845_),
    .A2(_06855_),
    .B1_N(_06850_),
    .Y(_07019_));
 sky130_vsdinv _37540_ (.A(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__a21oi_4 _37541_ (.A1(_07017_),
    .A2(_07018_),
    .B1(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__nand3_4 _37542_ (.A(_07017_),
    .B(_07020_),
    .C(_07018_),
    .Y(_07022_));
 sky130_vsdinv _37543_ (.A(_07022_),
    .Y(_07023_));
 sky130_fd_sc_hd__nor2_4 _37544_ (.A(_07021_),
    .B(_07023_),
    .Y(_07024_));
 sky130_vsdinv _37545_ (.A(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__o21ai_4 _37546_ (.A1(_06972_),
    .A2(_06974_),
    .B1(_07025_),
    .Y(_07026_));
 sky130_vsdinv _37547_ (.A(_06972_),
    .Y(_07027_));
 sky130_fd_sc_hd__nand3_4 _37548_ (.A(_07027_),
    .B(_07024_),
    .C(_06973_),
    .Y(_07028_));
 sky130_fd_sc_hd__nand2_4 _37549_ (.A(_07026_),
    .B(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__a21boi_4 _37550_ (.A1(_06871_),
    .A2(_06823_),
    .B1_N(_06825_),
    .Y(_07030_));
 sky130_fd_sc_hd__nand2_4 _37551_ (.A(_07029_),
    .B(_07030_),
    .Y(_07031_));
 sky130_vsdinv _37552_ (.A(_07030_),
    .Y(_07032_));
 sky130_fd_sc_hd__nand3_4 _37553_ (.A(_07026_),
    .B(_07032_),
    .C(_07028_),
    .Y(_07033_));
 sky130_fd_sc_hd__nand2_4 _37554_ (.A(_06168_),
    .B(_06896_),
    .Y(_07034_));
 sky130_fd_sc_hd__nand2_4 _37555_ (.A(_06009_),
    .B(_06894_),
    .Y(_07035_));
 sky130_fd_sc_hd__nand2_4 _37556_ (.A(_06143_),
    .B(_06888_),
    .Y(_07036_));
 sky130_fd_sc_hd__nand2_4 _37557_ (.A(_07035_),
    .B(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__buf_1 _37558_ (.A(_06637_),
    .X(_07038_));
 sky130_fd_sc_hd__nand4_4 _37559_ (.A(_05917_),
    .B(_06597_),
    .C(_06507_),
    .D(_07038_),
    .Y(_07039_));
 sky130_fd_sc_hd__nand2_4 _37560_ (.A(_07037_),
    .B(_07039_),
    .Y(_07040_));
 sky130_fd_sc_hd__xor2_4 _37561_ (.A(_07034_),
    .B(_07040_),
    .X(_07041_));
 sky130_vsdinv _37562_ (.A(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__buf_1 _37563_ (.A(\pcpi_mul.rs2[12] ),
    .X(_07043_));
 sky130_fd_sc_hd__buf_1 _37564_ (.A(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__buf_1 _37565_ (.A(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__nand2_4 _37566_ (.A(_06127_),
    .B(_07045_),
    .Y(_07046_));
 sky130_vsdinv _37567_ (.A(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__buf_1 _37568_ (.A(_05884_),
    .X(_07048_));
 sky130_fd_sc_hd__buf_1 _37569_ (.A(\pcpi_mul.rs2[13] ),
    .X(_07049_));
 sky130_fd_sc_hd__buf_1 _37570_ (.A(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__buf_1 _37571_ (.A(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__nand2_4 _37572_ (.A(_07048_),
    .B(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__buf_1 _37573_ (.A(\pcpi_mul.rs2[14] ),
    .X(_07053_));
 sky130_fd_sc_hd__buf_1 _37574_ (.A(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__buf_1 _37575_ (.A(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__nand2_4 _37576_ (.A(_05584_),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand2_4 _37577_ (.A(_07052_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__buf_1 _37578_ (.A(_07049_),
    .X(_07058_));
 sky130_fd_sc_hd__buf_1 _37579_ (.A(_07058_),
    .X(_07059_));
 sky130_fd_sc_hd__nand4_4 _37580_ (.A(_06634_),
    .B(_05885_),
    .C(_07059_),
    .D(_07055_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_4 _37581_ (.A(_07057_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__xor2_4 _37582_ (.A(_07047_),
    .B(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__xnor2_4 _37583_ (.A(_06885_),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__xor2_4 _37584_ (.A(_07042_),
    .B(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__a21o_4 _37585_ (.A1(_07031_),
    .A2(_07033_),
    .B1(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__nand3_4 _37586_ (.A(_07031_),
    .B(_07064_),
    .C(_07033_),
    .Y(_07066_));
 sky130_vsdinv _37587_ (.A(_06905_),
    .Y(_07067_));
 sky130_fd_sc_hd__a21oi_4 _37588_ (.A1(_07065_),
    .A2(_07066_),
    .B1(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__nand3_4 _37589_ (.A(_07065_),
    .B(_07067_),
    .C(_07066_),
    .Y(_07069_));
 sky130_vsdinv _37590_ (.A(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__or3_4 _37591_ (.A(_06935_),
    .B(_07068_),
    .C(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__o21ai_4 _37592_ (.A1(_07068_),
    .A2(_07070_),
    .B1(_06935_),
    .Y(_07072_));
 sky130_fd_sc_hd__a21boi_4 _37593_ (.A1(_06907_),
    .A2(_06914_),
    .B1_N(_06909_),
    .Y(_07073_));
 sky130_vsdinv _37594_ (.A(_07073_),
    .Y(_07074_));
 sky130_fd_sc_hd__a21o_4 _37595_ (.A1(_07071_),
    .A2(_07072_),
    .B1(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__nand3_4 _37596_ (.A(_07071_),
    .B(_07072_),
    .C(_07074_),
    .Y(_07076_));
 sky130_fd_sc_hd__nand2_4 _37597_ (.A(_07075_),
    .B(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__nand4_4 _37598_ (.A(_06734_),
    .B(_06733_),
    .C(_06738_),
    .D(_06911_),
    .Y(_07078_));
 sky130_fd_sc_hd__nand2_4 _37599_ (.A(_07077_),
    .B(_07078_),
    .Y(_07079_));
 sky130_vsdinv _37600_ (.A(_07078_),
    .Y(_07080_));
 sky130_fd_sc_hd__nand3_4 _37601_ (.A(_07075_),
    .B(_07080_),
    .C(_07076_),
    .Y(_07081_));
 sky130_fd_sc_hd__nand2_4 _37602_ (.A(_07079_),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__a21boi_4 _37603_ (.A1(_06918_),
    .A2(_06922_),
    .B1_N(_06920_),
    .Y(_07083_));
 sky130_fd_sc_hd__nand2_4 _37604_ (.A(_07082_),
    .B(_07083_),
    .Y(_07084_));
 sky130_vsdinv _37605_ (.A(_07083_),
    .Y(_07085_));
 sky130_fd_sc_hd__nand3_4 _37606_ (.A(_07079_),
    .B(_07081_),
    .C(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__nand2_4 _37607_ (.A(_07084_),
    .B(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__o21ai_4 _37608_ (.A1(_06931_),
    .A2(_06933_),
    .B1(_06930_),
    .Y(_07088_));
 sky130_fd_sc_hd__xnor2_4 _37609_ (.A(_07087_),
    .B(_07088_),
    .Y(_01419_));
 sky130_fd_sc_hd__and4_4 _37610_ (.A(_06873_),
    .B(_06876_),
    .C(_06874_),
    .D(_06934_),
    .X(_07089_));
 sky130_fd_sc_hd__o21ai_4 _37611_ (.A1(_06935_),
    .A2(_07068_),
    .B1(_07069_),
    .Y(_07090_));
 sky130_fd_sc_hd__maj3_4 _37612_ (.A(_07034_),
    .B(_07035_),
    .C(_07036_),
    .X(_07091_));
 sky130_fd_sc_hd__nand2_4 _37613_ (.A(_06248_),
    .B(_03492_),
    .Y(_07092_));
 sky130_fd_sc_hd__nand2_4 _37614_ (.A(_06347_),
    .B(_06947_),
    .Y(_07093_));
 sky130_fd_sc_hd__nand2_4 _37615_ (.A(_07092_),
    .B(_07093_),
    .Y(_07094_));
 sky130_fd_sc_hd__buf_1 _37616_ (.A(\pcpi_mul.rs2[7] ),
    .X(_07095_));
 sky130_fd_sc_hd__buf_1 _37617_ (.A(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__buf_1 _37618_ (.A(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__nand4_4 _37619_ (.A(_06156_),
    .B(_06256_),
    .C(_07097_),
    .D(_06483_),
    .Y(_07098_));
 sky130_fd_sc_hd__nand2_4 _37620_ (.A(_06980_),
    .B(_03477_),
    .Y(_07099_));
 sky130_vsdinv _37621_ (.A(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__a21o_4 _37622_ (.A1(_07094_),
    .A2(_07098_),
    .B1(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__nand3_4 _37623_ (.A(_07094_),
    .B(_07098_),
    .C(_07100_),
    .Y(_07102_));
 sky130_fd_sc_hd__nand2_4 _37624_ (.A(_07101_),
    .B(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__or2_4 _37625_ (.A(_07091_),
    .B(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__nand2_4 _37626_ (.A(_07103_),
    .B(_07091_),
    .Y(_07105_));
 sky130_fd_sc_hd__a21boi_4 _37627_ (.A1(_06944_),
    .A2(_06951_),
    .B1_N(_06948_),
    .Y(_07106_));
 sky130_vsdinv _37628_ (.A(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__a21o_4 _37629_ (.A1(_07104_),
    .A2(_07105_),
    .B1(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__nand3_4 _37630_ (.A(_07104_),
    .B(_07107_),
    .C(_07105_),
    .Y(_07109_));
 sky130_fd_sc_hd__nand2_4 _37631_ (.A(_07108_),
    .B(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__and2_4 _37632_ (.A(_07062_),
    .B(_06884_),
    .X(_07111_));
 sky130_fd_sc_hd__or2_4 _37633_ (.A(_06885_),
    .B(_07062_),
    .X(_07112_));
 sky130_fd_sc_hd__o21ai_4 _37634_ (.A1(_07042_),
    .A2(_07111_),
    .B1(_07112_),
    .Y(_07113_));
 sky130_vsdinv _37635_ (.A(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__nand2_4 _37636_ (.A(_07110_),
    .B(_07114_),
    .Y(_07115_));
 sky130_fd_sc_hd__nand3_4 _37637_ (.A(_07113_),
    .B(_07108_),
    .C(_07109_),
    .Y(_07116_));
 sky130_fd_sc_hd__a21oi_4 _37638_ (.A1(_06957_),
    .A2(_06959_),
    .B1(_06955_),
    .Y(_07117_));
 sky130_vsdinv _37639_ (.A(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__a21o_4 _37640_ (.A1(_07115_),
    .A2(_07116_),
    .B1(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__nand3_4 _37641_ (.A(_07115_),
    .B(_07118_),
    .C(_07116_),
    .Y(_07120_));
 sky130_fd_sc_hd__nand2_4 _37642_ (.A(_07119_),
    .B(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__a21boi_4 _37643_ (.A1(_06964_),
    .A2(_06967_),
    .B1_N(_06965_),
    .Y(_07122_));
 sky130_fd_sc_hd__nand2_4 _37644_ (.A(_07121_),
    .B(_07122_),
    .Y(_07123_));
 sky130_vsdinv _37645_ (.A(_07122_),
    .Y(_07124_));
 sky130_fd_sc_hd__nand3_4 _37646_ (.A(_07124_),
    .B(_07119_),
    .C(_07120_),
    .Y(_07125_));
 sky130_fd_sc_hd__nand2_4 _37647_ (.A(_07123_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__a21boi_4 _37648_ (.A1(_06979_),
    .A2(_06985_),
    .B1_N(_06982_),
    .Y(_07127_));
 sky130_fd_sc_hd__buf_1 _37649_ (.A(_06314_),
    .X(_07128_));
 sky130_fd_sc_hd__nand2_4 _37650_ (.A(_06981_),
    .B(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__buf_1 _37651_ (.A(_03298_),
    .X(_07130_));
 sky130_fd_sc_hd__buf_1 _37652_ (.A(_06134_),
    .X(_07131_));
 sky130_fd_sc_hd__buf_1 _37653_ (.A(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__nand2_4 _37654_ (.A(_07130_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_4 _37655_ (.A(_07129_),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__nand4_4 _37656_ (.A(_06568_),
    .B(_06572_),
    .C(_06430_),
    .D(_06432_),
    .Y(_07135_));
 sky130_fd_sc_hd__nand2_4 _37657_ (.A(_06996_),
    .B(_03454_),
    .Y(_07136_));
 sky130_fd_sc_hd__a21bo_4 _37658_ (.A1(_07134_),
    .A2(_07135_),
    .B1_N(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__nand4_4 _37659_ (.A(_06713_),
    .B(_07134_),
    .C(_07135_),
    .D(_03455_),
    .Y(_07138_));
 sky130_fd_sc_hd__nand2_4 _37660_ (.A(_07137_),
    .B(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__nor2_4 _37661_ (.A(_07127_),
    .B(_07139_),
    .Y(_07140_));
 sky130_vsdinv _37662_ (.A(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__a21boi_4 _37663_ (.A1(_07137_),
    .A2(_07138_),
    .B1_N(_07127_),
    .Y(_07142_));
 sky130_vsdinv _37664_ (.A(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__buf_1 _37665_ (.A(_05891_),
    .X(_07144_));
 sky130_fd_sc_hd__buf_1 _37666_ (.A(\pcpi_mul.rs1[13] ),
    .X(_07145_));
 sky130_fd_sc_hd__buf_1 _37667_ (.A(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__buf_1 _37668_ (.A(_07146_),
    .X(_07147_));
 sky130_fd_sc_hd__nand2_4 _37669_ (.A(_07147_),
    .B(_06073_),
    .Y(_07148_));
 sky130_fd_sc_hd__o21ai_4 _37670_ (.A1(_03315_),
    .A2(_07144_),
    .B1(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__buf_1 _37671_ (.A(_06851_),
    .X(_07150_));
 sky130_fd_sc_hd__buf_1 _37672_ (.A(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__buf_1 _37673_ (.A(_03313_),
    .X(_07152_));
 sky130_fd_sc_hd__buf_1 _37674_ (.A(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__buf_1 _37675_ (.A(_06705_),
    .X(_07154_));
 sky130_fd_sc_hd__nand4_4 _37676_ (.A(_07151_),
    .B(_07153_),
    .C(_07002_),
    .D(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__buf_1 _37677_ (.A(\pcpi_mul.rs1[15] ),
    .X(_07156_));
 sky130_fd_sc_hd__buf_1 _37678_ (.A(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__buf_1 _37679_ (.A(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__nand2_4 _37680_ (.A(_07158_),
    .B(_06021_),
    .Y(_07159_));
 sky130_vsdinv _37681_ (.A(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__a21o_4 _37682_ (.A1(_07149_),
    .A2(_07155_),
    .B1(_07160_),
    .X(_07161_));
 sky130_fd_sc_hd__nand3_4 _37683_ (.A(_07149_),
    .B(_07155_),
    .C(_07160_),
    .Y(_07162_));
 sky130_fd_sc_hd__and2_4 _37684_ (.A(_07161_),
    .B(_07162_),
    .X(_07163_));
 sky130_fd_sc_hd__buf_1 _37685_ (.A(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__a21o_4 _37686_ (.A1(_07141_),
    .A2(_07143_),
    .B1(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__nand3_4 _37687_ (.A(_07141_),
    .B(_07164_),
    .C(_07143_),
    .Y(_07166_));
 sky130_fd_sc_hd__a21oi_4 _37688_ (.A1(_07011_),
    .A2(_07009_),
    .B1(_06989_),
    .Y(_07167_));
 sky130_vsdinv _37689_ (.A(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__a21o_4 _37690_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07168_),
    .X(_07169_));
 sky130_fd_sc_hd__nand3_4 _37691_ (.A(_07165_),
    .B(_07168_),
    .C(_07166_),
    .Y(_07170_));
 sky130_fd_sc_hd__maj3_4 _37692_ (.A(_06997_),
    .B(_07003_),
    .C(_06994_),
    .X(_07171_));
 sky130_vsdinv _37693_ (.A(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__a21oi_4 _37694_ (.A1(_07169_),
    .A2(_07170_),
    .B1(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__nand3_4 _37695_ (.A(_07169_),
    .B(_07172_),
    .C(_07170_),
    .Y(_07174_));
 sky130_vsdinv _37696_ (.A(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__nor2_4 _37697_ (.A(_07173_),
    .B(_07175_),
    .Y(_07176_));
 sky130_vsdinv _37698_ (.A(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__nand2_4 _37699_ (.A(_07126_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand3_4 _37700_ (.A(_07123_),
    .B(_07125_),
    .C(_07176_),
    .Y(_07179_));
 sky130_fd_sc_hd__nand2_4 _37701_ (.A(_07178_),
    .B(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__o21ai_4 _37702_ (.A1(_07025_),
    .A2(_06972_),
    .B1(_06973_),
    .Y(_07181_));
 sky130_vsdinv _37703_ (.A(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__nand2_4 _37704_ (.A(_07180_),
    .B(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__nand3_4 _37705_ (.A(_07181_),
    .B(_07178_),
    .C(_07179_),
    .Y(_07184_));
 sky130_fd_sc_hd__nand2_4 _37706_ (.A(_07183_),
    .B(_07184_),
    .Y(_07185_));
 sky130_fd_sc_hd__nand2_4 _37707_ (.A(_05588_),
    .B(_03532_),
    .Y(_07186_));
 sky130_fd_sc_hd__buf_1 _37708_ (.A(_07054_),
    .X(_07187_));
 sky130_fd_sc_hd__nand2_4 _37709_ (.A(_05966_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__buf_1 _37710_ (.A(_07058_),
    .X(_07189_));
 sky130_fd_sc_hd__nand2_4 _37711_ (.A(_06127_),
    .B(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__nand2_4 _37712_ (.A(_07188_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__buf_1 _37713_ (.A(_07050_),
    .X(_07192_));
 sky130_fd_sc_hd__buf_1 _37714_ (.A(_07053_),
    .X(_07193_));
 sky130_fd_sc_hd__buf_1 _37715_ (.A(_07193_),
    .X(_07194_));
 sky130_fd_sc_hd__nand4_4 _37716_ (.A(_06371_),
    .B(_06133_),
    .C(_07192_),
    .D(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__buf_1 _37717_ (.A(_06007_),
    .X(_07196_));
 sky130_fd_sc_hd__buf_1 _37718_ (.A(_07044_),
    .X(_07197_));
 sky130_fd_sc_hd__nand2_4 _37719_ (.A(_07196_),
    .B(_07197_),
    .Y(_07198_));
 sky130_vsdinv _37720_ (.A(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__a21o_4 _37721_ (.A1(_07191_),
    .A2(_07195_),
    .B1(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__nand3_4 _37722_ (.A(_07191_),
    .B(_07195_),
    .C(_07199_),
    .Y(_07201_));
 sky130_fd_sc_hd__a21boi_4 _37723_ (.A1(_07057_),
    .A2(_07047_),
    .B1_N(_07060_),
    .Y(_07202_));
 sky130_fd_sc_hd__a21boi_4 _37724_ (.A1(_07200_),
    .A2(_07201_),
    .B1_N(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__buf_1 _37725_ (.A(\pcpi_mul.rs2[9] ),
    .X(_07204_));
 sky130_fd_sc_hd__buf_1 _37726_ (.A(_07204_),
    .X(_07205_));
 sky130_fd_sc_hd__nand2_4 _37727_ (.A(_06085_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand2_4 _37728_ (.A(_06072_),
    .B(_06748_),
    .Y(_07207_));
 sky130_fd_sc_hd__buf_1 _37729_ (.A(_06075_),
    .X(_07208_));
 sky130_fd_sc_hd__nand2_4 _37730_ (.A(_07208_),
    .B(_03501_),
    .Y(_07209_));
 sky130_fd_sc_hd__nand2_4 _37731_ (.A(_07207_),
    .B(_07209_),
    .Y(_07210_));
 sky130_fd_sc_hd__buf_1 _37732_ (.A(\pcpi_mul.rs2[10] ),
    .X(_07211_));
 sky130_fd_sc_hd__buf_1 _37733_ (.A(_07211_),
    .X(_07212_));
 sky130_fd_sc_hd__buf_1 _37734_ (.A(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__buf_1 _37735_ (.A(_06635_),
    .X(_07214_));
 sky130_fd_sc_hd__buf_1 _37736_ (.A(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__nand4_4 _37737_ (.A(_06011_),
    .B(_06317_),
    .C(_07213_),
    .D(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__nand2_4 _37738_ (.A(_07210_),
    .B(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__xor2_4 _37739_ (.A(_07206_),
    .B(_07217_),
    .X(_07218_));
 sky130_vsdinv _37740_ (.A(_07218_),
    .Y(_07219_));
 sky130_vsdinv _37741_ (.A(_07202_),
    .Y(_07220_));
 sky130_fd_sc_hd__and3_4 _37742_ (.A(_07220_),
    .B(_07201_),
    .C(_07200_),
    .X(_07221_));
 sky130_fd_sc_hd__or3_4 _37743_ (.A(_07203_),
    .B(_07219_),
    .C(_07221_),
    .X(_07222_));
 sky130_fd_sc_hd__o21ai_4 _37744_ (.A1(_07203_),
    .A2(_07221_),
    .B1(_07219_),
    .Y(_07223_));
 sky130_fd_sc_hd__nand2_4 _37745_ (.A(_07222_),
    .B(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__xor2_4 _37746_ (.A(_07186_),
    .B(_07224_),
    .X(_07225_));
 sky130_vsdinv _37747_ (.A(_07225_),
    .Y(_07226_));
 sky130_fd_sc_hd__nand2_4 _37748_ (.A(_07185_),
    .B(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__nand3_4 _37749_ (.A(_07183_),
    .B(_07225_),
    .C(_07184_),
    .Y(_07228_));
 sky130_fd_sc_hd__nand2_4 _37750_ (.A(_07227_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__nand2_4 _37751_ (.A(_07229_),
    .B(_07066_),
    .Y(_07230_));
 sky130_vsdinv _37752_ (.A(_07066_),
    .Y(_07231_));
 sky130_fd_sc_hd__nand3_4 _37753_ (.A(_07231_),
    .B(_07227_),
    .C(_07228_),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_4 _37754_ (.A(_07022_),
    .B(_07018_),
    .Y(_07233_));
 sky130_fd_sc_hd__xor2_4 _37755_ (.A(_07233_),
    .B(_07033_),
    .X(_07234_));
 sky130_vsdinv _37756_ (.A(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__a21o_4 _37757_ (.A1(_07230_),
    .A2(_07232_),
    .B1(_07235_),
    .X(_07236_));
 sky130_fd_sc_hd__nand3_4 _37758_ (.A(_07230_),
    .B(_07235_),
    .C(_07232_),
    .Y(_07237_));
 sky130_fd_sc_hd__nand2_4 _37759_ (.A(_07236_),
    .B(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__xnor2_4 _37760_ (.A(_07090_),
    .B(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__or2_4 _37761_ (.A(_07089_),
    .B(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__nand2_4 _37762_ (.A(_07239_),
    .B(_07089_),
    .Y(_07241_));
 sky130_fd_sc_hd__nand2_4 _37763_ (.A(_07081_),
    .B(_07076_),
    .Y(_07242_));
 sky130_fd_sc_hd__a21oi_4 _37764_ (.A1(_07240_),
    .A2(_07241_),
    .B1(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__nand3_4 _37765_ (.A(_07240_),
    .B(_07242_),
    .C(_07241_),
    .Y(_07244_));
 sky130_vsdinv _37766_ (.A(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__nor2_4 _37767_ (.A(_07243_),
    .B(_07245_),
    .Y(_07246_));
 sky130_vsdinv _37768_ (.A(_07086_),
    .Y(_07247_));
 sky130_fd_sc_hd__a21oi_4 _37769_ (.A1(_07088_),
    .A2(_07084_),
    .B1(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__xnor2_4 _37770_ (.A(_07246_),
    .B(_07248_),
    .Y(_01420_));
 sky130_fd_sc_hd__maj3_4 _37771_ (.A(_07206_),
    .B(_07207_),
    .C(_07209_),
    .X(_07249_));
 sky130_vsdinv _37772_ (.A(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_4 _37773_ (.A(_06444_),
    .B(_03492_),
    .Y(_07251_));
 sky130_fd_sc_hd__nand2_4 _37774_ (.A(_06447_),
    .B(_06947_),
    .Y(_07252_));
 sky130_fd_sc_hd__nand2_4 _37775_ (.A(_07251_),
    .B(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__nand4_4 _37776_ (.A(_06256_),
    .B(_06452_),
    .C(_07097_),
    .D(_06794_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand2_4 _37777_ (.A(_06456_),
    .B(_06797_),
    .Y(_07255_));
 sky130_vsdinv _37778_ (.A(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand3_4 _37779_ (.A(_07253_),
    .B(_07254_),
    .C(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__a21o_4 _37780_ (.A1(_07253_),
    .A2(_07254_),
    .B1(_07256_),
    .X(_07258_));
 sky130_fd_sc_hd__nand3_4 _37781_ (.A(_07250_),
    .B(_07257_),
    .C(_07258_),
    .Y(_07259_));
 sky130_fd_sc_hd__nand2_4 _37782_ (.A(_07258_),
    .B(_07257_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_4 _37783_ (.A(_07260_),
    .B(_07249_),
    .Y(_07261_));
 sky130_fd_sc_hd__a21boi_4 _37784_ (.A1(_07094_),
    .A2(_07100_),
    .B1_N(_07098_),
    .Y(_07262_));
 sky130_vsdinv _37785_ (.A(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__a21o_4 _37786_ (.A1(_07259_),
    .A2(_07261_),
    .B1(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__nand3_4 _37787_ (.A(_07259_),
    .B(_07263_),
    .C(_07261_),
    .Y(_07265_));
 sky130_vsdinv _37788_ (.A(_07221_),
    .Y(_07266_));
 sky130_fd_sc_hd__o21ai_4 _37789_ (.A1(_07203_),
    .A2(_07219_),
    .B1(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__a21oi_4 _37790_ (.A1(_07264_),
    .A2(_07265_),
    .B1(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__nand3_4 _37791_ (.A(_07264_),
    .B(_07267_),
    .C(_07265_),
    .Y(_07269_));
 sky130_vsdinv _37792_ (.A(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__maj3_4 _37793_ (.A(_07106_),
    .B(_07103_),
    .C(_07091_),
    .X(_07271_));
 sky130_fd_sc_hd__o21ai_4 _37794_ (.A1(_07268_),
    .A2(_07270_),
    .B1(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__a21o_4 _37795_ (.A1(_07264_),
    .A2(_07265_),
    .B1(_07267_),
    .X(_07273_));
 sky130_vsdinv _37796_ (.A(_07271_),
    .Y(_07274_));
 sky130_fd_sc_hd__nand3_4 _37797_ (.A(_07273_),
    .B(_07274_),
    .C(_07269_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand2_4 _37798_ (.A(_07272_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__nand3_4 _37799_ (.A(_07276_),
    .B(_07116_),
    .C(_07120_),
    .Y(_07277_));
 sky130_fd_sc_hd__nand2_4 _37800_ (.A(_07120_),
    .B(_07116_),
    .Y(_07278_));
 sky130_fd_sc_hd__nand3_4 _37801_ (.A(_07278_),
    .B(_07275_),
    .C(_07272_),
    .Y(_07279_));
 sky130_fd_sc_hd__buf_1 _37802_ (.A(_06846_),
    .X(_07280_));
 sky130_fd_sc_hd__nand2_4 _37803_ (.A(_07280_),
    .B(_06128_),
    .Y(_07281_));
 sky130_fd_sc_hd__nand2_4 _37804_ (.A(_06712_),
    .B(_06130_),
    .Y(_07282_));
 sky130_fd_sc_hd__nand2_4 _37805_ (.A(_07281_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__buf_1 _37806_ (.A(_06846_),
    .X(_07284_));
 sky130_fd_sc_hd__nand4_4 _37807_ (.A(_07284_),
    .B(_06712_),
    .C(_03465_),
    .D(_06220_),
    .Y(_07285_));
 sky130_fd_sc_hd__buf_1 _37808_ (.A(_03310_),
    .X(_07286_));
 sky130_fd_sc_hd__nand2_4 _37809_ (.A(_07286_),
    .B(_06232_),
    .Y(_07287_));
 sky130_vsdinv _37810_ (.A(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand3_4 _37811_ (.A(_07283_),
    .B(_07285_),
    .C(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__a21o_4 _37812_ (.A1(_07283_),
    .A2(_07285_),
    .B1(_07288_),
    .X(_07290_));
 sky130_fd_sc_hd__maj3_4 _37813_ (.A(_07136_),
    .B(_07129_),
    .C(_07133_),
    .X(_07291_));
 sky130_fd_sc_hd__a21boi_4 _37814_ (.A1(_07289_),
    .A2(_07290_),
    .B1_N(_07291_),
    .Y(_07292_));
 sky130_vsdinv _37815_ (.A(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__buf_1 _37816_ (.A(_03324_),
    .X(_07294_));
 sky130_fd_sc_hd__buf_1 _37817_ (.A(_07294_),
    .X(_07295_));
 sky130_fd_sc_hd__nand2_4 _37818_ (.A(_07295_),
    .B(_05956_),
    .Y(_07296_));
 sky130_fd_sc_hd__buf_1 _37819_ (.A(\pcpi_mul.rs1[14] ),
    .X(_07297_));
 sky130_fd_sc_hd__buf_1 _37820_ (.A(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__buf_1 _37821_ (.A(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__nand2_4 _37822_ (.A(_07299_),
    .B(_06003_),
    .Y(_07300_));
 sky130_fd_sc_hd__buf_1 _37823_ (.A(\pcpi_mul.rs1[15] ),
    .X(_07301_));
 sky130_fd_sc_hd__buf_1 _37824_ (.A(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__nand2_4 _37825_ (.A(_07302_),
    .B(_05947_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand2_4 _37826_ (.A(_07300_),
    .B(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__buf_1 _37827_ (.A(_07156_),
    .X(_07305_));
 sky130_fd_sc_hd__buf_1 _37828_ (.A(_07305_),
    .X(_07306_));
 sky130_fd_sc_hd__nand4_4 _37829_ (.A(_06993_),
    .B(_07306_),
    .C(_07002_),
    .D(_07154_),
    .Y(_07307_));
 sky130_fd_sc_hd__nand2_4 _37830_ (.A(_07304_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__xor2_4 _37831_ (.A(_07296_),
    .B(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__nand2_4 _37832_ (.A(_07290_),
    .B(_07289_),
    .Y(_07310_));
 sky130_fd_sc_hd__nor2_4 _37833_ (.A(_07291_),
    .B(_07310_),
    .Y(_07311_));
 sky130_vsdinv _37834_ (.A(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand3_4 _37835_ (.A(_07293_),
    .B(_07309_),
    .C(_07312_),
    .Y(_07313_));
 sky130_vsdinv _37836_ (.A(_07309_),
    .Y(_07314_));
 sky130_fd_sc_hd__o21ai_4 _37837_ (.A1(_07311_),
    .A2(_07292_),
    .B1(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__a21oi_4 _37838_ (.A1(_07143_),
    .A2(_07164_),
    .B1(_07140_),
    .Y(_07316_));
 sky130_vsdinv _37839_ (.A(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__a21o_4 _37840_ (.A1(_07313_),
    .A2(_07315_),
    .B1(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__nand3_4 _37841_ (.A(_07317_),
    .B(_07313_),
    .C(_07315_),
    .Y(_07319_));
 sky130_fd_sc_hd__a21boi_4 _37842_ (.A1(_07149_),
    .A2(_07160_),
    .B1_N(_07155_),
    .Y(_07320_));
 sky130_vsdinv _37843_ (.A(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__a21oi_4 _37844_ (.A1(_07318_),
    .A2(_07319_),
    .B1(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__nand3_4 _37845_ (.A(_07318_),
    .B(_07321_),
    .C(_07319_),
    .Y(_07323_));
 sky130_vsdinv _37846_ (.A(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__nor2_4 _37847_ (.A(_07322_),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__a21o_4 _37848_ (.A1(_07277_),
    .A2(_07279_),
    .B1(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__nand3_4 _37849_ (.A(_07277_),
    .B(_07279_),
    .C(_07325_),
    .Y(_07327_));
 sky130_fd_sc_hd__nand2_4 _37850_ (.A(_07326_),
    .B(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__a21boi_4 _37851_ (.A1(_07123_),
    .A2(_07176_),
    .B1_N(_07125_),
    .Y(_07329_));
 sky130_fd_sc_hd__nand2_4 _37852_ (.A(_07328_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand2_4 _37853_ (.A(_07179_),
    .B(_07125_),
    .Y(_07331_));
 sky130_fd_sc_hd__nand3_4 _37854_ (.A(_07331_),
    .B(_07327_),
    .C(_07326_),
    .Y(_07332_));
 sky130_fd_sc_hd__nand2_4 _37855_ (.A(_07330_),
    .B(_07332_),
    .Y(_07333_));
 sky130_vsdinv _37856_ (.A(_07186_),
    .Y(_07334_));
 sky130_fd_sc_hd__nand3_4 _37857_ (.A(_07222_),
    .B(_07223_),
    .C(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__nand2_4 _37858_ (.A(_05896_),
    .B(_03537_),
    .Y(_07336_));
 sky130_fd_sc_hd__buf_1 _37859_ (.A(_03530_),
    .X(_07337_));
 sky130_fd_sc_hd__nand2_4 _37860_ (.A(_05886_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand2_4 _37861_ (.A(_07336_),
    .B(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__nor2_4 _37862_ (.A(_07336_),
    .B(_07338_),
    .Y(_07340_));
 sky130_vsdinv _37863_ (.A(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__nand2_4 _37864_ (.A(_06945_),
    .B(_03496_),
    .Y(_07342_));
 sky130_fd_sc_hd__buf_1 _37865_ (.A(_03504_),
    .X(_07343_));
 sky130_fd_sc_hd__buf_1 _37866_ (.A(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__nand2_4 _37867_ (.A(_07208_),
    .B(_07344_),
    .Y(_07345_));
 sky130_fd_sc_hd__buf_1 _37868_ (.A(_03271_),
    .X(_07346_));
 sky130_fd_sc_hd__buf_1 _37869_ (.A(_06742_),
    .X(_07347_));
 sky130_fd_sc_hd__nand2_4 _37870_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__nand2_4 _37871_ (.A(_07345_),
    .B(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand4_4 _37872_ (.A(_06317_),
    .B(_06170_),
    .C(_03501_),
    .D(_06748_),
    .Y(_07350_));
 sky130_fd_sc_hd__nand2_4 _37873_ (.A(_07349_),
    .B(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__xnor2_4 _37874_ (.A(_07342_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__buf_1 _37875_ (.A(_03524_),
    .X(_07353_));
 sky130_fd_sc_hd__nand2_4 _37876_ (.A(_06380_),
    .B(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__buf_1 _37877_ (.A(\pcpi_mul.rs2[13] ),
    .X(_07355_));
 sky130_fd_sc_hd__buf_1 _37878_ (.A(_07355_),
    .X(_07356_));
 sky130_fd_sc_hd__nand2_4 _37879_ (.A(_06226_),
    .B(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__nand2_4 _37880_ (.A(_07354_),
    .B(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__buf_1 _37881_ (.A(_05899_),
    .X(_07359_));
 sky130_fd_sc_hd__buf_1 _37882_ (.A(_06383_),
    .X(_07360_));
 sky130_fd_sc_hd__buf_1 _37883_ (.A(\pcpi_mul.rs2[14] ),
    .X(_07361_));
 sky130_fd_sc_hd__buf_8 _37884_ (.A(_07361_),
    .X(_07362_));
 sky130_fd_sc_hd__nand4_4 _37885_ (.A(_07359_),
    .B(_07360_),
    .C(_03517_),
    .D(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__buf_1 _37886_ (.A(\pcpi_mul.rs1[4] ),
    .X(_07364_));
 sky130_fd_sc_hd__buf_1 _37887_ (.A(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__buf_1 _37888_ (.A(_07043_),
    .X(_07366_));
 sky130_fd_sc_hd__nand2_4 _37889_ (.A(_07365_),
    .B(_07366_),
    .Y(_07367_));
 sky130_vsdinv _37890_ (.A(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__nand3_4 _37891_ (.A(_07358_),
    .B(_07363_),
    .C(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__nand2_4 _37892_ (.A(_07358_),
    .B(_07363_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand2_4 _37893_ (.A(_07370_),
    .B(_07367_),
    .Y(_07371_));
 sky130_fd_sc_hd__a21boi_4 _37894_ (.A1(_07191_),
    .A2(_07199_),
    .B1_N(_07195_),
    .Y(_07372_));
 sky130_fd_sc_hd__a21boi_4 _37895_ (.A1(_07369_),
    .A2(_07371_),
    .B1_N(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__nand2_4 _37896_ (.A(_07371_),
    .B(_07369_),
    .Y(_07374_));
 sky130_fd_sc_hd__nor2_4 _37897_ (.A(_07372_),
    .B(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__nor2_4 _37898_ (.A(_07373_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__xnor2_4 _37899_ (.A(_07352_),
    .B(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__a21o_4 _37900_ (.A1(_07339_),
    .A2(_07341_),
    .B1(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__nand2_4 _37901_ (.A(_07341_),
    .B(_07339_),
    .Y(_07379_));
 sky130_vsdinv _37902_ (.A(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__nand2_4 _37903_ (.A(_07377_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__nand2_4 _37904_ (.A(_07378_),
    .B(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__xor2_4 _37905_ (.A(_07335_),
    .B(_07382_),
    .X(_07383_));
 sky130_vsdinv _37906_ (.A(_07383_),
    .Y(_07384_));
 sky130_fd_sc_hd__nand2_4 _37907_ (.A(_07333_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__nand3_4 _37908_ (.A(_07330_),
    .B(_07332_),
    .C(_07383_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand2_4 _37909_ (.A(_07385_),
    .B(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__nand2_4 _37910_ (.A(_07387_),
    .B(_07228_),
    .Y(_07388_));
 sky130_vsdinv _37911_ (.A(_07228_),
    .Y(_07389_));
 sky130_fd_sc_hd__nand3_4 _37912_ (.A(_07389_),
    .B(_07385_),
    .C(_07386_),
    .Y(_07390_));
 sky130_fd_sc_hd__nand2_4 _37913_ (.A(_07388_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__nand2_4 _37914_ (.A(_07174_),
    .B(_07170_),
    .Y(_07392_));
 sky130_fd_sc_hd__xor2_4 _37915_ (.A(_07392_),
    .B(_07184_),
    .X(_07393_));
 sky130_fd_sc_hd__nand2_4 _37916_ (.A(_07391_),
    .B(_07393_),
    .Y(_07394_));
 sky130_vsdinv _37917_ (.A(_07393_),
    .Y(_07395_));
 sky130_fd_sc_hd__nand3_4 _37918_ (.A(_07388_),
    .B(_07395_),
    .C(_07390_),
    .Y(_07396_));
 sky130_fd_sc_hd__nand2_4 _37919_ (.A(_07394_),
    .B(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__a21boi_4 _37920_ (.A1(_07230_),
    .A2(_07235_),
    .B1_N(_07232_),
    .Y(_07398_));
 sky130_fd_sc_hd__nand2_4 _37921_ (.A(_07397_),
    .B(_07398_),
    .Y(_07399_));
 sky130_fd_sc_hd__nand2_4 _37922_ (.A(_07237_),
    .B(_07232_),
    .Y(_07400_));
 sky130_fd_sc_hd__nand3_4 _37923_ (.A(_07400_),
    .B(_07396_),
    .C(_07394_),
    .Y(_07401_));
 sky130_fd_sc_hd__nand4_4 _37924_ (.A(_07032_),
    .B(_07026_),
    .C(_07028_),
    .D(_07233_),
    .Y(_07402_));
 sky130_vsdinv _37925_ (.A(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__a21o_4 _37926_ (.A1(_07399_),
    .A2(_07401_),
    .B1(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__nand3_4 _37927_ (.A(_07399_),
    .B(_07401_),
    .C(_07403_),
    .Y(_07405_));
 sky130_vsdinv _37928_ (.A(_07089_),
    .Y(_07406_));
 sky130_fd_sc_hd__a21oi_4 _37929_ (.A1(_07236_),
    .A2(_07237_),
    .B1(_07090_),
    .Y(_07407_));
 sky130_fd_sc_hd__nand3_4 _37930_ (.A(_07090_),
    .B(_07236_),
    .C(_07237_),
    .Y(_07408_));
 sky130_fd_sc_hd__o21ai_4 _37931_ (.A1(_07406_),
    .A2(_07407_),
    .B1(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__a21oi_4 _37932_ (.A1(_07404_),
    .A2(_07405_),
    .B1(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__nand3_4 _37933_ (.A(_07409_),
    .B(_07404_),
    .C(_07405_),
    .Y(_07411_));
 sky130_vsdinv _37934_ (.A(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__nor2_4 _37935_ (.A(_07410_),
    .B(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__o21ai_4 _37936_ (.A1(_07243_),
    .A2(_07248_),
    .B1(_07244_),
    .Y(_07414_));
 sky130_fd_sc_hd__buf_1 _37937_ (.A(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__xor2_4 _37938_ (.A(_07413_),
    .B(_07415_),
    .X(_01421_));
 sky130_fd_sc_hd__buf_1 _37939_ (.A(_03303_),
    .X(_07416_));
 sky130_fd_sc_hd__nand2_4 _37940_ (.A(_07416_),
    .B(_06138_),
    .Y(_07417_));
 sky130_fd_sc_hd__nand2_4 _37941_ (.A(_07286_),
    .B(_06318_),
    .Y(_07418_));
 sky130_fd_sc_hd__nand2_4 _37942_ (.A(_07417_),
    .B(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__nand4_4 _37943_ (.A(_07416_),
    .B(_07286_),
    .C(_06318_),
    .D(_06229_),
    .Y(_07420_));
 sky130_fd_sc_hd__buf_1 _37944_ (.A(\pcpi_mul.rs1[14] ),
    .X(_07421_));
 sky130_fd_sc_hd__buf_1 _37945_ (.A(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__nand2_4 _37946_ (.A(_07422_),
    .B(_06551_),
    .Y(_07423_));
 sky130_vsdinv _37947_ (.A(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__a21o_4 _37948_ (.A1(_07419_),
    .A2(_07420_),
    .B1(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__nand3_4 _37949_ (.A(_07419_),
    .B(_07420_),
    .C(_07424_),
    .Y(_07426_));
 sky130_fd_sc_hd__a21boi_4 _37950_ (.A1(_07283_),
    .A2(_07288_),
    .B1_N(_07285_),
    .Y(_07427_));
 sky130_fd_sc_hd__a21boi_4 _37951_ (.A1(_07425_),
    .A2(_07426_),
    .B1_N(_07427_),
    .Y(_07428_));
 sky130_vsdinv _37952_ (.A(_07427_),
    .Y(_07429_));
 sky130_fd_sc_hd__nand3_4 _37953_ (.A(_07429_),
    .B(_07426_),
    .C(_07425_),
    .Y(_07430_));
 sky130_vsdinv _37954_ (.A(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__buf_1 _37955_ (.A(_03317_),
    .X(_07432_));
 sky130_fd_sc_hd__nand2_4 _37956_ (.A(_07432_),
    .B(_06705_),
    .Y(_07433_));
 sky130_fd_sc_hd__buf_1 _37957_ (.A(\pcpi_mul.rs1[16] ),
    .X(_07434_));
 sky130_fd_sc_hd__buf_1 _37958_ (.A(_07434_),
    .X(_07435_));
 sky130_fd_sc_hd__nand2_4 _37959_ (.A(_07435_),
    .B(_07001_),
    .Y(_07436_));
 sky130_fd_sc_hd__nand2_4 _37960_ (.A(_07433_),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__buf_1 _37961_ (.A(\pcpi_mul.rs1[15] ),
    .X(_07438_));
 sky130_fd_sc_hd__buf_1 _37962_ (.A(_07438_),
    .X(_07439_));
 sky130_fd_sc_hd__buf_1 _37963_ (.A(_06012_),
    .X(_07440_));
 sky130_fd_sc_hd__nand4_4 _37964_ (.A(_07439_),
    .B(_07294_),
    .C(_07440_),
    .D(_05939_),
    .Y(_07441_));
 sky130_fd_sc_hd__buf_1 _37965_ (.A(\pcpi_mul.rs1[17] ),
    .X(_07442_));
 sky130_fd_sc_hd__buf_1 _37966_ (.A(_07442_),
    .X(_07443_));
 sky130_fd_sc_hd__buf_1 _37967_ (.A(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__nand2_4 _37968_ (.A(_07444_),
    .B(_05955_),
    .Y(_07445_));
 sky130_vsdinv _37969_ (.A(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__a21o_4 _37970_ (.A1(_07437_),
    .A2(_07441_),
    .B1(_07446_),
    .X(_07447_));
 sky130_fd_sc_hd__nand3_4 _37971_ (.A(_07437_),
    .B(_07441_),
    .C(_07446_),
    .Y(_07448_));
 sky130_fd_sc_hd__and2_4 _37972_ (.A(_07447_),
    .B(_07448_),
    .X(_07449_));
 sky130_vsdinv _37973_ (.A(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__o21ai_4 _37974_ (.A1(_07428_),
    .A2(_07431_),
    .B1(_07450_),
    .Y(_07451_));
 sky130_vsdinv _37975_ (.A(_07428_),
    .Y(_07452_));
 sky130_fd_sc_hd__nand3_4 _37976_ (.A(_07452_),
    .B(_07449_),
    .C(_07430_),
    .Y(_07453_));
 sky130_fd_sc_hd__o21ai_4 _37977_ (.A1(_07292_),
    .A2(_07314_),
    .B1(_07312_),
    .Y(_07454_));
 sky130_fd_sc_hd__a21o_4 _37978_ (.A1(_07451_),
    .A2(_07453_),
    .B1(_07454_),
    .X(_07455_));
 sky130_fd_sc_hd__nand3_4 _37979_ (.A(_07454_),
    .B(_07451_),
    .C(_07453_),
    .Y(_07456_));
 sky130_fd_sc_hd__nand2_4 _37980_ (.A(_07455_),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__maj3_4 _37981_ (.A(_07300_),
    .B(_07303_),
    .C(_07296_),
    .X(_07458_));
 sky130_fd_sc_hd__nand2_4 _37982_ (.A(_07457_),
    .B(_07458_),
    .Y(_07459_));
 sky130_vsdinv _37983_ (.A(_07458_),
    .Y(_07460_));
 sky130_fd_sc_hd__nand3_4 _37984_ (.A(_07455_),
    .B(_07456_),
    .C(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__and2_4 _37985_ (.A(_07459_),
    .B(_07461_),
    .X(_07462_));
 sky130_vsdinv _37986_ (.A(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__buf_1 _37987_ (.A(\pcpi_mul.rs1[9] ),
    .X(_07464_));
 sky130_fd_sc_hd__buf_1 _37988_ (.A(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__nand2_4 _37989_ (.A(_07465_),
    .B(_06482_),
    .Y(_07466_));
 sky130_fd_sc_hd__buf_1 _37990_ (.A(_03480_),
    .X(_07467_));
 sky130_fd_sc_hd__nand2_4 _37991_ (.A(_06567_),
    .B(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__nand2_4 _37992_ (.A(_07466_),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__buf_1 _37993_ (.A(_06593_),
    .X(_07470_));
 sky130_fd_sc_hd__nand4_4 _37994_ (.A(_06350_),
    .B(_06977_),
    .C(_06791_),
    .D(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nand2_4 _37995_ (.A(_07280_),
    .B(_06949_),
    .Y(_07472_));
 sky130_vsdinv _37996_ (.A(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__a21o_4 _37997_ (.A1(_07469_),
    .A2(_07471_),
    .B1(_07473_),
    .X(_07474_));
 sky130_fd_sc_hd__nand3_4 _37998_ (.A(_07469_),
    .B(_07471_),
    .C(_07473_),
    .Y(_07475_));
 sky130_fd_sc_hd__nand2_4 _37999_ (.A(_07474_),
    .B(_07475_),
    .Y(_07476_));
 sky130_fd_sc_hd__maj3_4 _38000_ (.A(_07342_),
    .B(_07345_),
    .C(_07348_),
    .X(_07477_));
 sky130_fd_sc_hd__nand2_4 _38001_ (.A(_07476_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__o21ai_4 _38002_ (.A1(_07342_),
    .A2(_07351_),
    .B1(_07350_),
    .Y(_07479_));
 sky130_fd_sc_hd__nand3_4 _38003_ (.A(_07479_),
    .B(_07475_),
    .C(_07474_),
    .Y(_07480_));
 sky130_fd_sc_hd__nand2_4 _38004_ (.A(_07478_),
    .B(_07480_),
    .Y(_07481_));
 sky130_fd_sc_hd__a21boi_4 _38005_ (.A1(_07253_),
    .A2(_07256_),
    .B1_N(_07254_),
    .Y(_07482_));
 sky130_fd_sc_hd__nand2_4 _38006_ (.A(_07481_),
    .B(_07482_),
    .Y(_07483_));
 sky130_vsdinv _38007_ (.A(_07482_),
    .Y(_07484_));
 sky130_fd_sc_hd__nand3_4 _38008_ (.A(_07478_),
    .B(_07480_),
    .C(_07484_),
    .Y(_07485_));
 sky130_fd_sc_hd__nand2_4 _38009_ (.A(_07483_),
    .B(_07485_),
    .Y(_07486_));
 sky130_vsdinv _38010_ (.A(_07375_),
    .Y(_07487_));
 sky130_fd_sc_hd__o21ai_4 _38011_ (.A1(_07352_),
    .A2(_07373_),
    .B1(_07487_),
    .Y(_07488_));
 sky130_vsdinv _38012_ (.A(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__nand2_4 _38013_ (.A(_07486_),
    .B(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__nand3_4 _38014_ (.A(_07488_),
    .B(_07483_),
    .C(_07485_),
    .Y(_07491_));
 sky130_fd_sc_hd__nand2_4 _38015_ (.A(_07490_),
    .B(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__maj3_4 _38016_ (.A(_07262_),
    .B(_07260_),
    .C(_07249_),
    .X(_07493_));
 sky130_fd_sc_hd__nand2_4 _38017_ (.A(_07492_),
    .B(_07493_),
    .Y(_07494_));
 sky130_vsdinv _38018_ (.A(_07493_),
    .Y(_07495_));
 sky130_fd_sc_hd__nand3_4 _38019_ (.A(_07490_),
    .B(_07495_),
    .C(_07491_),
    .Y(_07496_));
 sky130_fd_sc_hd__nand2_4 _38020_ (.A(_07494_),
    .B(_07496_),
    .Y(_07497_));
 sky130_fd_sc_hd__a21oi_4 _38021_ (.A1(_07273_),
    .A2(_07274_),
    .B1(_07270_),
    .Y(_07498_));
 sky130_fd_sc_hd__nand2_4 _38022_ (.A(_07497_),
    .B(_07498_),
    .Y(_07499_));
 sky130_fd_sc_hd__o21ai_4 _38023_ (.A1(_07271_),
    .A2(_07268_),
    .B1(_07269_),
    .Y(_07500_));
 sky130_fd_sc_hd__nand3_4 _38024_ (.A(_07500_),
    .B(_07496_),
    .C(_07494_),
    .Y(_07501_));
 sky130_fd_sc_hd__nand2_4 _38025_ (.A(_07499_),
    .B(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__nand2_4 _38026_ (.A(_07463_),
    .B(_07502_),
    .Y(_07503_));
 sky130_fd_sc_hd__nand3_4 _38027_ (.A(_07462_),
    .B(_07501_),
    .C(_07499_),
    .Y(_07504_));
 sky130_fd_sc_hd__nand2_4 _38028_ (.A(_07503_),
    .B(_07504_),
    .Y(_07505_));
 sky130_vsdinv _38029_ (.A(_07335_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand3_4 _38030_ (.A(_07378_),
    .B(_07506_),
    .C(_07381_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand2_4 _38031_ (.A(_07505_),
    .B(_07507_),
    .Y(_07508_));
 sky130_vsdinv _38032_ (.A(_07507_),
    .Y(_07509_));
 sky130_fd_sc_hd__nand3_4 _38033_ (.A(_07503_),
    .B(_07509_),
    .C(_07504_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand2_4 _38034_ (.A(_07508_),
    .B(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__a21boi_4 _38035_ (.A1(_07277_),
    .A2(_07325_),
    .B1_N(_07279_),
    .Y(_07512_));
 sky130_fd_sc_hd__nand2_4 _38036_ (.A(_07511_),
    .B(_07512_),
    .Y(_07513_));
 sky130_vsdinv _38037_ (.A(_07512_),
    .Y(_07514_));
 sky130_fd_sc_hd__nand3_4 _38038_ (.A(_07508_),
    .B(_07514_),
    .C(_07510_),
    .Y(_07515_));
 sky130_fd_sc_hd__nand2_4 _38039_ (.A(_07513_),
    .B(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__nand2_4 _38040_ (.A(_07196_),
    .B(_07055_),
    .Y(_07517_));
 sky130_fd_sc_hd__buf_1 _38041_ (.A(_07058_),
    .X(_07518_));
 sky130_fd_sc_hd__nand2_4 _38042_ (.A(_06142_),
    .B(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__nand2_4 _38043_ (.A(_07517_),
    .B(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__buf_1 _38044_ (.A(_07355_),
    .X(_07521_));
 sky130_fd_sc_hd__buf_1 _38045_ (.A(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__buf_1 _38046_ (.A(_03525_),
    .X(_07523_));
 sky130_fd_sc_hd__nand4_4 _38047_ (.A(_06227_),
    .B(_06072_),
    .C(_07522_),
    .D(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__buf_1 _38048_ (.A(_03267_),
    .X(_07525_));
 sky130_fd_sc_hd__buf_1 _38049_ (.A(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__nand2_4 _38050_ (.A(_07526_),
    .B(_07045_),
    .Y(_07527_));
 sky130_vsdinv _38051_ (.A(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__nand3_4 _38052_ (.A(_07520_),
    .B(_07524_),
    .C(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__nand2_4 _38053_ (.A(_07520_),
    .B(_07524_),
    .Y(_07530_));
 sky130_fd_sc_hd__nand2_4 _38054_ (.A(_07530_),
    .B(_07527_),
    .Y(_07531_));
 sky130_fd_sc_hd__a21boi_4 _38055_ (.A1(_07358_),
    .A2(_07368_),
    .B1_N(_07363_),
    .Y(_07532_));
 sky130_fd_sc_hd__a21boi_4 _38056_ (.A1(_07529_),
    .A2(_07531_),
    .B1_N(_07532_),
    .Y(_07533_));
 sky130_fd_sc_hd__nand2_4 _38057_ (.A(_07531_),
    .B(_07529_),
    .Y(_07534_));
 sky130_fd_sc_hd__nor2_4 _38058_ (.A(_07532_),
    .B(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__nand2_4 _38059_ (.A(_06347_),
    .B(_03496_),
    .Y(_07536_));
 sky130_fd_sc_hd__buf_1 _38060_ (.A(_06636_),
    .X(_07537_));
 sky130_fd_sc_hd__nand2_4 _38061_ (.A(_06245_),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand2_4 _38062_ (.A(_06945_),
    .B(_06632_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_4 _38063_ (.A(_07538_),
    .B(_07539_),
    .Y(_07540_));
 sky130_fd_sc_hd__buf_1 _38064_ (.A(_07211_),
    .X(_07541_));
 sky130_fd_sc_hd__buf_1 _38065_ (.A(_07541_),
    .X(_07542_));
 sky130_fd_sc_hd__buf_1 _38066_ (.A(_06635_),
    .X(_07543_));
 sky130_fd_sc_hd__buf_1 _38067_ (.A(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__nand4_4 _38068_ (.A(_06245_),
    .B(_06248_),
    .C(_07542_),
    .D(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__nand2_4 _38069_ (.A(_07540_),
    .B(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__xor2_4 _38070_ (.A(_07536_),
    .B(_07546_),
    .X(_07547_));
 sky130_vsdinv _38071_ (.A(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__o21ai_4 _38072_ (.A1(_07533_),
    .A2(_07535_),
    .B1(_07548_),
    .Y(_07549_));
 sky130_vsdinv _38073_ (.A(_07535_),
    .Y(_07550_));
 sky130_vsdinv _38074_ (.A(_07533_),
    .Y(_07551_));
 sky130_fd_sc_hd__nand3_4 _38075_ (.A(_07550_),
    .B(_07551_),
    .C(_07547_),
    .Y(_07552_));
 sky130_fd_sc_hd__buf_1 _38076_ (.A(_03534_),
    .X(_07553_));
 sky130_fd_sc_hd__buf_1 _38077_ (.A(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__nand2_4 _38078_ (.A(_06371_),
    .B(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__buf_1 _38079_ (.A(_03539_),
    .X(_07556_));
 sky130_fd_sc_hd__buf_1 _38080_ (.A(_07556_),
    .X(_07557_));
 sky130_fd_sc_hd__nand2_4 _38081_ (.A(_05895_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__nand2_4 _38082_ (.A(_07555_),
    .B(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__nand4_4 _38083_ (.A(_05585_),
    .B(_05886_),
    .C(_03537_),
    .D(_03542_),
    .Y(_07560_));
 sky130_fd_sc_hd__buf_1 _38084_ (.A(\pcpi_mul.rs2[15] ),
    .X(_07561_));
 sky130_fd_sc_hd__buf_1 _38085_ (.A(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__buf_1 _38086_ (.A(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__nand2_4 _38087_ (.A(_06381_),
    .B(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__a21bo_4 _38088_ (.A1(_07559_),
    .A2(_07560_),
    .B1_N(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__nand4_4 _38089_ (.A(_05902_),
    .B(_07559_),
    .C(_07560_),
    .D(_03532_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_4 _38090_ (.A(_07565_),
    .B(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__xor2_4 _38091_ (.A(_07341_),
    .B(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__a21o_4 _38092_ (.A1(_07549_),
    .A2(_07552_),
    .B1(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__nand3_4 _38093_ (.A(_07568_),
    .B(_07549_),
    .C(_07552_),
    .Y(_07570_));
 sky130_fd_sc_hd__nand2_4 _38094_ (.A(_07569_),
    .B(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__xor2_4 _38095_ (.A(_07571_),
    .B(_07381_),
    .X(_07572_));
 sky130_vsdinv _38096_ (.A(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__nand2_4 _38097_ (.A(_07516_),
    .B(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__nand3_4 _38098_ (.A(_07513_),
    .B(_07572_),
    .C(_07515_),
    .Y(_07575_));
 sky130_fd_sc_hd__buf_1 _38099_ (.A(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__nand2_4 _38100_ (.A(_07574_),
    .B(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__nand2_4 _38101_ (.A(_07577_),
    .B(_07386_),
    .Y(_07578_));
 sky130_vsdinv _38102_ (.A(_07386_),
    .Y(_07579_));
 sky130_fd_sc_hd__nand3_4 _38103_ (.A(_07574_),
    .B(_07579_),
    .C(_07576_),
    .Y(_07580_));
 sky130_fd_sc_hd__nand2_4 _38104_ (.A(_07578_),
    .B(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__nand2_4 _38105_ (.A(_07323_),
    .B(_07319_),
    .Y(_07582_));
 sky130_fd_sc_hd__xor2_4 _38106_ (.A(_07582_),
    .B(_07332_),
    .X(_07583_));
 sky130_fd_sc_hd__nand2_4 _38107_ (.A(_07581_),
    .B(_07583_),
    .Y(_07584_));
 sky130_vsdinv _38108_ (.A(_07583_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand3_4 _38109_ (.A(_07578_),
    .B(_07585_),
    .C(_07580_),
    .Y(_07586_));
 sky130_fd_sc_hd__nand2_4 _38110_ (.A(_07584_),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__a21boi_4 _38111_ (.A1(_07388_),
    .A2(_07395_),
    .B1_N(_07390_),
    .Y(_07588_));
 sky130_fd_sc_hd__nand2_4 _38112_ (.A(_07587_),
    .B(_07588_),
    .Y(_07589_));
 sky130_vsdinv _38113_ (.A(_07588_),
    .Y(_07590_));
 sky130_fd_sc_hd__nand3_4 _38114_ (.A(_07590_),
    .B(_07584_),
    .C(_07586_),
    .Y(_07591_));
 sky130_fd_sc_hd__nand2_4 _38115_ (.A(_07589_),
    .B(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__nand4_4 _38116_ (.A(_07181_),
    .B(_07178_),
    .C(_07179_),
    .D(_07392_),
    .Y(_07593_));
 sky130_fd_sc_hd__nand2_4 _38117_ (.A(_07592_),
    .B(_07593_),
    .Y(_07594_));
 sky130_vsdinv _38118_ (.A(_07593_),
    .Y(_07595_));
 sky130_fd_sc_hd__nand3_4 _38119_ (.A(_07589_),
    .B(_07595_),
    .C(_07591_),
    .Y(_07596_));
 sky130_fd_sc_hd__nand2_4 _38120_ (.A(_07594_),
    .B(_07596_),
    .Y(_07597_));
 sky130_fd_sc_hd__nand2_4 _38121_ (.A(_07405_),
    .B(_07401_),
    .Y(_07598_));
 sky130_vsdinv _38122_ (.A(_07598_),
    .Y(_07599_));
 sky130_fd_sc_hd__nand2_4 _38123_ (.A(_07597_),
    .B(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__nand3_4 _38124_ (.A(_07594_),
    .B(_07596_),
    .C(_07598_),
    .Y(_07601_));
 sky130_fd_sc_hd__nand2_4 _38125_ (.A(_07600_),
    .B(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__a21oi_4 _38126_ (.A1(_07415_),
    .A2(_07413_),
    .B1(_07412_),
    .Y(_07603_));
 sky130_fd_sc_hd__xor2_4 _38127_ (.A(_07602_),
    .B(_07603_),
    .X(_01422_));
 sky130_fd_sc_hd__nand2_4 _38128_ (.A(_07000_),
    .B(_07128_),
    .Y(_07604_));
 sky130_fd_sc_hd__buf_1 _38129_ (.A(_07298_),
    .X(_07605_));
 sky130_fd_sc_hd__nand2_4 _38130_ (.A(_07605_),
    .B(_07132_),
    .Y(_07606_));
 sky130_fd_sc_hd__nand2_4 _38131_ (.A(_07604_),
    .B(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__nand4_4 _38132_ (.A(_07000_),
    .B(_07605_),
    .C(_06427_),
    .D(_06696_),
    .Y(_07608_));
 sky130_fd_sc_hd__nand2_4 _38133_ (.A(_07306_),
    .B(_06328_),
    .Y(_07609_));
 sky130_vsdinv _38134_ (.A(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__nand3_4 _38135_ (.A(_07607_),
    .B(_07608_),
    .C(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__a21o_4 _38136_ (.A1(_07607_),
    .A2(_07608_),
    .B1(_07610_),
    .X(_07612_));
 sky130_fd_sc_hd__a21boi_4 _38137_ (.A1(_07419_),
    .A2(_07424_),
    .B1_N(_07420_),
    .Y(_07613_));
 sky130_vsdinv _38138_ (.A(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__a21o_4 _38139_ (.A1(_07611_),
    .A2(_07612_),
    .B1(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__nand3_4 _38140_ (.A(_07614_),
    .B(_07611_),
    .C(_07612_),
    .Y(_07616_));
 sky130_fd_sc_hd__nand2_4 _38141_ (.A(_07615_),
    .B(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__buf_1 _38142_ (.A(_05891_),
    .X(_07618_));
 sky130_fd_sc_hd__buf_1 _38143_ (.A(_07618_),
    .X(_07619_));
 sky130_fd_sc_hd__buf_1 _38144_ (.A(_07434_),
    .X(_07620_));
 sky130_fd_sc_hd__buf_1 _38145_ (.A(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__nand2_4 _38146_ (.A(_07621_),
    .B(_06003_),
    .Y(_07622_));
 sky130_fd_sc_hd__o21ai_4 _38147_ (.A1(_03333_),
    .A2(_07619_),
    .B1(_07622_),
    .Y(_07623_));
 sky130_fd_sc_hd__buf_1 _38148_ (.A(_07434_),
    .X(_07624_));
 sky130_fd_sc_hd__buf_1 _38149_ (.A(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__buf_1 _38150_ (.A(_03331_),
    .X(_07626_));
 sky130_fd_sc_hd__buf_1 _38151_ (.A(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__nand4_4 _38152_ (.A(_07625_),
    .B(_07627_),
    .C(_06165_),
    .D(_06706_),
    .Y(_07628_));
 sky130_fd_sc_hd__buf_1 _38153_ (.A(_03335_),
    .X(_07629_));
 sky130_fd_sc_hd__buf_1 _38154_ (.A(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__nand2_4 _38155_ (.A(_07630_),
    .B(_06021_),
    .Y(_07631_));
 sky130_vsdinv _38156_ (.A(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__a21oi_4 _38157_ (.A1(_07623_),
    .A2(_07628_),
    .B1(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand3_4 _38158_ (.A(_07623_),
    .B(_07628_),
    .C(_07632_),
    .Y(_07634_));
 sky130_vsdinv _38159_ (.A(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__nor2_4 _38160_ (.A(_07633_),
    .B(_07635_),
    .Y(_07636_));
 sky130_vsdinv _38161_ (.A(_07636_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_4 _38162_ (.A(_07617_),
    .B(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand3_4 _38163_ (.A(_07615_),
    .B(_07636_),
    .C(_07616_),
    .Y(_07639_));
 sky130_fd_sc_hd__nand2_4 _38164_ (.A(_07638_),
    .B(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__o21ai_4 _38165_ (.A1(_07428_),
    .A2(_07450_),
    .B1(_07430_),
    .Y(_07641_));
 sky130_vsdinv _38166_ (.A(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__nand2_4 _38167_ (.A(_07640_),
    .B(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__nand3_4 _38168_ (.A(_07638_),
    .B(_07641_),
    .C(_07639_),
    .Y(_07644_));
 sky130_fd_sc_hd__nand2_4 _38169_ (.A(_07643_),
    .B(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__a21boi_4 _38170_ (.A1(_07437_),
    .A2(_07446_),
    .B1_N(_07441_),
    .Y(_07646_));
 sky130_fd_sc_hd__nand2_4 _38171_ (.A(_07645_),
    .B(_07646_),
    .Y(_07647_));
 sky130_vsdinv _38172_ (.A(_07646_),
    .Y(_07648_));
 sky130_fd_sc_hd__nand3_4 _38173_ (.A(_07643_),
    .B(_07644_),
    .C(_07648_),
    .Y(_07649_));
 sky130_fd_sc_hd__and2_4 _38174_ (.A(_07647_),
    .B(_07649_),
    .X(_07650_));
 sky130_vsdinv _38175_ (.A(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__o21ai_4 _38176_ (.A1(_07533_),
    .A2(_07548_),
    .B1(_07550_),
    .Y(_07652_));
 sky130_fd_sc_hd__buf_1 _38177_ (.A(_03293_),
    .X(_07653_));
 sky130_fd_sc_hd__buf_1 _38178_ (.A(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__nand2_4 _38179_ (.A(_07654_),
    .B(_06939_),
    .Y(_07655_));
 sky130_fd_sc_hd__nand2_4 _38180_ (.A(_06571_),
    .B(_07467_),
    .Y(_07656_));
 sky130_fd_sc_hd__nand2_4 _38181_ (.A(_07655_),
    .B(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__nand4_4 _38182_ (.A(_06977_),
    .B(_07284_),
    .C(_06600_),
    .D(_06594_),
    .Y(_07658_));
 sky130_fd_sc_hd__nand2_4 _38183_ (.A(_07657_),
    .B(_07658_),
    .Y(_07659_));
 sky130_fd_sc_hd__buf_1 _38184_ (.A(_06848_),
    .X(_07660_));
 sky130_fd_sc_hd__nand2_4 _38185_ (.A(_07660_),
    .B(_06606_),
    .Y(_07661_));
 sky130_fd_sc_hd__nand2_4 _38186_ (.A(_07659_),
    .B(_07661_),
    .Y(_07662_));
 sky130_vsdinv _38187_ (.A(_07661_),
    .Y(_07663_));
 sky130_fd_sc_hd__nand3_4 _38188_ (.A(_07657_),
    .B(_07658_),
    .C(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__nand2_4 _38189_ (.A(_07662_),
    .B(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__maj3_4 _38190_ (.A(_07536_),
    .B(_07538_),
    .C(_07539_),
    .X(_07666_));
 sky130_fd_sc_hd__nand2_4 _38191_ (.A(_07665_),
    .B(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__buf_1 _38192_ (.A(_07343_),
    .X(_07668_));
 sky130_fd_sc_hd__buf_1 _38193_ (.A(_07668_),
    .X(_07669_));
 sky130_fd_sc_hd__a22oi_4 _38194_ (.A1(_06171_),
    .A2(_07669_),
    .B1(_06156_),
    .B2(_06507_),
    .Y(_07670_));
 sky130_fd_sc_hd__o21ai_4 _38195_ (.A1(_07536_),
    .A2(_07670_),
    .B1(_07545_),
    .Y(_07671_));
 sky130_fd_sc_hd__nand3_4 _38196_ (.A(_07671_),
    .B(_07664_),
    .C(_07662_),
    .Y(_07672_));
 sky130_fd_sc_hd__a21boi_4 _38197_ (.A1(_07469_),
    .A2(_07473_),
    .B1_N(_07471_),
    .Y(_07673_));
 sky130_vsdinv _38198_ (.A(_07673_),
    .Y(_07674_));
 sky130_fd_sc_hd__nand3_4 _38199_ (.A(_07667_),
    .B(_07672_),
    .C(_07674_),
    .Y(_07675_));
 sky130_fd_sc_hd__nand2_4 _38200_ (.A(_07667_),
    .B(_07672_),
    .Y(_07676_));
 sky130_fd_sc_hd__nand2_4 _38201_ (.A(_07676_),
    .B(_07673_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand3_4 _38202_ (.A(_07652_),
    .B(_07675_),
    .C(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__a21oi_4 _38203_ (.A1(_07551_),
    .A2(_07547_),
    .B1(_07535_),
    .Y(_07679_));
 sky130_fd_sc_hd__nand2_4 _38204_ (.A(_07677_),
    .B(_07675_),
    .Y(_07680_));
 sky130_fd_sc_hd__nand2_4 _38205_ (.A(_07679_),
    .B(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__nand2_4 _38206_ (.A(_07678_),
    .B(_07681_),
    .Y(_07682_));
 sky130_fd_sc_hd__a21boi_4 _38207_ (.A1(_07478_),
    .A2(_07484_),
    .B1_N(_07480_),
    .Y(_07683_));
 sky130_fd_sc_hd__nand2_4 _38208_ (.A(_07682_),
    .B(_07683_),
    .Y(_07684_));
 sky130_vsdinv _38209_ (.A(_07683_),
    .Y(_07685_));
 sky130_fd_sc_hd__nand3_4 _38210_ (.A(_07678_),
    .B(_07681_),
    .C(_07685_),
    .Y(_07686_));
 sky130_fd_sc_hd__nand2_4 _38211_ (.A(_07684_),
    .B(_07686_),
    .Y(_07687_));
 sky130_vsdinv _38212_ (.A(_07491_),
    .Y(_07688_));
 sky130_fd_sc_hd__a21oi_4 _38213_ (.A1(_07490_),
    .A2(_07495_),
    .B1(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__nand2_4 _38214_ (.A(_07687_),
    .B(_07689_),
    .Y(_07690_));
 sky130_fd_sc_hd__a21o_4 _38215_ (.A1(_07490_),
    .A2(_07495_),
    .B1(_07688_),
    .X(_07691_));
 sky130_fd_sc_hd__nand3_4 _38216_ (.A(_07691_),
    .B(_07686_),
    .C(_07684_),
    .Y(_07692_));
 sky130_fd_sc_hd__nand2_4 _38217_ (.A(_07690_),
    .B(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__nand2_4 _38218_ (.A(_07651_),
    .B(_07693_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand3_4 _38219_ (.A(_07650_),
    .B(_07692_),
    .C(_07690_),
    .Y(_07695_));
 sky130_fd_sc_hd__nand2_4 _38220_ (.A(_07694_),
    .B(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__nand4_4 _38221_ (.A(_07380_),
    .B(_07377_),
    .C(_07569_),
    .D(_07570_),
    .Y(_07697_));
 sky130_fd_sc_hd__nand2_4 _38222_ (.A(_07696_),
    .B(_07697_),
    .Y(_07698_));
 sky130_vsdinv _38223_ (.A(_07697_),
    .Y(_07699_));
 sky130_fd_sc_hd__nand3_4 _38224_ (.A(_07694_),
    .B(_07699_),
    .C(_07695_),
    .Y(_07700_));
 sky130_fd_sc_hd__nand2_4 _38225_ (.A(_07698_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__a21boi_4 _38226_ (.A1(_07462_),
    .A2(_07499_),
    .B1_N(_07501_),
    .Y(_07702_));
 sky130_fd_sc_hd__nand2_4 _38227_ (.A(_07701_),
    .B(_07702_),
    .Y(_07703_));
 sky130_vsdinv _38228_ (.A(_07702_),
    .Y(_07704_));
 sky130_fd_sc_hd__nand3_4 _38229_ (.A(_07698_),
    .B(_07704_),
    .C(_07700_),
    .Y(_07705_));
 sky130_fd_sc_hd__nand2_4 _38230_ (.A(_07703_),
    .B(_07705_),
    .Y(_07706_));
 sky130_fd_sc_hd__nand2_4 _38231_ (.A(_05589_),
    .B(_03546_),
    .Y(_07707_));
 sky130_fd_sc_hd__maj3_4 _38232_ (.A(_07564_),
    .B(_07555_),
    .C(_07558_),
    .X(_07708_));
 sky130_fd_sc_hd__buf_1 _38233_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07709_));
 sky130_fd_sc_hd__buf_1 _38234_ (.A(_07709_),
    .X(_07710_));
 sky130_fd_sc_hd__nand2_4 _38235_ (.A(_06050_),
    .B(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__buf_1 _38236_ (.A(\pcpi_mul.rs2[16] ),
    .X(_07712_));
 sky130_fd_sc_hd__buf_1 _38237_ (.A(_07712_),
    .X(_07713_));
 sky130_fd_sc_hd__nand2_4 _38238_ (.A(_05900_),
    .B(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__nand2_4 _38239_ (.A(_07711_),
    .B(_07714_),
    .Y(_07715_));
 sky130_fd_sc_hd__buf_1 _38240_ (.A(_03539_),
    .X(_07716_));
 sky130_fd_sc_hd__buf_1 _38241_ (.A(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__nand4_4 _38242_ (.A(_06746_),
    .B(_06127_),
    .C(_03536_),
    .D(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__buf_1 _38243_ (.A(\pcpi_mul.rs2[15] ),
    .X(_07719_));
 sky130_fd_sc_hd__buf_1 _38244_ (.A(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__nand2_4 _38245_ (.A(_05916_),
    .B(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__a21bo_4 _38246_ (.A1(_07715_),
    .A2(_07718_),
    .B1_N(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__nand4_4 _38247_ (.A(_05944_),
    .B(_07715_),
    .C(_07718_),
    .D(_07337_),
    .Y(_07723_));
 sky130_fd_sc_hd__nand2_4 _38248_ (.A(_07722_),
    .B(_07723_),
    .Y(_07724_));
 sky130_fd_sc_hd__nor2_4 _38249_ (.A(_07708_),
    .B(_07724_),
    .Y(_07725_));
 sky130_vsdinv _38250_ (.A(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__nand2_4 _38251_ (.A(_07724_),
    .B(_07708_),
    .Y(_07727_));
 sky130_fd_sc_hd__nand3_4 _38252_ (.A(_07565_),
    .B(_07340_),
    .C(_07566_),
    .Y(_07728_));
 sky130_vsdinv _38253_ (.A(_07728_),
    .Y(_07729_));
 sky130_fd_sc_hd__a21o_4 _38254_ (.A1(_07726_),
    .A2(_07727_),
    .B1(_07729_),
    .X(_07730_));
 sky130_fd_sc_hd__nand3_4 _38255_ (.A(_07726_),
    .B(_07729_),
    .C(_07727_),
    .Y(_07731_));
 sky130_fd_sc_hd__a21boi_4 _38256_ (.A1(_07520_),
    .A2(_07528_),
    .B1_N(_07524_),
    .Y(_07732_));
 sky130_fd_sc_hd__buf_1 _38257_ (.A(\pcpi_mul.rs2[14] ),
    .X(_07733_));
 sky130_fd_sc_hd__buf_1 _38258_ (.A(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__nand2_4 _38259_ (.A(_06010_),
    .B(_07734_),
    .Y(_07735_));
 sky130_fd_sc_hd__buf_1 _38260_ (.A(_03268_),
    .X(_07736_));
 sky130_fd_sc_hd__buf_1 _38261_ (.A(_03516_),
    .X(_07737_));
 sky130_fd_sc_hd__nand2_4 _38262_ (.A(_07736_),
    .B(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand2_4 _38263_ (.A(_07735_),
    .B(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__buf_1 _38264_ (.A(_06141_),
    .X(_07740_));
 sky130_fd_sc_hd__buf_1 _38265_ (.A(_07054_),
    .X(_07741_));
 sky130_fd_sc_hd__nand4_4 _38266_ (.A(_07740_),
    .B(_06160_),
    .C(_07518_),
    .D(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__nand2_4 _38267_ (.A(_07739_),
    .B(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__buf_1 _38268_ (.A(_07044_),
    .X(_07744_));
 sky130_fd_sc_hd__nand2_4 _38269_ (.A(_06170_),
    .B(_07744_),
    .Y(_07745_));
 sky130_fd_sc_hd__nand2_4 _38270_ (.A(_07743_),
    .B(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__buf_1 _38271_ (.A(_07045_),
    .X(_07747_));
 sky130_fd_sc_hd__nand4_4 _38272_ (.A(_06171_),
    .B(_07739_),
    .C(_07742_),
    .D(_07747_),
    .Y(_07748_));
 sky130_fd_sc_hd__nand2_4 _38273_ (.A(_07746_),
    .B(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__nor2_4 _38274_ (.A(_07732_),
    .B(_07749_),
    .Y(_07750_));
 sky130_vsdinv _38275_ (.A(_07750_),
    .Y(_07751_));
 sky130_fd_sc_hd__nand2_4 _38276_ (.A(_07749_),
    .B(_07732_),
    .Y(_07752_));
 sky130_fd_sc_hd__buf_1 _38277_ (.A(_06450_),
    .X(_07753_));
 sky130_fd_sc_hd__buf_1 _38278_ (.A(\pcpi_mul.rs2[9] ),
    .X(_07754_));
 sky130_fd_sc_hd__nand2_4 _38279_ (.A(_07753_),
    .B(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__buf_1 _38280_ (.A(_07343_),
    .X(_07756_));
 sky130_fd_sc_hd__nand2_4 _38281_ (.A(_06942_),
    .B(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__buf_1 _38282_ (.A(_06254_),
    .X(_07758_));
 sky130_fd_sc_hd__nand2_4 _38283_ (.A(_07758_),
    .B(_06887_),
    .Y(_07759_));
 sky130_fd_sc_hd__nand2_4 _38284_ (.A(_07757_),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__buf_1 _38285_ (.A(_03279_),
    .X(_07761_));
 sky130_fd_sc_hd__buf_1 _38286_ (.A(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__nand4_4 _38287_ (.A(_06545_),
    .B(_07762_),
    .C(_07347_),
    .D(_07756_),
    .Y(_07763_));
 sky130_fd_sc_hd__nand2_4 _38288_ (.A(_07760_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__xor2_4 _38289_ (.A(_07755_),
    .B(_07764_),
    .X(_07765_));
 sky130_fd_sc_hd__a21o_4 _38290_ (.A1(_07751_),
    .A2(_07752_),
    .B1(_07765_),
    .X(_07766_));
 sky130_fd_sc_hd__nand3_4 _38291_ (.A(_07751_),
    .B(_07765_),
    .C(_07752_),
    .Y(_07767_));
 sky130_fd_sc_hd__and2_4 _38292_ (.A(_07766_),
    .B(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__a21o_4 _38293_ (.A1(_07730_),
    .A2(_07731_),
    .B1(_07768_),
    .X(_07769_));
 sky130_fd_sc_hd__nand4_4 _38294_ (.A(_07730_),
    .B(_07766_),
    .C(_07731_),
    .D(_07767_),
    .Y(_07770_));
 sky130_fd_sc_hd__nand2_4 _38295_ (.A(_07769_),
    .B(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__nand2_4 _38296_ (.A(_07771_),
    .B(_07570_),
    .Y(_07772_));
 sky130_vsdinv _38297_ (.A(_07570_),
    .Y(_07773_));
 sky130_fd_sc_hd__nand3_4 _38298_ (.A(_07769_),
    .B(_07773_),
    .C(_07770_),
    .Y(_07774_));
 sky130_fd_sc_hd__nand2_4 _38299_ (.A(_07772_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__xor2_4 _38300_ (.A(_07707_),
    .B(_07775_),
    .X(_07776_));
 sky130_vsdinv _38301_ (.A(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__nand2_4 _38302_ (.A(_07706_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__nand3_4 _38303_ (.A(_07703_),
    .B(_07776_),
    .C(_07705_),
    .Y(_07779_));
 sky130_fd_sc_hd__buf_1 _38304_ (.A(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__nand2_4 _38305_ (.A(_07778_),
    .B(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__nand2_4 _38306_ (.A(_07781_),
    .B(_07576_),
    .Y(_07782_));
 sky130_vsdinv _38307_ (.A(_07575_),
    .Y(_07783_));
 sky130_fd_sc_hd__nand3_4 _38308_ (.A(_07783_),
    .B(_07780_),
    .C(_07778_),
    .Y(_07784_));
 sky130_fd_sc_hd__nand2_4 _38309_ (.A(_07782_),
    .B(_07784_),
    .Y(_07785_));
 sky130_fd_sc_hd__a21boi_4 _38310_ (.A1(_07455_),
    .A2(_07460_),
    .B1_N(_07456_),
    .Y(_07786_));
 sky130_fd_sc_hd__a21oi_4 _38311_ (.A1(_07515_),
    .A2(_07510_),
    .B1(_07786_),
    .Y(_07787_));
 sky130_vsdinv _38312_ (.A(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__nand3_4 _38313_ (.A(_07515_),
    .B(_07510_),
    .C(_07786_),
    .Y(_07789_));
 sky130_fd_sc_hd__nand2_4 _38314_ (.A(_07788_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__nand2_4 _38315_ (.A(_07785_),
    .B(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__nand4_4 _38316_ (.A(_07788_),
    .B(_07782_),
    .C(_07789_),
    .D(_07784_),
    .Y(_07792_));
 sky130_fd_sc_hd__nand2_4 _38317_ (.A(_07791_),
    .B(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__a21boi_4 _38318_ (.A1(_07578_),
    .A2(_07585_),
    .B1_N(_07580_),
    .Y(_07794_));
 sky130_fd_sc_hd__nand2_4 _38319_ (.A(_07793_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__nand2_4 _38320_ (.A(_07586_),
    .B(_07580_),
    .Y(_07796_));
 sky130_fd_sc_hd__nand3_4 _38321_ (.A(_07796_),
    .B(_07791_),
    .C(_07792_),
    .Y(_07797_));
 sky130_fd_sc_hd__nand2_4 _38322_ (.A(_07795_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__nand4_4 _38323_ (.A(_07331_),
    .B(_07327_),
    .C(_07326_),
    .D(_07582_),
    .Y(_07799_));
 sky130_fd_sc_hd__nand2_4 _38324_ (.A(_07798_),
    .B(_07799_),
    .Y(_07800_));
 sky130_vsdinv _38325_ (.A(_07799_),
    .Y(_07801_));
 sky130_fd_sc_hd__nand3_4 _38326_ (.A(_07795_),
    .B(_07797_),
    .C(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__nand2_4 _38327_ (.A(_07800_),
    .B(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__a21boi_4 _38328_ (.A1(_07589_),
    .A2(_07595_),
    .B1_N(_07591_),
    .Y(_07804_));
 sky130_fd_sc_hd__nand2_4 _38329_ (.A(_07803_),
    .B(_07804_),
    .Y(_07805_));
 sky130_fd_sc_hd__nand2_4 _38330_ (.A(_07596_),
    .B(_07591_),
    .Y(_07806_));
 sky130_fd_sc_hd__nand3_4 _38331_ (.A(_07806_),
    .B(_07800_),
    .C(_07802_),
    .Y(_07807_));
 sky130_fd_sc_hd__and2_4 _38332_ (.A(_07805_),
    .B(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__nand3_4 _38333_ (.A(_07413_),
    .B(_07601_),
    .C(_07600_),
    .Y(_07809_));
 sky130_vsdinv _38334_ (.A(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__nand2_4 _38335_ (.A(_07601_),
    .B(_07411_),
    .Y(_07811_));
 sky130_fd_sc_hd__nand2_4 _38336_ (.A(_07811_),
    .B(_07600_),
    .Y(_07812_));
 sky130_fd_sc_hd__a21boi_4 _38337_ (.A1(_07415_),
    .A2(_07810_),
    .B1_N(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__xnor2_4 _38338_ (.A(_07808_),
    .B(_07813_),
    .Y(_01423_));
 sky130_vsdinv _38339_ (.A(_07755_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21boi_4 _38340_ (.A1(_07760_),
    .A2(_07814_),
    .B1_N(_07763_),
    .Y(_07815_));
 sky130_vsdinv _38341_ (.A(_07815_),
    .Y(_07816_));
 sky130_fd_sc_hd__nand2_4 _38342_ (.A(_06843_),
    .B(_03491_),
    .Y(_07817_));
 sky130_fd_sc_hd__buf_1 _38343_ (.A(\pcpi_mul.rs1[12] ),
    .X(_07818_));
 sky130_fd_sc_hd__buf_1 _38344_ (.A(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__nand2_4 _38345_ (.A(_07819_),
    .B(_06477_),
    .Y(_07820_));
 sky130_fd_sc_hd__nand2_4 _38346_ (.A(_07817_),
    .B(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__buf_1 _38347_ (.A(_06570_),
    .X(_07822_));
 sky130_fd_sc_hd__nand4_4 _38348_ (.A(_07822_),
    .B(_06849_),
    .C(_07467_),
    .D(_06482_),
    .Y(_07823_));
 sky130_fd_sc_hd__buf_1 _38349_ (.A(_06998_),
    .X(_07824_));
 sky130_fd_sc_hd__nand2_4 _38350_ (.A(_07824_),
    .B(_03476_),
    .Y(_07825_));
 sky130_vsdinv _38351_ (.A(_07825_),
    .Y(_07826_));
 sky130_fd_sc_hd__nand3_4 _38352_ (.A(_07821_),
    .B(_07823_),
    .C(_07826_),
    .Y(_07827_));
 sky130_fd_sc_hd__nand2_4 _38353_ (.A(_07821_),
    .B(_07823_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand2_4 _38354_ (.A(_07828_),
    .B(_07825_),
    .Y(_07829_));
 sky130_fd_sc_hd__nand3_4 _38355_ (.A(_07816_),
    .B(_07827_),
    .C(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__nand2_4 _38356_ (.A(_07829_),
    .B(_07827_),
    .Y(_07831_));
 sky130_fd_sc_hd__nand2_4 _38357_ (.A(_07831_),
    .B(_07815_),
    .Y(_07832_));
 sky130_fd_sc_hd__nand2_4 _38358_ (.A(_07830_),
    .B(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__a21boi_4 _38359_ (.A1(_07657_),
    .A2(_07663_),
    .B1_N(_07658_),
    .Y(_07834_));
 sky130_fd_sc_hd__nand2_4 _38360_ (.A(_07833_),
    .B(_07834_),
    .Y(_07835_));
 sky130_vsdinv _38361_ (.A(_07834_),
    .Y(_07836_));
 sky130_fd_sc_hd__nand3_4 _38362_ (.A(_07830_),
    .B(_07832_),
    .C(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__nand2_4 _38363_ (.A(_07835_),
    .B(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__a21oi_4 _38364_ (.A1(_07765_),
    .A2(_07752_),
    .B1(_07750_),
    .Y(_07839_));
 sky130_fd_sc_hd__nand2_4 _38365_ (.A(_07838_),
    .B(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__a21o_4 _38366_ (.A1(_07765_),
    .A2(_07752_),
    .B1(_07750_),
    .X(_07841_));
 sky130_fd_sc_hd__nand3_4 _38367_ (.A(_07841_),
    .B(_07837_),
    .C(_07835_),
    .Y(_07842_));
 sky130_fd_sc_hd__nand2_4 _38368_ (.A(_07840_),
    .B(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__a21boi_4 _38369_ (.A1(_07667_),
    .A2(_07674_),
    .B1_N(_07672_),
    .Y(_07844_));
 sky130_fd_sc_hd__nand2_4 _38370_ (.A(_07843_),
    .B(_07844_),
    .Y(_07845_));
 sky130_vsdinv _38371_ (.A(_07844_),
    .Y(_07846_));
 sky130_fd_sc_hd__nand3_4 _38372_ (.A(_07840_),
    .B(_07842_),
    .C(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand2_4 _38373_ (.A(_07845_),
    .B(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__a21boi_4 _38374_ (.A1(_07685_),
    .A2(_07681_),
    .B1_N(_07678_),
    .Y(_07849_));
 sky130_fd_sc_hd__nand2_4 _38375_ (.A(_07848_),
    .B(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__nand2_4 _38376_ (.A(_07686_),
    .B(_07678_),
    .Y(_07851_));
 sky130_fd_sc_hd__nand3_4 _38377_ (.A(_07851_),
    .B(_07845_),
    .C(_07847_),
    .Y(_07852_));
 sky130_fd_sc_hd__nand2_4 _38378_ (.A(_07850_),
    .B(_07852_),
    .Y(_07853_));
 sky130_vsdinv _38379_ (.A(_07616_),
    .Y(_07854_));
 sky130_fd_sc_hd__a21oi_4 _38380_ (.A1(_07615_),
    .A2(_07636_),
    .B1(_07854_),
    .Y(_07855_));
 sky130_vsdinv _38381_ (.A(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__nand2_4 _38382_ (.A(_07153_),
    .B(_06696_),
    .Y(_07857_));
 sky130_fd_sc_hd__buf_1 _38383_ (.A(_07157_),
    .X(_07858_));
 sky130_fd_sc_hd__nand2_4 _38384_ (.A(_07858_),
    .B(_06427_),
    .Y(_07859_));
 sky130_fd_sc_hd__nand2_4 _38385_ (.A(_07857_),
    .B(_07859_),
    .Y(_07860_));
 sky130_fd_sc_hd__nand4_4 _38386_ (.A(_07153_),
    .B(_07306_),
    .C(_06430_),
    .D(_06432_),
    .Y(_07861_));
 sky130_fd_sc_hd__nand2_4 _38387_ (.A(_07625_),
    .B(_03454_),
    .Y(_07862_));
 sky130_vsdinv _38388_ (.A(_07862_),
    .Y(_07863_));
 sky130_fd_sc_hd__a21o_4 _38389_ (.A1(_07860_),
    .A2(_07861_),
    .B1(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__nand3_4 _38390_ (.A(_07860_),
    .B(_07861_),
    .C(_07863_),
    .Y(_07865_));
 sky130_fd_sc_hd__a21boi_4 _38391_ (.A1(_07607_),
    .A2(_07610_),
    .B1_N(_07608_),
    .Y(_07866_));
 sky130_fd_sc_hd__a21boi_4 _38392_ (.A1(_07864_),
    .A2(_07865_),
    .B1_N(_07866_),
    .Y(_07867_));
 sky130_vsdinv _38393_ (.A(_07867_),
    .Y(_07868_));
 sky130_fd_sc_hd__nand2_4 _38394_ (.A(_07444_),
    .B(_06015_),
    .Y(_07869_));
 sky130_fd_sc_hd__buf_1 _38395_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07870_));
 sky130_fd_sc_hd__buf_1 _38396_ (.A(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__nand2_4 _38397_ (.A(_07871_),
    .B(_06013_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_4 _38398_ (.A(_07869_),
    .B(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__buf_1 _38399_ (.A(_07442_),
    .X(_07874_));
 sky130_fd_sc_hd__buf_1 _38400_ (.A(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__nand4_4 _38401_ (.A(_07875_),
    .B(_03337_),
    .C(_03435_),
    .D(_05939_),
    .Y(_07876_));
 sky130_fd_sc_hd__buf_1 _38402_ (.A(_03340_),
    .X(_07877_));
 sky130_fd_sc_hd__buf_1 _38403_ (.A(_07877_),
    .X(_07878_));
 sky130_fd_sc_hd__nand2_4 _38404_ (.A(_07878_),
    .B(_03419_),
    .Y(_07879_));
 sky130_vsdinv _38405_ (.A(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__a21oi_4 _38406_ (.A1(_07873_),
    .A2(_07876_),
    .B1(_07880_),
    .Y(_07881_));
 sky130_fd_sc_hd__nand3_4 _38407_ (.A(_07873_),
    .B(_07876_),
    .C(_07880_),
    .Y(_07882_));
 sky130_vsdinv _38408_ (.A(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__nor2_4 _38409_ (.A(_07881_),
    .B(_07883_),
    .Y(_07884_));
 sky130_vsdinv _38410_ (.A(_07866_),
    .Y(_07885_));
 sky130_fd_sc_hd__nand3_4 _38411_ (.A(_07885_),
    .B(_07865_),
    .C(_07864_),
    .Y(_07886_));
 sky130_fd_sc_hd__nand3_4 _38412_ (.A(_07868_),
    .B(_07884_),
    .C(_07886_),
    .Y(_07887_));
 sky130_vsdinv _38413_ (.A(_07886_),
    .Y(_07888_));
 sky130_vsdinv _38414_ (.A(_07884_),
    .Y(_07889_));
 sky130_fd_sc_hd__o21ai_4 _38415_ (.A1(_07867_),
    .A2(_07888_),
    .B1(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__nand3_4 _38416_ (.A(_07856_),
    .B(_07887_),
    .C(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__nand2_4 _38417_ (.A(_07890_),
    .B(_07887_),
    .Y(_07892_));
 sky130_fd_sc_hd__nand2_4 _38418_ (.A(_07892_),
    .B(_07855_),
    .Y(_07893_));
 sky130_fd_sc_hd__a21boi_4 _38419_ (.A1(_07623_),
    .A2(_07632_),
    .B1_N(_07628_),
    .Y(_07894_));
 sky130_vsdinv _38420_ (.A(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__a21oi_4 _38421_ (.A1(_07891_),
    .A2(_07893_),
    .B1(_07895_),
    .Y(_07896_));
 sky130_vsdinv _38422_ (.A(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__nand3_4 _38423_ (.A(_07891_),
    .B(_07893_),
    .C(_07895_),
    .Y(_07898_));
 sky130_fd_sc_hd__nand2_4 _38424_ (.A(_07897_),
    .B(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__nand2_4 _38425_ (.A(_07853_),
    .B(_07899_),
    .Y(_07900_));
 sky130_vsdinv _38426_ (.A(_07898_),
    .Y(_07901_));
 sky130_fd_sc_hd__nor2_4 _38427_ (.A(_07896_),
    .B(_07901_),
    .Y(_07902_));
 sky130_fd_sc_hd__nand3_4 _38428_ (.A(_07902_),
    .B(_07852_),
    .C(_07850_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand2_4 _38429_ (.A(_07900_),
    .B(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__nand2_4 _38430_ (.A(_07904_),
    .B(_07774_),
    .Y(_07905_));
 sky130_vsdinv _38431_ (.A(_07774_),
    .Y(_07906_));
 sky130_fd_sc_hd__nand3_4 _38432_ (.A(_07900_),
    .B(_07903_),
    .C(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__nand2_4 _38433_ (.A(_07905_),
    .B(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__a21boi_4 _38434_ (.A1(_07650_),
    .A2(_07690_),
    .B1_N(_07692_),
    .Y(_07909_));
 sky130_fd_sc_hd__nand2_4 _38435_ (.A(_07908_),
    .B(_07909_),
    .Y(_07910_));
 sky130_vsdinv _38436_ (.A(_07909_),
    .Y(_07911_));
 sky130_fd_sc_hd__nand3_4 _38437_ (.A(_07905_),
    .B(_07911_),
    .C(_07907_),
    .Y(_07912_));
 sky130_fd_sc_hd__nand2_4 _38438_ (.A(_07910_),
    .B(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__maj3_4 _38439_ (.A(_07721_),
    .B(_07711_),
    .C(_07714_),
    .X(_07914_));
 sky130_fd_sc_hd__buf_1 _38440_ (.A(_07716_),
    .X(_07915_));
 sky130_fd_sc_hd__nand2_4 _38441_ (.A(_06133_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__buf_1 _38442_ (.A(_03535_),
    .X(_07917_));
 sky130_fd_sc_hd__nand2_4 _38443_ (.A(_06227_),
    .B(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__nand2_4 _38444_ (.A(_07916_),
    .B(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__buf_1 _38445_ (.A(_07713_),
    .X(_07920_));
 sky130_fd_sc_hd__buf_1 _38446_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07921_));
 sky130_fd_sc_hd__buf_1 _38447_ (.A(_07921_),
    .X(_07922_));
 sky130_fd_sc_hd__buf_1 _38448_ (.A(_07922_),
    .X(_07923_));
 sky130_fd_sc_hd__nand4_4 _38449_ (.A(_05901_),
    .B(_05916_),
    .C(_07920_),
    .D(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__nand2_4 _38450_ (.A(_06011_),
    .B(_07563_),
    .Y(_07925_));
 sky130_fd_sc_hd__a21bo_4 _38451_ (.A1(_07919_),
    .A2(_07924_),
    .B1_N(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__nand4_4 _38452_ (.A(_05953_),
    .B(_07919_),
    .C(_07924_),
    .D(_03532_),
    .Y(_07927_));
 sky130_fd_sc_hd__nand2_4 _38453_ (.A(_07926_),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__nor2_4 _38454_ (.A(_07914_),
    .B(_07928_),
    .Y(_07929_));
 sky130_vsdinv _38455_ (.A(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__nand2_4 _38456_ (.A(_07928_),
    .B(_07914_),
    .Y(_07931_));
 sky130_fd_sc_hd__nand3_4 _38457_ (.A(_07930_),
    .B(_07725_),
    .C(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__a21o_4 _38458_ (.A1(_07930_),
    .A2(_07931_),
    .B1(_07725_),
    .X(_07933_));
 sky130_fd_sc_hd__maj3_4 _38459_ (.A(_07745_),
    .B(_07735_),
    .C(_07738_),
    .X(_07934_));
 sky130_fd_sc_hd__nand2_4 _38460_ (.A(_06019_),
    .B(_07353_),
    .Y(_07935_));
 sky130_fd_sc_hd__nand2_4 _38461_ (.A(_06325_),
    .B(_07356_),
    .Y(_07936_));
 sky130_fd_sc_hd__nand2_4 _38462_ (.A(_07935_),
    .B(_07936_),
    .Y(_07937_));
 sky130_fd_sc_hd__buf_1 _38463_ (.A(_06159_),
    .X(_07938_));
 sky130_fd_sc_hd__buf_1 _38464_ (.A(_03271_),
    .X(_07939_));
 sky130_fd_sc_hd__buf_1 _38465_ (.A(_03516_),
    .X(_07940_));
 sky130_fd_sc_hd__buf_1 _38466_ (.A(_07361_),
    .X(_07941_));
 sky130_fd_sc_hd__nand4_4 _38467_ (.A(_07938_),
    .B(_07939_),
    .C(_07940_),
    .D(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__nand2_4 _38468_ (.A(_07937_),
    .B(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_4 _38469_ (.A(_06247_),
    .B(_07366_),
    .Y(_07944_));
 sky130_fd_sc_hd__nand2_4 _38470_ (.A(_07943_),
    .B(_07944_),
    .Y(_07945_));
 sky130_vsdinv _38471_ (.A(_07944_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand3_4 _38472_ (.A(_07937_),
    .B(_07942_),
    .C(_07946_),
    .Y(_07947_));
 sky130_fd_sc_hd__nand2_4 _38473_ (.A(_07945_),
    .B(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__nor2_4 _38474_ (.A(_07934_),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__nand2_4 _38475_ (.A(_07948_),
    .B(_07934_),
    .Y(_07950_));
 sky130_vsdinv _38476_ (.A(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__buf_1 _38477_ (.A(_06566_),
    .X(_07952_));
 sky130_fd_sc_hd__nand2_4 _38478_ (.A(_07952_),
    .B(_07754_),
    .Y(_07953_));
 sky130_vsdinv _38479_ (.A(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__nand2_4 _38480_ (.A(_07762_),
    .B(_06893_),
    .Y(_07955_));
 sky130_fd_sc_hd__buf_1 _38481_ (.A(_07211_),
    .X(_07956_));
 sky130_fd_sc_hd__nand2_4 _38482_ (.A(_07465_),
    .B(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__nand2_4 _38483_ (.A(_07955_),
    .B(_07957_),
    .Y(_07958_));
 sky130_fd_sc_hd__buf_1 _38484_ (.A(_07761_),
    .X(_07959_));
 sky130_fd_sc_hd__nand4_4 _38485_ (.A(_07959_),
    .B(_07465_),
    .C(_07347_),
    .D(_07756_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand2_4 _38486_ (.A(_07958_),
    .B(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__xor2_4 _38487_ (.A(_07954_),
    .B(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__o21ai_4 _38488_ (.A1(_07949_),
    .A2(_07951_),
    .B1(_07962_),
    .Y(_07963_));
 sky130_vsdinv _38489_ (.A(_07949_),
    .Y(_07964_));
 sky130_vsdinv _38490_ (.A(_07962_),
    .Y(_07965_));
 sky130_fd_sc_hd__nand3_4 _38491_ (.A(_07964_),
    .B(_07965_),
    .C(_07950_),
    .Y(_07966_));
 sky130_fd_sc_hd__and2_4 _38492_ (.A(_07963_),
    .B(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__a21o_4 _38493_ (.A1(_07932_),
    .A2(_07933_),
    .B1(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__nand4_4 _38494_ (.A(_07966_),
    .B(_07933_),
    .C(_07963_),
    .D(_07932_),
    .Y(_07969_));
 sky130_fd_sc_hd__nand2_4 _38495_ (.A(_07968_),
    .B(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__nand2_4 _38496_ (.A(_07770_),
    .B(_07731_),
    .Y(_07971_));
 sky130_vsdinv _38497_ (.A(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__nand2_4 _38498_ (.A(_07970_),
    .B(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__nand3_4 _38499_ (.A(_07968_),
    .B(_07971_),
    .C(_07969_),
    .Y(_07974_));
 sky130_fd_sc_hd__buf_1 _38500_ (.A(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__buf_1 _38501_ (.A(_03551_),
    .X(_07976_));
 sky130_fd_sc_hd__buf_1 _38502_ (.A(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__nand2_4 _38503_ (.A(_05895_),
    .B(_07977_),
    .Y(_07978_));
 sky130_fd_sc_hd__buf_1 _38504_ (.A(\pcpi_mul.rs2[18] ),
    .X(_07979_));
 sky130_fd_sc_hd__buf_1 _38505_ (.A(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__nand2_4 _38506_ (.A(_06276_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__xnor2_4 _38507_ (.A(_07978_),
    .B(_07981_),
    .Y(_07982_));
 sky130_vsdinv _38508_ (.A(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__a21oi_4 _38509_ (.A1(_07973_),
    .A2(_07975_),
    .B1(_07983_),
    .Y(_07984_));
 sky130_fd_sc_hd__nand3_4 _38510_ (.A(_07973_),
    .B(_07983_),
    .C(_07974_),
    .Y(_07985_));
 sky130_vsdinv _38511_ (.A(_07985_),
    .Y(_07986_));
 sky130_vsdinv _38512_ (.A(_07707_),
    .Y(_07987_));
 sky130_fd_sc_hd__nand3_4 _38513_ (.A(_07772_),
    .B(_07774_),
    .C(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__o21ai_4 _38514_ (.A1(_07984_),
    .A2(_07986_),
    .B1(_07988_),
    .Y(_07989_));
 sky130_vsdinv _38515_ (.A(_07988_),
    .Y(_07990_));
 sky130_fd_sc_hd__a21o_4 _38516_ (.A1(_07973_),
    .A2(_07975_),
    .B1(_07983_),
    .X(_07991_));
 sky130_fd_sc_hd__nand3_4 _38517_ (.A(_07990_),
    .B(_07985_),
    .C(_07991_),
    .Y(_07992_));
 sky130_fd_sc_hd__nand2_4 _38518_ (.A(_07989_),
    .B(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__nand2_4 _38519_ (.A(_07913_),
    .B(_07993_),
    .Y(_07994_));
 sky130_vsdinv _38520_ (.A(_07993_),
    .Y(_07995_));
 sky130_fd_sc_hd__nand3_4 _38521_ (.A(_07995_),
    .B(_07912_),
    .C(_07910_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_4 _38522_ (.A(_07994_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__nand2_4 _38523_ (.A(_07997_),
    .B(_07780_),
    .Y(_07998_));
 sky130_vsdinv _38524_ (.A(_07779_),
    .Y(_07999_));
 sky130_fd_sc_hd__nand3_4 _38525_ (.A(_07999_),
    .B(_07996_),
    .C(_07994_),
    .Y(_08000_));
 sky130_fd_sc_hd__nand2_4 _38526_ (.A(_07998_),
    .B(_08000_),
    .Y(_08001_));
 sky130_fd_sc_hd__a21boi_4 _38527_ (.A1(_07643_),
    .A2(_07648_),
    .B1_N(_07644_),
    .Y(_08002_));
 sky130_fd_sc_hd__nand2_4 _38528_ (.A(_07705_),
    .B(_07700_),
    .Y(_08003_));
 sky130_fd_sc_hd__xor2_4 _38529_ (.A(_08002_),
    .B(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__nand2_4 _38530_ (.A(_08001_),
    .B(_08004_),
    .Y(_08005_));
 sky130_vsdinv _38531_ (.A(_08004_),
    .Y(_08006_));
 sky130_fd_sc_hd__nand3_4 _38532_ (.A(_08006_),
    .B(_08000_),
    .C(_07998_),
    .Y(_08007_));
 sky130_fd_sc_hd__nand2_4 _38533_ (.A(_08005_),
    .B(_08007_),
    .Y(_08008_));
 sky130_fd_sc_hd__a21boi_4 _38534_ (.A1(_07778_),
    .A2(_07780_),
    .B1_N(_07576_),
    .Y(_08009_));
 sky130_fd_sc_hd__o21ai_4 _38535_ (.A1(_07790_),
    .A2(_08009_),
    .B1(_07784_),
    .Y(_08010_));
 sky130_vsdinv _38536_ (.A(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__nand2_4 _38537_ (.A(_08008_),
    .B(_08011_),
    .Y(_08012_));
 sky130_fd_sc_hd__nand3_4 _38538_ (.A(_08010_),
    .B(_08005_),
    .C(_08007_),
    .Y(_08013_));
 sky130_fd_sc_hd__nand2_4 _38539_ (.A(_08012_),
    .B(_08013_),
    .Y(_08014_));
 sky130_fd_sc_hd__nand2_4 _38540_ (.A(_08014_),
    .B(_07788_),
    .Y(_08015_));
 sky130_fd_sc_hd__nand3_4 _38541_ (.A(_08012_),
    .B(_07787_),
    .C(_08013_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand2_4 _38542_ (.A(_08015_),
    .B(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__a21boi_4 _38543_ (.A1(_07795_),
    .A2(_07801_),
    .B1_N(_07797_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand2_4 _38544_ (.A(_08017_),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand2_4 _38545_ (.A(_07802_),
    .B(_07797_),
    .Y(_08020_));
 sky130_fd_sc_hd__nand3_4 _38546_ (.A(_08020_),
    .B(_08016_),
    .C(_08015_),
    .Y(_08021_));
 sky130_fd_sc_hd__and2_4 _38547_ (.A(_08019_),
    .B(_08021_),
    .X(_08022_));
 sky130_fd_sc_hd__nand2_4 _38548_ (.A(_07415_),
    .B(_07810_),
    .Y(_08023_));
 sky130_fd_sc_hd__a21bo_4 _38549_ (.A1(_08023_),
    .A2(_07812_),
    .B1_N(_07808_),
    .X(_08024_));
 sky130_fd_sc_hd__nand2_4 _38550_ (.A(_08024_),
    .B(_07807_),
    .Y(_08025_));
 sky130_fd_sc_hd__xor2_4 _38551_ (.A(_08022_),
    .B(_08025_),
    .X(_01424_));
 sky130_fd_sc_hd__buf_1 _38552_ (.A(_03317_),
    .X(_08026_));
 sky130_fd_sc_hd__nand2_4 _38553_ (.A(_08026_),
    .B(_06431_),
    .Y(_08027_));
 sky130_fd_sc_hd__buf_1 _38554_ (.A(_05962_),
    .X(_08028_));
 sky130_fd_sc_hd__nand2_4 _38555_ (.A(_07624_),
    .B(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__nand2_4 _38556_ (.A(_08027_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__nand4_4 _38557_ (.A(_07432_),
    .B(_07620_),
    .C(_06059_),
    .D(_06431_),
    .Y(_08031_));
 sky130_fd_sc_hd__buf_1 _38558_ (.A(_03331_),
    .X(_08032_));
 sky130_fd_sc_hd__nand2_4 _38559_ (.A(_08032_),
    .B(_05967_),
    .Y(_08033_));
 sky130_vsdinv _38560_ (.A(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__a21o_4 _38561_ (.A1(_08030_),
    .A2(_08031_),
    .B1(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__nand3_4 _38562_ (.A(_08030_),
    .B(_08031_),
    .C(_08034_),
    .Y(_08036_));
 sky130_fd_sc_hd__a21boi_4 _38563_ (.A1(_07860_),
    .A2(_07863_),
    .B1_N(_07861_),
    .Y(_08037_));
 sky130_fd_sc_hd__a21boi_4 _38564_ (.A1(_08035_),
    .A2(_08036_),
    .B1_N(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__nand2_4 _38565_ (.A(_08035_),
    .B(_08036_),
    .Y(_08039_));
 sky130_fd_sc_hd__nor2_4 _38566_ (.A(_08037_),
    .B(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__nor2_4 _38567_ (.A(_08038_),
    .B(_08040_),
    .Y(_08041_));
 sky130_fd_sc_hd__buf_1 _38568_ (.A(_07870_),
    .X(_08042_));
 sky130_fd_sc_hd__buf_1 _38569_ (.A(_03442_),
    .X(_08043_));
 sky130_fd_sc_hd__nand2_4 _38570_ (.A(_08042_),
    .B(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__buf_1 _38571_ (.A(\pcpi_mul.rs1[19] ),
    .X(_08045_));
 sky130_fd_sc_hd__buf_1 _38572_ (.A(_08045_),
    .X(_08046_));
 sky130_fd_sc_hd__buf_1 _38573_ (.A(_06012_),
    .X(_08047_));
 sky130_fd_sc_hd__nand2_4 _38574_ (.A(_08046_),
    .B(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__nand2_4 _38575_ (.A(_08044_),
    .B(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__buf_1 _38576_ (.A(\pcpi_mul.rs1[18] ),
    .X(_08050_));
 sky130_fd_sc_hd__buf_1 _38577_ (.A(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__buf_1 _38578_ (.A(_07877_),
    .X(_08052_));
 sky130_fd_sc_hd__nand4_4 _38579_ (.A(_08051_),
    .B(_08052_),
    .C(_07440_),
    .D(_03443_),
    .Y(_08053_));
 sky130_fd_sc_hd__buf_1 _38580_ (.A(\pcpi_mul.rs1[20] ),
    .X(_08054_));
 sky130_fd_sc_hd__buf_1 _38581_ (.A(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__buf_1 _38582_ (.A(_08055_),
    .X(_08056_));
 sky130_fd_sc_hd__nand2_4 _38583_ (.A(_08056_),
    .B(_03419_),
    .Y(_08057_));
 sky130_vsdinv _38584_ (.A(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__a21o_4 _38585_ (.A1(_08049_),
    .A2(_08053_),
    .B1(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__nand3_4 _38586_ (.A(_08049_),
    .B(_08053_),
    .C(_08058_),
    .Y(_08060_));
 sky130_fd_sc_hd__and2_4 _38587_ (.A(_08059_),
    .B(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__nand2_4 _38588_ (.A(_08041_),
    .B(_08061_),
    .Y(_08062_));
 sky130_vsdinv _38589_ (.A(_08061_),
    .Y(_08063_));
 sky130_fd_sc_hd__o21ai_4 _38590_ (.A1(_08038_),
    .A2(_08040_),
    .B1(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__o21a_4 _38591_ (.A1(_07867_),
    .A2(_07889_),
    .B1(_07886_),
    .X(_08065_));
 sky130_vsdinv _38592_ (.A(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__a21o_4 _38593_ (.A1(_08062_),
    .A2(_08064_),
    .B1(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__a21boi_4 _38594_ (.A1(_07873_),
    .A2(_07880_),
    .B1_N(_07876_),
    .Y(_08068_));
 sky130_vsdinv _38595_ (.A(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__nand3_4 _38596_ (.A(_08066_),
    .B(_08064_),
    .C(_08062_),
    .Y(_08070_));
 sky130_fd_sc_hd__nand3_4 _38597_ (.A(_08067_),
    .B(_08069_),
    .C(_08070_),
    .Y(_08071_));
 sky130_vsdinv _38598_ (.A(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21oi_4 _38599_ (.A1(_08067_),
    .A2(_08070_),
    .B1(_08069_),
    .Y(_08073_));
 sky130_fd_sc_hd__a21boi_4 _38600_ (.A1(_07840_),
    .A2(_07846_),
    .B1_N(_07842_),
    .Y(_08074_));
 sky130_vsdinv _38601_ (.A(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__a21boi_4 _38602_ (.A1(_07958_),
    .A2(_07954_),
    .B1_N(_07960_),
    .Y(_08076_));
 sky130_vsdinv _38603_ (.A(_08076_),
    .Y(_08077_));
 sky130_fd_sc_hd__nand2_4 _38604_ (.A(_07819_),
    .B(_06788_),
    .Y(_08078_));
 sky130_fd_sc_hd__nand2_4 _38605_ (.A(_07824_),
    .B(_06946_),
    .Y(_08079_));
 sky130_fd_sc_hd__nand2_4 _38606_ (.A(_08078_),
    .B(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__buf_1 _38607_ (.A(\pcpi_mul.rs2[8] ),
    .X(_08081_));
 sky130_fd_sc_hd__buf_1 _38608_ (.A(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__nand4_4 _38609_ (.A(_07660_),
    .B(_07150_),
    .C(_07096_),
    .D(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__nand2_4 _38610_ (.A(_07298_),
    .B(_03476_),
    .Y(_08084_));
 sky130_vsdinv _38611_ (.A(_08084_),
    .Y(_08085_));
 sky130_fd_sc_hd__nand3_4 _38612_ (.A(_08080_),
    .B(_08083_),
    .C(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__nand2_4 _38613_ (.A(_08080_),
    .B(_08083_),
    .Y(_08087_));
 sky130_fd_sc_hd__nand2_4 _38614_ (.A(_08087_),
    .B(_08084_),
    .Y(_08088_));
 sky130_fd_sc_hd__nand3_4 _38615_ (.A(_08077_),
    .B(_08086_),
    .C(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__nand2_4 _38616_ (.A(_08088_),
    .B(_08086_),
    .Y(_08090_));
 sky130_fd_sc_hd__nand2_4 _38617_ (.A(_08090_),
    .B(_08076_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand2_4 _38618_ (.A(_08089_),
    .B(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__a21boi_4 _38619_ (.A1(_07821_),
    .A2(_07826_),
    .B1_N(_07823_),
    .Y(_08093_));
 sky130_fd_sc_hd__nand2_4 _38620_ (.A(_08092_),
    .B(_08093_),
    .Y(_08094_));
 sky130_vsdinv _38621_ (.A(_08093_),
    .Y(_08095_));
 sky130_fd_sc_hd__nand3_4 _38622_ (.A(_08089_),
    .B(_08091_),
    .C(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__nand2_4 _38623_ (.A(_08094_),
    .B(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__a21oi_4 _38624_ (.A1(_07965_),
    .A2(_07950_),
    .B1(_07949_),
    .Y(_08098_));
 sky130_fd_sc_hd__nand2_4 _38625_ (.A(_08097_),
    .B(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__o21ai_4 _38626_ (.A1(_07962_),
    .A2(_07951_),
    .B1(_07964_),
    .Y(_08100_));
 sky130_fd_sc_hd__nand3_4 _38627_ (.A(_08100_),
    .B(_08096_),
    .C(_08094_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand2_4 _38628_ (.A(_08099_),
    .B(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__a21boi_4 _38629_ (.A1(_07832_),
    .A2(_07836_),
    .B1_N(_07830_),
    .Y(_08103_));
 sky130_fd_sc_hd__nand2_4 _38630_ (.A(_08102_),
    .B(_08103_),
    .Y(_08104_));
 sky130_vsdinv _38631_ (.A(_08103_),
    .Y(_08105_));
 sky130_fd_sc_hd__nand3_4 _38632_ (.A(_08099_),
    .B(_08101_),
    .C(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__nand3_4 _38633_ (.A(_08075_),
    .B(_08104_),
    .C(_08106_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand2_4 _38634_ (.A(_08104_),
    .B(_08106_),
    .Y(_08108_));
 sky130_fd_sc_hd__nand2_4 _38635_ (.A(_08108_),
    .B(_08074_),
    .Y(_08109_));
 sky130_fd_sc_hd__nand2_4 _38636_ (.A(_08107_),
    .B(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__o21ai_4 _38637_ (.A1(_08072_),
    .A2(_08073_),
    .B1(_08110_),
    .Y(_08111_));
 sky130_vsdinv _38638_ (.A(_08073_),
    .Y(_08112_));
 sky130_fd_sc_hd__nand4_4 _38639_ (.A(_08071_),
    .B(_08112_),
    .C(_08107_),
    .D(_08109_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand2_4 _38640_ (.A(_08111_),
    .B(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_4 _38641_ (.A(_08114_),
    .B(_07975_),
    .Y(_08115_));
 sky130_vsdinv _38642_ (.A(_07975_),
    .Y(_08116_));
 sky130_fd_sc_hd__nand3_4 _38643_ (.A(_08111_),
    .B(_08113_),
    .C(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__nand2_4 _38644_ (.A(_08115_),
    .B(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__a21boi_4 _38645_ (.A1(_07902_),
    .A2(_07850_),
    .B1_N(_07852_),
    .Y(_08119_));
 sky130_fd_sc_hd__nand2_4 _38646_ (.A(_08118_),
    .B(_08119_),
    .Y(_08120_));
 sky130_vsdinv _38647_ (.A(_08119_),
    .Y(_08121_));
 sky130_fd_sc_hd__nand3_4 _38648_ (.A(_08115_),
    .B(_08121_),
    .C(_08117_),
    .Y(_08122_));
 sky130_fd_sc_hd__nand2_4 _38649_ (.A(_08120_),
    .B(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__buf_1 _38650_ (.A(\pcpi_mul.rs2[17] ),
    .X(_08124_));
 sky130_fd_sc_hd__buf_1 _38651_ (.A(_08124_),
    .X(_08125_));
 sky130_fd_sc_hd__nand2_4 _38652_ (.A(_06008_),
    .B(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__buf_1 _38653_ (.A(\pcpi_mul.rs2[16] ),
    .X(_08127_));
 sky130_fd_sc_hd__buf_1 _38654_ (.A(_08127_),
    .X(_08128_));
 sky130_fd_sc_hd__nand2_4 _38655_ (.A(_06142_),
    .B(_08128_),
    .Y(_08129_));
 sky130_fd_sc_hd__nand2_4 _38656_ (.A(_08126_),
    .B(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__nand4_4 _38657_ (.A(_06227_),
    .B(_06223_),
    .C(_07917_),
    .D(_07915_),
    .Y(_08131_));
 sky130_fd_sc_hd__buf_1 _38658_ (.A(_07719_),
    .X(_08132_));
 sky130_fd_sc_hd__nand2_4 _38659_ (.A(_07208_),
    .B(_08132_),
    .Y(_08133_));
 sky130_vsdinv _38660_ (.A(_08133_),
    .Y(_08134_));
 sky130_fd_sc_hd__a21o_4 _38661_ (.A1(_08130_),
    .A2(_08131_),
    .B1(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__nand3_4 _38662_ (.A(_08130_),
    .B(_08131_),
    .C(_08134_),
    .Y(_08136_));
 sky130_fd_sc_hd__nor2_4 _38663_ (.A(_07978_),
    .B(_07981_),
    .Y(_08137_));
 sky130_fd_sc_hd__a21o_4 _38664_ (.A1(_08135_),
    .A2(_08136_),
    .B1(_08137_),
    .X(_08138_));
 sky130_fd_sc_hd__nand3_4 _38665_ (.A(_08135_),
    .B(_08137_),
    .C(_08136_),
    .Y(_08139_));
 sky130_fd_sc_hd__nand2_4 _38666_ (.A(_08138_),
    .B(_08139_),
    .Y(_08140_));
 sky130_fd_sc_hd__maj3_4 _38667_ (.A(_07925_),
    .B(_07916_),
    .C(_07918_),
    .X(_08141_));
 sky130_fd_sc_hd__nand2_4 _38668_ (.A(_08140_),
    .B(_08141_),
    .Y(_08142_));
 sky130_vsdinv _38669_ (.A(_08141_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand3_4 _38670_ (.A(_08138_),
    .B(_08143_),
    .C(_08139_),
    .Y(_08144_));
 sky130_fd_sc_hd__a21oi_4 _38671_ (.A1(_08142_),
    .A2(_08144_),
    .B1(_07929_),
    .Y(_08145_));
 sky130_fd_sc_hd__nand3_4 _38672_ (.A(_08142_),
    .B(_07929_),
    .C(_08144_),
    .Y(_08146_));
 sky130_vsdinv _38673_ (.A(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__nand2_4 _38674_ (.A(_06084_),
    .B(_03525_),
    .Y(_08148_));
 sky130_fd_sc_hd__nand2_4 _38675_ (.A(_03275_),
    .B(_07521_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand2_4 _38676_ (.A(_08148_),
    .B(_08149_),
    .Y(_08150_));
 sky130_fd_sc_hd__nand4_4 _38677_ (.A(_07939_),
    .B(_06251_),
    .C(_07737_),
    .D(_07734_),
    .Y(_08151_));
 sky130_fd_sc_hd__nand2_4 _38678_ (.A(_06342_),
    .B(_07044_),
    .Y(_08152_));
 sky130_vsdinv _38679_ (.A(_08152_),
    .Y(_08153_));
 sky130_fd_sc_hd__nand3_4 _38680_ (.A(_08150_),
    .B(_08151_),
    .C(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__nand2_4 _38681_ (.A(_08150_),
    .B(_08151_),
    .Y(_08155_));
 sky130_fd_sc_hd__nand2_4 _38682_ (.A(_08155_),
    .B(_08152_),
    .Y(_08156_));
 sky130_fd_sc_hd__a21boi_4 _38683_ (.A1(_07937_),
    .A2(_07946_),
    .B1_N(_07942_),
    .Y(_08157_));
 sky130_fd_sc_hd__a21boi_4 _38684_ (.A1(_08154_),
    .A2(_08156_),
    .B1_N(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__nand2_4 _38685_ (.A(_08156_),
    .B(_08154_),
    .Y(_08159_));
 sky130_fd_sc_hd__nor2_4 _38686_ (.A(_08157_),
    .B(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand2_4 _38687_ (.A(_03298_),
    .B(_07204_),
    .Y(_08161_));
 sky130_fd_sc_hd__buf_1 _38688_ (.A(_03504_),
    .X(_08162_));
 sky130_fd_sc_hd__nand2_4 _38689_ (.A(_06349_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__buf_1 _38690_ (.A(_03499_),
    .X(_08164_));
 sky130_fd_sc_hd__nand2_4 _38691_ (.A(_06832_),
    .B(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__nand2_4 _38692_ (.A(_08163_),
    .B(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__buf_1 _38693_ (.A(_03289_),
    .X(_08167_));
 sky130_fd_sc_hd__buf_1 _38694_ (.A(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__buf_1 _38695_ (.A(_06832_),
    .X(_08169_));
 sky130_fd_sc_hd__nand4_4 _38696_ (.A(_08168_),
    .B(_08169_),
    .C(_06743_),
    .D(_07668_),
    .Y(_08170_));
 sky130_fd_sc_hd__nand2_4 _38697_ (.A(_08166_),
    .B(_08170_),
    .Y(_08171_));
 sky130_fd_sc_hd__xor2_4 _38698_ (.A(_08161_),
    .B(_08171_),
    .X(_08172_));
 sky130_vsdinv _38699_ (.A(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__o21ai_4 _38700_ (.A1(_08158_),
    .A2(_08160_),
    .B1(_08173_),
    .Y(_08174_));
 sky130_vsdinv _38701_ (.A(_08160_),
    .Y(_08175_));
 sky130_vsdinv _38702_ (.A(_08158_),
    .Y(_08176_));
 sky130_fd_sc_hd__nand3_4 _38703_ (.A(_08175_),
    .B(_08176_),
    .C(_08172_),
    .Y(_08177_));
 sky130_fd_sc_hd__nand2_4 _38704_ (.A(_08174_),
    .B(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__o21ai_4 _38705_ (.A1(_08145_),
    .A2(_08147_),
    .B1(_08178_),
    .Y(_08179_));
 sky130_vsdinv _38706_ (.A(_08145_),
    .Y(_08180_));
 sky130_vsdinv _38707_ (.A(_08178_),
    .Y(_08181_));
 sky130_fd_sc_hd__nand3_4 _38708_ (.A(_08180_),
    .B(_08181_),
    .C(_08146_),
    .Y(_08182_));
 sky130_fd_sc_hd__nand2_4 _38709_ (.A(_08179_),
    .B(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__a21boi_4 _38710_ (.A1(_07967_),
    .A2(_07933_),
    .B1_N(_07932_),
    .Y(_08184_));
 sky130_fd_sc_hd__nand2_4 _38711_ (.A(_08183_),
    .B(_08184_),
    .Y(_08185_));
 sky130_vsdinv _38712_ (.A(_08184_),
    .Y(_08186_));
 sky130_fd_sc_hd__nand3_4 _38713_ (.A(_08186_),
    .B(_08179_),
    .C(_08182_),
    .Y(_08187_));
 sky130_fd_sc_hd__nand2_4 _38714_ (.A(_08185_),
    .B(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__nand2_4 _38715_ (.A(_06381_),
    .B(_03545_),
    .Y(_08189_));
 sky130_fd_sc_hd__buf_1 _38716_ (.A(\pcpi_mul.rs2[19] ),
    .X(_08190_));
 sky130_fd_sc_hd__buf_1 _38717_ (.A(_08190_),
    .X(_08191_));
 sky130_fd_sc_hd__nand2_4 _38718_ (.A(_05885_),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__buf_1 _38719_ (.A(\pcpi_mul.rs2[20] ),
    .X(_08193_));
 sky130_fd_sc_hd__buf_1 _38720_ (.A(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__nand2_4 _38721_ (.A(_05961_),
    .B(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__nand2_4 _38722_ (.A(_08192_),
    .B(_08195_),
    .Y(_08196_));
 sky130_fd_sc_hd__buf_1 _38723_ (.A(\pcpi_mul.rs2[20] ),
    .X(_08197_));
 sky130_fd_sc_hd__buf_1 _38724_ (.A(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__nand4_4 _38725_ (.A(_06634_),
    .B(_07048_),
    .C(_08191_),
    .D(_08198_),
    .Y(_08199_));
 sky130_fd_sc_hd__nand2_4 _38726_ (.A(_08196_),
    .B(_08199_),
    .Y(_08200_));
 sky130_fd_sc_hd__xor2_4 _38727_ (.A(_08189_),
    .B(_08200_),
    .X(_08201_));
 sky130_vsdinv _38728_ (.A(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_4 _38729_ (.A(_08188_),
    .B(_08202_),
    .Y(_08203_));
 sky130_fd_sc_hd__nand3_4 _38730_ (.A(_08185_),
    .B(_08201_),
    .C(_08187_),
    .Y(_08204_));
 sky130_fd_sc_hd__a21oi_4 _38731_ (.A1(_08203_),
    .A2(_08204_),
    .B1(_07986_),
    .Y(_08205_));
 sky130_fd_sc_hd__nand3_4 _38732_ (.A(_08203_),
    .B(_07986_),
    .C(_08204_),
    .Y(_08206_));
 sky130_vsdinv _38733_ (.A(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__nor2_4 _38734_ (.A(_08205_),
    .B(_08207_),
    .Y(_08208_));
 sky130_vsdinv _38735_ (.A(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand2_4 _38736_ (.A(_08123_),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__nand3_4 _38737_ (.A(_08120_),
    .B(_08208_),
    .C(_08122_),
    .Y(_08211_));
 sky130_fd_sc_hd__nand2_4 _38738_ (.A(_07996_),
    .B(_07992_),
    .Y(_08212_));
 sky130_fd_sc_hd__a21oi_4 _38739_ (.A1(_08210_),
    .A2(_08211_),
    .B1(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__nand3_4 _38740_ (.A(_08212_),
    .B(_08210_),
    .C(_08211_),
    .Y(_08214_));
 sky130_vsdinv _38741_ (.A(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__a21boi_4 _38742_ (.A1(_07893_),
    .A2(_07895_),
    .B1_N(_07891_),
    .Y(_08216_));
 sky130_fd_sc_hd__a21boi_4 _38743_ (.A1(_07905_),
    .A2(_07911_),
    .B1_N(_07907_),
    .Y(_08217_));
 sky130_fd_sc_hd__xnor2_4 _38744_ (.A(_08216_),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__o21ai_4 _38745_ (.A1(_08213_),
    .A2(_08215_),
    .B1(_08218_),
    .Y(_08219_));
 sky130_fd_sc_hd__nand2_4 _38746_ (.A(_08210_),
    .B(_08211_),
    .Y(_08220_));
 sky130_vsdinv _38747_ (.A(_08212_),
    .Y(_08221_));
 sky130_fd_sc_hd__nand2_4 _38748_ (.A(_08220_),
    .B(_08221_),
    .Y(_08222_));
 sky130_vsdinv _38749_ (.A(_08218_),
    .Y(_08223_));
 sky130_fd_sc_hd__nand3_4 _38750_ (.A(_08222_),
    .B(_08223_),
    .C(_08214_),
    .Y(_08224_));
 sky130_fd_sc_hd__nand2_4 _38751_ (.A(_08219_),
    .B(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__a21boi_4 _38752_ (.A1(_08006_),
    .A2(_07998_),
    .B1_N(_08000_),
    .Y(_08226_));
 sky130_fd_sc_hd__nand2_4 _38753_ (.A(_08225_),
    .B(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__nand2_4 _38754_ (.A(_08007_),
    .B(_08000_),
    .Y(_08228_));
 sky130_fd_sc_hd__nand3_4 _38755_ (.A(_08228_),
    .B(_08224_),
    .C(_08219_),
    .Y(_08229_));
 sky130_fd_sc_hd__nand2_4 _38756_ (.A(_08227_),
    .B(_08229_),
    .Y(_08230_));
 sky130_fd_sc_hd__a21oi_4 _38757_ (.A1(_07705_),
    .A2(_07700_),
    .B1(_08002_),
    .Y(_08231_));
 sky130_vsdinv _38758_ (.A(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__nand2_4 _38759_ (.A(_08230_),
    .B(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand3_4 _38760_ (.A(_08227_),
    .B(_08229_),
    .C(_08231_),
    .Y(_08234_));
 sky130_fd_sc_hd__nand2_4 _38761_ (.A(_08233_),
    .B(_08234_),
    .Y(_08235_));
 sky130_fd_sc_hd__nand2_4 _38762_ (.A(_08016_),
    .B(_08013_),
    .Y(_08236_));
 sky130_vsdinv _38763_ (.A(_08236_),
    .Y(_08237_));
 sky130_fd_sc_hd__nand2_4 _38764_ (.A(_08235_),
    .B(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__nand3_4 _38765_ (.A(_08233_),
    .B(_08236_),
    .C(_08234_),
    .Y(_08239_));
 sky130_fd_sc_hd__and2_4 _38766_ (.A(_08238_),
    .B(_08239_),
    .X(_08240_));
 sky130_vsdinv _38767_ (.A(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__nand4_4 _38768_ (.A(_07807_),
    .B(_07805_),
    .C(_08019_),
    .D(_08021_),
    .Y(_08242_));
 sky130_fd_sc_hd__nor2_4 _38769_ (.A(_08242_),
    .B(_07809_),
    .Y(_08243_));
 sky130_vsdinv _38770_ (.A(_07807_),
    .Y(_08244_));
 sky130_fd_sc_hd__a21boi_4 _38771_ (.A1(_08244_),
    .A2(_08019_),
    .B1_N(_08021_),
    .Y(_08245_));
 sky130_fd_sc_hd__o21ai_4 _38772_ (.A1(_07812_),
    .A2(_08242_),
    .B1(_08245_),
    .Y(_08246_));
 sky130_fd_sc_hd__a21oi_4 _38773_ (.A1(_07414_),
    .A2(_08243_),
    .B1(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__xor2_4 _38774_ (.A(_08241_),
    .B(_08247_),
    .X(_01425_));
 sky130_fd_sc_hd__nand2_4 _38775_ (.A(_08211_),
    .B(_08206_),
    .Y(_08248_));
 sky130_vsdinv _38776_ (.A(_08248_),
    .Y(_08249_));
 sky130_fd_sc_hd__a21boi_4 _38777_ (.A1(_08099_),
    .A2(_08105_),
    .B1_N(_08101_),
    .Y(_08250_));
 sky130_vsdinv _38778_ (.A(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__o21ai_4 _38779_ (.A1(_08158_),
    .A2(_08173_),
    .B1(_08175_),
    .Y(_08252_));
 sky130_vsdinv _38780_ (.A(_08161_),
    .Y(_08253_));
 sky130_fd_sc_hd__nor2_4 _38781_ (.A(_08163_),
    .B(_08165_),
    .Y(_08254_));
 sky130_fd_sc_hd__a21o_4 _38782_ (.A1(_08166_),
    .A2(_08253_),
    .B1(_08254_),
    .X(_08255_));
 sky130_vsdinv _38783_ (.A(_08255_),
    .Y(_08256_));
 sky130_fd_sc_hd__buf_1 _38784_ (.A(_06592_),
    .X(_08257_));
 sky130_fd_sc_hd__nand2_4 _38785_ (.A(_07146_),
    .B(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__buf_1 _38786_ (.A(_06598_),
    .X(_08259_));
 sky130_fd_sc_hd__nand2_4 _38787_ (.A(_07298_),
    .B(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__nand2_4 _38788_ (.A(_08258_),
    .B(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__nand4_4 _38789_ (.A(_06852_),
    .B(_07152_),
    .C(_06376_),
    .D(_03491_),
    .Y(_08262_));
 sky130_fd_sc_hd__nand2_4 _38790_ (.A(_08261_),
    .B(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__nand2_4 _38791_ (.A(_07301_),
    .B(_06796_),
    .Y(_08264_));
 sky130_fd_sc_hd__nand2_4 _38792_ (.A(_08263_),
    .B(_08264_),
    .Y(_08265_));
 sky130_vsdinv _38793_ (.A(_08264_),
    .Y(_08266_));
 sky130_fd_sc_hd__nand3_4 _38794_ (.A(_08261_),
    .B(_08262_),
    .C(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__nand2_4 _38795_ (.A(_08265_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand2_4 _38796_ (.A(_08256_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__a21boi_4 _38797_ (.A1(_08080_),
    .A2(_08085_),
    .B1_N(_08083_),
    .Y(_08270_));
 sky130_vsdinv _38798_ (.A(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__nand3_4 _38799_ (.A(_08255_),
    .B(_08267_),
    .C(_08265_),
    .Y(_08272_));
 sky130_fd_sc_hd__nand3_4 _38800_ (.A(_08269_),
    .B(_08271_),
    .C(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__nand2_4 _38801_ (.A(_08269_),
    .B(_08272_),
    .Y(_08274_));
 sky130_fd_sc_hd__nand2_4 _38802_ (.A(_08274_),
    .B(_08270_),
    .Y(_08275_));
 sky130_fd_sc_hd__nand3_4 _38803_ (.A(_08252_),
    .B(_08273_),
    .C(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__nand2_4 _38804_ (.A(_08275_),
    .B(_08273_),
    .Y(_08277_));
 sky130_fd_sc_hd__a21oi_4 _38805_ (.A1(_08176_),
    .A2(_08172_),
    .B1(_08160_),
    .Y(_08278_));
 sky130_fd_sc_hd__nand2_4 _38806_ (.A(_08277_),
    .B(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__a21boi_4 _38807_ (.A1(_08091_),
    .A2(_08095_),
    .B1_N(_08089_),
    .Y(_08280_));
 sky130_vsdinv _38808_ (.A(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__nand3_4 _38809_ (.A(_08276_),
    .B(_08279_),
    .C(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__nand2_4 _38810_ (.A(_08276_),
    .B(_08279_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand2_4 _38811_ (.A(_08283_),
    .B(_08280_),
    .Y(_08284_));
 sky130_fd_sc_hd__nand3_4 _38812_ (.A(_08251_),
    .B(_08282_),
    .C(_08284_),
    .Y(_08285_));
 sky130_fd_sc_hd__nand2_4 _38813_ (.A(_08284_),
    .B(_08282_),
    .Y(_08286_));
 sky130_fd_sc_hd__nand2_4 _38814_ (.A(_08286_),
    .B(_08250_),
    .Y(_08287_));
 sky130_fd_sc_hd__nand2_4 _38815_ (.A(_08285_),
    .B(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__buf_1 _38816_ (.A(_03323_),
    .X(_08289_));
 sky130_fd_sc_hd__nand2_4 _38817_ (.A(_08289_),
    .B(_06137_),
    .Y(_08290_));
 sky130_fd_sc_hd__buf_1 _38818_ (.A(_07442_),
    .X(_08291_));
 sky130_fd_sc_hd__nand2_4 _38819_ (.A(_08291_),
    .B(_03464_),
    .Y(_08292_));
 sky130_fd_sc_hd__nand2_4 _38820_ (.A(_08290_),
    .B(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__buf_1 _38821_ (.A(_03323_),
    .X(_08294_));
 sky130_fd_sc_hd__nand4_4 _38822_ (.A(_08294_),
    .B(_07874_),
    .C(_06135_),
    .D(_06137_),
    .Y(_08295_));
 sky130_fd_sc_hd__nand2_4 _38823_ (.A(_07629_),
    .B(_06231_),
    .Y(_08296_));
 sky130_vsdinv _38824_ (.A(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__a21o_4 _38825_ (.A1(_08293_),
    .A2(_08295_),
    .B1(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__nand3_4 _38826_ (.A(_08293_),
    .B(_08295_),
    .C(_08297_),
    .Y(_08299_));
 sky130_fd_sc_hd__a21boi_4 _38827_ (.A1(_08030_),
    .A2(_08034_),
    .B1_N(_08031_),
    .Y(_08300_));
 sky130_fd_sc_hd__a21boi_4 _38828_ (.A1(_08298_),
    .A2(_08299_),
    .B1_N(_08300_),
    .Y(_08301_));
 sky130_vsdinv _38829_ (.A(_08300_),
    .Y(_08302_));
 sky130_fd_sc_hd__nand3_4 _38830_ (.A(_08302_),
    .B(_08299_),
    .C(_08298_),
    .Y(_08303_));
 sky130_vsdinv _38831_ (.A(_08303_),
    .Y(_08304_));
 sky130_fd_sc_hd__nand2_4 _38832_ (.A(_03342_),
    .B(_05910_),
    .Y(_08305_));
 sky130_fd_sc_hd__o21ai_4 _38833_ (.A1(_03348_),
    .A2(_07144_),
    .B1(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__buf_1 _38834_ (.A(_08046_),
    .X(_08307_));
 sky130_fd_sc_hd__buf_1 _38835_ (.A(_03346_),
    .X(_08308_));
 sky130_fd_sc_hd__buf_1 _38836_ (.A(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__buf_1 _38837_ (.A(_08047_),
    .X(_08310_));
 sky130_fd_sc_hd__buf_1 _38838_ (.A(_06080_),
    .X(_08311_));
 sky130_fd_sc_hd__nand4_4 _38839_ (.A(_08307_),
    .B(_08309_),
    .C(_08310_),
    .D(_08311_),
    .Y(_08312_));
 sky130_fd_sc_hd__buf_1 _38840_ (.A(\pcpi_mul.rs1[21] ),
    .X(_08313_));
 sky130_fd_sc_hd__buf_1 _38841_ (.A(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__buf_1 _38842_ (.A(_08314_),
    .X(_08315_));
 sky130_fd_sc_hd__nand2_4 _38843_ (.A(_08315_),
    .B(_05955_),
    .Y(_08316_));
 sky130_vsdinv _38844_ (.A(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__a21oi_4 _38845_ (.A1(_08306_),
    .A2(_08312_),
    .B1(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__nand3_4 _38846_ (.A(_08306_),
    .B(_08312_),
    .C(_08317_),
    .Y(_08319_));
 sky130_vsdinv _38847_ (.A(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__nor2_4 _38848_ (.A(_08318_),
    .B(_08320_),
    .Y(_08321_));
 sky130_vsdinv _38849_ (.A(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__o21ai_4 _38850_ (.A1(_08301_),
    .A2(_08304_),
    .B1(_08322_),
    .Y(_08323_));
 sky130_vsdinv _38851_ (.A(_08301_),
    .Y(_08324_));
 sky130_fd_sc_hd__nand3_4 _38852_ (.A(_08324_),
    .B(_08321_),
    .C(_08303_),
    .Y(_08325_));
 sky130_fd_sc_hd__nand2_4 _38853_ (.A(_08323_),
    .B(_08325_),
    .Y(_08326_));
 sky130_vsdinv _38854_ (.A(_08040_),
    .Y(_08327_));
 sky130_fd_sc_hd__o21ai_4 _38855_ (.A1(_08038_),
    .A2(_08063_),
    .B1(_08327_),
    .Y(_08328_));
 sky130_vsdinv _38856_ (.A(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__nand2_4 _38857_ (.A(_08326_),
    .B(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__nand3_4 _38858_ (.A(_08323_),
    .B(_08328_),
    .C(_08325_),
    .Y(_08331_));
 sky130_fd_sc_hd__nand2_4 _38859_ (.A(_08330_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__a21boi_4 _38860_ (.A1(_08049_),
    .A2(_08058_),
    .B1_N(_08053_),
    .Y(_08333_));
 sky130_fd_sc_hd__nand2_4 _38861_ (.A(_08332_),
    .B(_08333_),
    .Y(_08334_));
 sky130_vsdinv _38862_ (.A(_08333_),
    .Y(_08335_));
 sky130_fd_sc_hd__nand3_4 _38863_ (.A(_08330_),
    .B(_08335_),
    .C(_08331_),
    .Y(_08336_));
 sky130_fd_sc_hd__and2_4 _38864_ (.A(_08334_),
    .B(_08336_),
    .X(_08337_));
 sky130_vsdinv _38865_ (.A(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__nand2_4 _38866_ (.A(_08288_),
    .B(_08338_),
    .Y(_08339_));
 sky130_fd_sc_hd__nand3_4 _38867_ (.A(_08337_),
    .B(_08285_),
    .C(_08287_),
    .Y(_08340_));
 sky130_fd_sc_hd__nand2_4 _38868_ (.A(_08339_),
    .B(_08340_),
    .Y(_08341_));
 sky130_fd_sc_hd__nand2_4 _38869_ (.A(_08341_),
    .B(_08187_),
    .Y(_08342_));
 sky130_vsdinv _38870_ (.A(_08187_),
    .Y(_08343_));
 sky130_fd_sc_hd__nand3_4 _38871_ (.A(_08339_),
    .B(_08343_),
    .C(_08340_),
    .Y(_08344_));
 sky130_fd_sc_hd__nand2_4 _38872_ (.A(_08342_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__nand2_4 _38873_ (.A(_08113_),
    .B(_08107_),
    .Y(_08346_));
 sky130_vsdinv _38874_ (.A(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__nand2_4 _38875_ (.A(_08345_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nand3_4 _38876_ (.A(_08342_),
    .B(_08346_),
    .C(_08344_),
    .Y(_08349_));
 sky130_fd_sc_hd__nand2_4 _38877_ (.A(_08348_),
    .B(_08349_),
    .Y(_08350_));
 sky130_vsdinv _38878_ (.A(_08139_),
    .Y(_08351_));
 sky130_fd_sc_hd__a21oi_4 _38879_ (.A1(_08138_),
    .A2(_08143_),
    .B1(_08351_),
    .Y(_08352_));
 sky130_vsdinv _38880_ (.A(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand2_4 _38881_ (.A(_07740_),
    .B(_03541_),
    .Y(_08354_));
 sky130_fd_sc_hd__nand2_4 _38882_ (.A(_07526_),
    .B(_08128_),
    .Y(_08355_));
 sky130_fd_sc_hd__nand2_4 _38883_ (.A(_08354_),
    .B(_08355_),
    .Y(_08356_));
 sky130_fd_sc_hd__buf_1 _38884_ (.A(_03535_),
    .X(_08357_));
 sky130_fd_sc_hd__buf_1 _38885_ (.A(_07716_),
    .X(_08358_));
 sky130_fd_sc_hd__nand4_4 _38886_ (.A(_06072_),
    .B(_07208_),
    .C(_08357_),
    .D(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__nand2_4 _38887_ (.A(_06938_),
    .B(_08132_),
    .Y(_08360_));
 sky130_vsdinv _38888_ (.A(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__a21o_4 _38889_ (.A1(_08356_),
    .A2(_08359_),
    .B1(_08361_),
    .X(_08362_));
 sky130_fd_sc_hd__nand3_4 _38890_ (.A(_08356_),
    .B(_08359_),
    .C(_08361_),
    .Y(_08363_));
 sky130_fd_sc_hd__nand2_4 _38891_ (.A(_08362_),
    .B(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__maj3_4 _38892_ (.A(_08189_),
    .B(_08192_),
    .C(_08195_),
    .X(_08365_));
 sky130_fd_sc_hd__nand2_4 _38893_ (.A(_08364_),
    .B(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__o21ai_4 _38894_ (.A1(_08189_),
    .A2(_08200_),
    .B1(_08199_),
    .Y(_08367_));
 sky130_fd_sc_hd__nand3_4 _38895_ (.A(_08367_),
    .B(_08363_),
    .C(_08362_),
    .Y(_08368_));
 sky130_fd_sc_hd__a21boi_4 _38896_ (.A1(_08130_),
    .A2(_08134_),
    .B1_N(_08131_),
    .Y(_08369_));
 sky130_vsdinv _38897_ (.A(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__nand3_4 _38898_ (.A(_08366_),
    .B(_08368_),
    .C(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__nand2_4 _38899_ (.A(_08366_),
    .B(_08368_),
    .Y(_08372_));
 sky130_fd_sc_hd__nand2_4 _38900_ (.A(_08372_),
    .B(_08369_),
    .Y(_08373_));
 sky130_fd_sc_hd__nand3_4 _38901_ (.A(_08353_),
    .B(_08371_),
    .C(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__nand2_4 _38902_ (.A(_08373_),
    .B(_08371_),
    .Y(_08375_));
 sky130_fd_sc_hd__nand2_4 _38903_ (.A(_08375_),
    .B(_08352_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand2_4 _38904_ (.A(_08374_),
    .B(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__nand2_4 _38905_ (.A(_03275_),
    .B(_07193_),
    .Y(_08378_));
 sky130_fd_sc_hd__nand2_4 _38906_ (.A(_06549_),
    .B(_07050_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand2_4 _38907_ (.A(_08378_),
    .B(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__buf_1 _38908_ (.A(_06154_),
    .X(_08381_));
 sky130_fd_sc_hd__nand4_4 _38909_ (.A(_08381_),
    .B(_06346_),
    .C(_03517_),
    .D(_07362_),
    .Y(_08382_));
 sky130_fd_sc_hd__buf_1 _38910_ (.A(_03511_),
    .X(_08383_));
 sky130_fd_sc_hd__nand2_4 _38911_ (.A(_06349_),
    .B(_08383_),
    .Y(_08384_));
 sky130_vsdinv _38912_ (.A(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__a21o_4 _38913_ (.A1(_08380_),
    .A2(_08382_),
    .B1(_08385_),
    .X(_08386_));
 sky130_fd_sc_hd__nand3_4 _38914_ (.A(_08380_),
    .B(_08382_),
    .C(_08385_),
    .Y(_08387_));
 sky130_fd_sc_hd__a21boi_4 _38915_ (.A1(_08150_),
    .A2(_08153_),
    .B1_N(_08151_),
    .Y(_08388_));
 sky130_fd_sc_hd__a21boi_4 _38916_ (.A1(_08386_),
    .A2(_08387_),
    .B1_N(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__nand2_4 _38917_ (.A(_08386_),
    .B(_08387_),
    .Y(_08390_));
 sky130_fd_sc_hd__nor2_4 _38918_ (.A(_08388_),
    .B(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__buf_1 _38919_ (.A(_06848_),
    .X(_08392_));
 sky130_fd_sc_hd__nand2_4 _38920_ (.A(_08392_),
    .B(_07754_),
    .Y(_08393_));
 sky130_fd_sc_hd__buf_1 _38921_ (.A(_07653_),
    .X(_08394_));
 sky130_fd_sc_hd__nand2_4 _38922_ (.A(_08394_),
    .B(_07756_),
    .Y(_08395_));
 sky130_fd_sc_hd__nand2_4 _38923_ (.A(_06847_),
    .B(_06887_),
    .Y(_08396_));
 sky130_fd_sc_hd__nand2_4 _38924_ (.A(_08395_),
    .B(_08396_),
    .Y(_08397_));
 sky130_fd_sc_hd__nand4_4 _38925_ (.A(_06977_),
    .B(_07280_),
    .C(_06743_),
    .D(_07344_),
    .Y(_08398_));
 sky130_fd_sc_hd__nand2_4 _38926_ (.A(_08397_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__xor2_4 _38927_ (.A(_08393_),
    .B(_08399_),
    .X(_08400_));
 sky130_vsdinv _38928_ (.A(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__o21a_4 _38929_ (.A1(_08389_),
    .A2(_08391_),
    .B1(_08401_),
    .X(_08402_));
 sky130_vsdinv _38930_ (.A(_08391_),
    .Y(_08403_));
 sky130_vsdinv _38931_ (.A(_08389_),
    .Y(_08404_));
 sky130_fd_sc_hd__nand3_4 _38932_ (.A(_08403_),
    .B(_08404_),
    .C(_08400_),
    .Y(_08405_));
 sky130_vsdinv _38933_ (.A(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__nor2_4 _38934_ (.A(_08402_),
    .B(_08406_),
    .Y(_08407_));
 sky130_vsdinv _38935_ (.A(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__nand2_4 _38936_ (.A(_08377_),
    .B(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__nand3_4 _38937_ (.A(_08407_),
    .B(_08374_),
    .C(_08376_),
    .Y(_08410_));
 sky130_fd_sc_hd__nand2_4 _38938_ (.A(_08409_),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__o21ai_4 _38939_ (.A1(_08178_),
    .A2(_08145_),
    .B1(_08146_),
    .Y(_08412_));
 sky130_vsdinv _38940_ (.A(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__nand2_4 _38941_ (.A(_08411_),
    .B(_08413_),
    .Y(_08414_));
 sky130_fd_sc_hd__nand3_4 _38942_ (.A(_08409_),
    .B(_08412_),
    .C(_08410_),
    .Y(_08415_));
 sky130_fd_sc_hd__nand2_4 _38943_ (.A(_08414_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__nand2_4 _38944_ (.A(_05589_),
    .B(_03566_),
    .Y(_08417_));
 sky130_fd_sc_hd__nand2_4 _38945_ (.A(_06370_),
    .B(_03557_),
    .Y(_08418_));
 sky130_fd_sc_hd__nand2_4 _38946_ (.A(_03253_),
    .B(_03552_),
    .Y(_08419_));
 sky130_fd_sc_hd__nand2_4 _38947_ (.A(_08418_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__nand4_4 _38948_ (.A(_06050_),
    .B(_03253_),
    .C(_07976_),
    .D(_03557_),
    .Y(_08421_));
 sky130_fd_sc_hd__nand2_4 _38949_ (.A(_07360_),
    .B(_03544_),
    .Y(_08422_));
 sky130_vsdinv _38950_ (.A(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__a21o_4 _38951_ (.A1(_08420_),
    .A2(_08421_),
    .B1(_08423_),
    .X(_08424_));
 sky130_fd_sc_hd__nand3_4 _38952_ (.A(_08420_),
    .B(_08421_),
    .C(_08423_),
    .Y(_08425_));
 sky130_fd_sc_hd__nand2_4 _38953_ (.A(_08424_),
    .B(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__xor2_4 _38954_ (.A(_08417_),
    .B(_08426_),
    .X(_08427_));
 sky130_vsdinv _38955_ (.A(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__nand2_4 _38956_ (.A(_08416_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__nand3_4 _38957_ (.A(_08414_),
    .B(_08427_),
    .C(_08415_),
    .Y(_08430_));
 sky130_fd_sc_hd__nand2_4 _38958_ (.A(_08429_),
    .B(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__nand2_4 _38959_ (.A(_08431_),
    .B(_08204_),
    .Y(_08432_));
 sky130_vsdinv _38960_ (.A(_08204_),
    .Y(_08433_));
 sky130_fd_sc_hd__nand3_4 _38961_ (.A(_08433_),
    .B(_08429_),
    .C(_08430_),
    .Y(_08434_));
 sky130_fd_sc_hd__and2_4 _38962_ (.A(_08432_),
    .B(_08434_),
    .X(_08435_));
 sky130_vsdinv _38963_ (.A(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__nand2_4 _38964_ (.A(_08350_),
    .B(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand3_4 _38965_ (.A(_08348_),
    .B(_08435_),
    .C(_08349_),
    .Y(_08438_));
 sky130_fd_sc_hd__nand2_4 _38966_ (.A(_08437_),
    .B(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__nand2_4 _38967_ (.A(_08249_),
    .B(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__nand3_4 _38968_ (.A(_08248_),
    .B(_08438_),
    .C(_08437_),
    .Y(_08441_));
 sky130_fd_sc_hd__nand2_4 _38969_ (.A(_08440_),
    .B(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a21boi_4 _38970_ (.A1(_08067_),
    .A2(_08069_),
    .B1_N(_08070_),
    .Y(_08443_));
 sky130_fd_sc_hd__a21oi_4 _38971_ (.A1(_08122_),
    .A2(_08117_),
    .B1(_08443_),
    .Y(_08444_));
 sky130_vsdinv _38972_ (.A(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__nand3_4 _38973_ (.A(_08122_),
    .B(_08117_),
    .C(_08443_),
    .Y(_08446_));
 sky130_fd_sc_hd__nand2_4 _38974_ (.A(_08445_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__nand2_4 _38975_ (.A(_08442_),
    .B(_08447_),
    .Y(_08448_));
 sky130_vsdinv _38976_ (.A(_08447_),
    .Y(_08449_));
 sky130_fd_sc_hd__nand3_4 _38977_ (.A(_08440_),
    .B(_08449_),
    .C(_08441_),
    .Y(_08450_));
 sky130_fd_sc_hd__nand2_4 _38978_ (.A(_08448_),
    .B(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__o21ai_4 _38979_ (.A1(_08218_),
    .A2(_08213_),
    .B1(_08214_),
    .Y(_08452_));
 sky130_vsdinv _38980_ (.A(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_4 _38981_ (.A(_08451_),
    .B(_08453_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand3_4 _38982_ (.A(_08448_),
    .B(_08452_),
    .C(_08450_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand2_4 _38983_ (.A(_08454_),
    .B(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__a21oi_4 _38984_ (.A1(_07912_),
    .A2(_07907_),
    .B1(_08216_),
    .Y(_08457_));
 sky130_vsdinv _38985_ (.A(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__nand2_4 _38986_ (.A(_08456_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__nand3_4 _38987_ (.A(_08454_),
    .B(_08457_),
    .C(_08455_),
    .Y(_08460_));
 sky130_fd_sc_hd__nand2_4 _38988_ (.A(_08459_),
    .B(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__a21boi_4 _38989_ (.A1(_08227_),
    .A2(_08231_),
    .B1_N(_08229_),
    .Y(_08462_));
 sky130_fd_sc_hd__nand2_4 _38990_ (.A(_08461_),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nand2_4 _38991_ (.A(_08234_),
    .B(_08229_),
    .Y(_08464_));
 sky130_fd_sc_hd__nand3_4 _38992_ (.A(_08464_),
    .B(_08460_),
    .C(_08459_),
    .Y(_08465_));
 sky130_fd_sc_hd__and2_4 _38993_ (.A(_08463_),
    .B(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__o21ai_4 _38994_ (.A1(_08241_),
    .A2(_08247_),
    .B1(_08239_),
    .Y(_08467_));
 sky130_fd_sc_hd__xor2_4 _38995_ (.A(_08466_),
    .B(_08467_),
    .X(_01426_));
 sky130_fd_sc_hd__nand2_4 _38996_ (.A(_08438_),
    .B(_08434_),
    .Y(_08468_));
 sky130_vsdinv _38997_ (.A(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__buf_1 _38998_ (.A(_06991_),
    .X(_08470_));
 sky130_fd_sc_hd__nand2_4 _38999_ (.A(_08470_),
    .B(_06482_),
    .Y(_08471_));
 sky130_fd_sc_hd__nand2_4 _39000_ (.A(_03318_),
    .B(_07467_),
    .Y(_08472_));
 sky130_fd_sc_hd__nand2_4 _39001_ (.A(_08471_),
    .B(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__nand4_4 _39002_ (.A(_07299_),
    .B(_07439_),
    .C(_06791_),
    .D(_07470_),
    .Y(_08474_));
 sky130_fd_sc_hd__nand2_4 _39003_ (.A(_07294_),
    .B(_06949_),
    .Y(_08475_));
 sky130_vsdinv _39004_ (.A(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__a21o_4 _39005_ (.A1(_08473_),
    .A2(_08474_),
    .B1(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__nand3_4 _39006_ (.A(_08473_),
    .B(_08474_),
    .C(_08476_),
    .Y(_08478_));
 sky130_fd_sc_hd__nand2_4 _39007_ (.A(_08477_),
    .B(_08478_),
    .Y(_08479_));
 sky130_vsdinv _39008_ (.A(_08393_),
    .Y(_08480_));
 sky130_fd_sc_hd__a21boi_4 _39009_ (.A1(_08397_),
    .A2(_08480_),
    .B1_N(_08398_),
    .Y(_08481_));
 sky130_fd_sc_hd__nand2_4 _39010_ (.A(_08479_),
    .B(_08481_),
    .Y(_08482_));
 sky130_vsdinv _39011_ (.A(_08481_),
    .Y(_08483_));
 sky130_fd_sc_hd__nand3_4 _39012_ (.A(_08483_),
    .B(_08478_),
    .C(_08477_),
    .Y(_08484_));
 sky130_fd_sc_hd__a21boi_4 _39013_ (.A1(_08261_),
    .A2(_08266_),
    .B1_N(_08262_),
    .Y(_08485_));
 sky130_vsdinv _39014_ (.A(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__a21o_4 _39015_ (.A1(_08482_),
    .A2(_08484_),
    .B1(_08486_),
    .X(_08487_));
 sky130_fd_sc_hd__nand3_4 _39016_ (.A(_08482_),
    .B(_08484_),
    .C(_08486_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand2_4 _39017_ (.A(_08487_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__a21oi_4 _39018_ (.A1(_08404_),
    .A2(_08400_),
    .B1(_08391_),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_4 _39019_ (.A(_08489_),
    .B(_08490_),
    .Y(_08491_));
 sky130_fd_sc_hd__o21ai_4 _39020_ (.A1(_08389_),
    .A2(_08401_),
    .B1(_08403_),
    .Y(_08492_));
 sky130_fd_sc_hd__nand3_4 _39021_ (.A(_08492_),
    .B(_08488_),
    .C(_08487_),
    .Y(_08493_));
 sky130_fd_sc_hd__nand2_4 _39022_ (.A(_08491_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__a21boi_4 _39023_ (.A1(_08269_),
    .A2(_08271_),
    .B1_N(_08272_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand2_4 _39024_ (.A(_08494_),
    .B(_08495_),
    .Y(_08496_));
 sky130_vsdinv _39025_ (.A(_08495_),
    .Y(_08497_));
 sky130_fd_sc_hd__nand3_4 _39026_ (.A(_08491_),
    .B(_08493_),
    .C(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__nand2_4 _39027_ (.A(_08496_),
    .B(_08498_),
    .Y(_08499_));
 sky130_fd_sc_hd__nand2_4 _39028_ (.A(_08282_),
    .B(_08276_),
    .Y(_08500_));
 sky130_vsdinv _39029_ (.A(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__nand2_4 _39030_ (.A(_08499_),
    .B(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__nand3_4 _39031_ (.A(_08500_),
    .B(_08496_),
    .C(_08498_),
    .Y(_08503_));
 sky130_fd_sc_hd__nand2_4 _39032_ (.A(_08502_),
    .B(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__buf_1 _39033_ (.A(_03470_),
    .X(_08505_));
 sky130_fd_sc_hd__nand2_4 _39034_ (.A(_03332_),
    .B(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__buf_1 _39035_ (.A(_06134_),
    .X(_08507_));
 sky130_fd_sc_hd__nand2_4 _39036_ (.A(_07629_),
    .B(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__nand2_4 _39037_ (.A(_08506_),
    .B(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__buf_1 _39038_ (.A(_03335_),
    .X(_08510_));
 sky130_fd_sc_hd__nand4_4 _39039_ (.A(_07626_),
    .B(_08510_),
    .C(_08028_),
    .D(_06322_),
    .Y(_08511_));
 sky130_fd_sc_hd__nand2_4 _39040_ (.A(_08046_),
    .B(_03453_),
    .Y(_08512_));
 sky130_vsdinv _39041_ (.A(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__a21o_4 _39042_ (.A1(_08509_),
    .A2(_08511_),
    .B1(_08513_),
    .X(_08514_));
 sky130_fd_sc_hd__nand3_4 _39043_ (.A(_08509_),
    .B(_08511_),
    .C(_08513_),
    .Y(_08515_));
 sky130_fd_sc_hd__a21boi_4 _39044_ (.A1(_08293_),
    .A2(_08297_),
    .B1_N(_08295_),
    .Y(_08516_));
 sky130_fd_sc_hd__a21boi_4 _39045_ (.A1(_08514_),
    .A2(_08515_),
    .B1_N(_08516_),
    .Y(_08517_));
 sky130_vsdinv _39046_ (.A(_08516_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand3_4 _39047_ (.A(_08518_),
    .B(_08515_),
    .C(_08514_),
    .Y(_08519_));
 sky130_vsdinv _39048_ (.A(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__nor2_4 _39049_ (.A(_08517_),
    .B(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__buf_1 _39050_ (.A(_08054_),
    .X(_08522_));
 sky130_fd_sc_hd__buf_1 _39051_ (.A(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__nand2_4 _39052_ (.A(_08523_),
    .B(_05910_),
    .Y(_08524_));
 sky130_fd_sc_hd__o21ai_4 _39053_ (.A1(_03355_),
    .A2(_07619_),
    .B1(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__buf_1 _39054_ (.A(_08056_),
    .X(_08526_));
 sky130_fd_sc_hd__buf_1 _39055_ (.A(_08313_),
    .X(_08527_));
 sky130_fd_sc_hd__buf_1 _39056_ (.A(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__nand4_4 _39057_ (.A(_08526_),
    .B(_08528_),
    .C(_07002_),
    .D(_07154_),
    .Y(_08529_));
 sky130_fd_sc_hd__buf_1 _39058_ (.A(\pcpi_mul.rs1[22] ),
    .X(_08530_));
 sky130_fd_sc_hd__buf_1 _39059_ (.A(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__nand2_4 _39060_ (.A(_08531_),
    .B(_06086_),
    .Y(_08532_));
 sky130_vsdinv _39061_ (.A(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__a21oi_4 _39062_ (.A1(_08525_),
    .A2(_08529_),
    .B1(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__nand3_4 _39063_ (.A(_08525_),
    .B(_08529_),
    .C(_08533_),
    .Y(_08535_));
 sky130_vsdinv _39064_ (.A(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__nor2_4 _39065_ (.A(_08534_),
    .B(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__nand2_4 _39066_ (.A(_08521_),
    .B(_08537_),
    .Y(_08538_));
 sky130_vsdinv _39067_ (.A(_08537_),
    .Y(_08539_));
 sky130_fd_sc_hd__o21ai_4 _39068_ (.A1(_08517_),
    .A2(_08520_),
    .B1(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__nand2_4 _39069_ (.A(_08538_),
    .B(_08540_),
    .Y(_08541_));
 sky130_fd_sc_hd__a21oi_4 _39070_ (.A1(_08324_),
    .A2(_08321_),
    .B1(_08304_),
    .Y(_08542_));
 sky130_fd_sc_hd__nand2_4 _39071_ (.A(_08541_),
    .B(_08542_),
    .Y(_08543_));
 sky130_vsdinv _39072_ (.A(_08542_),
    .Y(_08544_));
 sky130_fd_sc_hd__nand3_4 _39073_ (.A(_08544_),
    .B(_08538_),
    .C(_08540_),
    .Y(_08545_));
 sky130_fd_sc_hd__nand2_4 _39074_ (.A(_08543_),
    .B(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__a21boi_4 _39075_ (.A1(_08306_),
    .A2(_08317_),
    .B1_N(_08312_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand2_4 _39076_ (.A(_08546_),
    .B(_08547_),
    .Y(_08548_));
 sky130_vsdinv _39077_ (.A(_08547_),
    .Y(_08549_));
 sky130_fd_sc_hd__nand3_4 _39078_ (.A(_08543_),
    .B(_08545_),
    .C(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__nand2_4 _39079_ (.A(_08548_),
    .B(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__nand2_4 _39080_ (.A(_08504_),
    .B(_08551_),
    .Y(_08552_));
 sky130_vsdinv _39081_ (.A(_08551_),
    .Y(_08553_));
 sky130_fd_sc_hd__nand3_4 _39082_ (.A(_08553_),
    .B(_08502_),
    .C(_08503_),
    .Y(_08554_));
 sky130_fd_sc_hd__nand2_4 _39083_ (.A(_08552_),
    .B(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__nand2_4 _39084_ (.A(_08555_),
    .B(_08415_),
    .Y(_08556_));
 sky130_vsdinv _39085_ (.A(_08415_),
    .Y(_08557_));
 sky130_fd_sc_hd__nand3_4 _39086_ (.A(_08552_),
    .B(_08557_),
    .C(_08554_),
    .Y(_08558_));
 sky130_fd_sc_hd__nand2_4 _39087_ (.A(_08556_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__a21boi_4 _39088_ (.A1(_08337_),
    .A2(_08287_),
    .B1_N(_08285_),
    .Y(_08560_));
 sky130_fd_sc_hd__nand2_4 _39089_ (.A(_08559_),
    .B(_08560_),
    .Y(_08561_));
 sky130_vsdinv _39090_ (.A(_08560_),
    .Y(_08562_));
 sky130_fd_sc_hd__nand3_4 _39091_ (.A(_08556_),
    .B(_08562_),
    .C(_08558_),
    .Y(_08563_));
 sky130_fd_sc_hd__nand2_4 _39092_ (.A(_08561_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__buf_1 _39093_ (.A(_03268_),
    .X(_08565_));
 sky130_fd_sc_hd__buf_1 _39094_ (.A(_07921_),
    .X(_08566_));
 sky130_fd_sc_hd__nand2_4 _39095_ (.A(_08565_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__buf_1 _39096_ (.A(_07712_),
    .X(_08568_));
 sky130_fd_sc_hd__nand2_4 _39097_ (.A(_06244_),
    .B(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__nand2_4 _39098_ (.A(_08567_),
    .B(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__buf_1 _39099_ (.A(\pcpi_mul.rs2[16] ),
    .X(_08571_));
 sky130_fd_sc_hd__buf_1 _39100_ (.A(_08571_),
    .X(_08572_));
 sky130_fd_sc_hd__nand4_4 _39101_ (.A(_07938_),
    .B(_07939_),
    .C(_08572_),
    .D(_07710_),
    .Y(_08573_));
 sky130_fd_sc_hd__nand2_4 _39102_ (.A(_08381_),
    .B(_07562_),
    .Y(_08574_));
 sky130_vsdinv _39103_ (.A(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__a21o_4 _39104_ (.A1(_08570_),
    .A2(_08573_),
    .B1(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__nand3_4 _39105_ (.A(_08570_),
    .B(_08573_),
    .C(_08575_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand2_4 _39106_ (.A(_08576_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__a21boi_4 _39107_ (.A1(_08420_),
    .A2(_08423_),
    .B1_N(_08421_),
    .Y(_08579_));
 sky130_fd_sc_hd__nand2_4 _39108_ (.A(_08578_),
    .B(_08579_),
    .Y(_08580_));
 sky130_vsdinv _39109_ (.A(_08579_),
    .Y(_08581_));
 sky130_fd_sc_hd__nand3_4 _39110_ (.A(_08581_),
    .B(_08577_),
    .C(_08576_),
    .Y(_08582_));
 sky130_fd_sc_hd__nand2_4 _39111_ (.A(_08580_),
    .B(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__a21boi_4 _39112_ (.A1(_08356_),
    .A2(_08361_),
    .B1_N(_08359_),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_4 _39113_ (.A(_08583_),
    .B(_08584_),
    .Y(_08585_));
 sky130_vsdinv _39114_ (.A(_08584_),
    .Y(_08586_));
 sky130_fd_sc_hd__nand3_4 _39115_ (.A(_08580_),
    .B(_08582_),
    .C(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__nand2_4 _39116_ (.A(_08585_),
    .B(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__a21boi_4 _39117_ (.A1(_08366_),
    .A2(_08370_),
    .B1_N(_08368_),
    .Y(_08589_));
 sky130_fd_sc_hd__nand2_4 _39118_ (.A(_08588_),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__nand2_4 _39119_ (.A(_08371_),
    .B(_08368_),
    .Y(_08591_));
 sky130_fd_sc_hd__nand3_4 _39120_ (.A(_08591_),
    .B(_08587_),
    .C(_08585_),
    .Y(_08592_));
 sky130_fd_sc_hd__nand4_4 _39121_ (.A(_03280_),
    .B(_06349_),
    .C(_07521_),
    .D(_03525_),
    .Y(_08593_));
 sky130_fd_sc_hd__nand2_4 _39122_ (.A(_06549_),
    .B(_07193_),
    .Y(_08594_));
 sky130_fd_sc_hd__nand2_4 _39123_ (.A(_08167_),
    .B(_07050_),
    .Y(_08595_));
 sky130_fd_sc_hd__nand2_4 _39124_ (.A(_08594_),
    .B(_08595_),
    .Y(_08596_));
 sky130_fd_sc_hd__a2bb2o_4 _39125_ (.A1_N(_03295_),
    .A2_N(_06882_),
    .B1(_08593_),
    .B2(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__buf_1 _39126_ (.A(_08383_),
    .X(_08598_));
 sky130_fd_sc_hd__nand4_4 _39127_ (.A(_06981_),
    .B(_08596_),
    .C(_08593_),
    .D(_08598_),
    .Y(_08599_));
 sky130_fd_sc_hd__nand2_4 _39128_ (.A(_08597_),
    .B(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__a21boi_4 _39129_ (.A1(_08380_),
    .A2(_08385_),
    .B1_N(_08382_),
    .Y(_08601_));
 sky130_fd_sc_hd__nand2_4 _39130_ (.A(_08600_),
    .B(_08601_),
    .Y(_08602_));
 sky130_vsdinv _39131_ (.A(_08601_),
    .Y(_08603_));
 sky130_fd_sc_hd__nand3_4 _39132_ (.A(_08603_),
    .B(_08597_),
    .C(_08599_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand2_4 _39133_ (.A(_07146_),
    .B(_03495_),
    .Y(_08605_));
 sky130_fd_sc_hd__buf_1 _39134_ (.A(\pcpi_mul.rs1[11] ),
    .X(_08606_));
 sky130_fd_sc_hd__buf_1 _39135_ (.A(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__nand2_4 _39136_ (.A(_08607_),
    .B(_07543_),
    .Y(_08608_));
 sky130_fd_sc_hd__nand2_4 _39137_ (.A(_08392_),
    .B(_07212_),
    .Y(_08609_));
 sky130_fd_sc_hd__nand2_4 _39138_ (.A(_08608_),
    .B(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__nand4_4 _39139_ (.A(_06571_),
    .B(_06995_),
    .C(_07956_),
    .D(_06893_),
    .Y(_08611_));
 sky130_fd_sc_hd__nand2_4 _39140_ (.A(_08610_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__xor2_4 _39141_ (.A(_08605_),
    .B(_08612_),
    .X(_08613_));
 sky130_fd_sc_hd__a21oi_4 _39142_ (.A1(_08602_),
    .A2(_08604_),
    .B1(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__nand3_4 _39143_ (.A(_08602_),
    .B(_08613_),
    .C(_08604_),
    .Y(_08615_));
 sky130_vsdinv _39144_ (.A(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__nor2_4 _39145_ (.A(_08614_),
    .B(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__a21oi_4 _39146_ (.A1(_08590_),
    .A2(_08592_),
    .B1(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__nand3_4 _39147_ (.A(_08590_),
    .B(_08592_),
    .C(_08617_),
    .Y(_08619_));
 sky130_vsdinv _39148_ (.A(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__a21boi_4 _39149_ (.A1(_08407_),
    .A2(_08376_),
    .B1_N(_08374_),
    .Y(_08621_));
 sky130_fd_sc_hd__o21ai_4 _39150_ (.A1(_08618_),
    .A2(_08620_),
    .B1(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__nand2_4 _39151_ (.A(_08410_),
    .B(_08374_),
    .Y(_08623_));
 sky130_vsdinv _39152_ (.A(_08618_),
    .Y(_08624_));
 sky130_fd_sc_hd__nand3_4 _39153_ (.A(_08623_),
    .B(_08624_),
    .C(_08619_),
    .Y(_08625_));
 sky130_fd_sc_hd__nand2_4 _39154_ (.A(_08622_),
    .B(_08625_),
    .Y(_08626_));
 sky130_fd_sc_hd__nand4_4 _39155_ (.A(_05588_),
    .B(_08424_),
    .C(_03566_),
    .D(_08425_),
    .Y(_08627_));
 sky130_vsdinv _39156_ (.A(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__buf_1 _39157_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08629_));
 sky130_fd_sc_hd__buf_1 _39158_ (.A(_08629_),
    .X(_08630_));
 sky130_fd_sc_hd__buf_1 _39159_ (.A(_08630_),
    .X(_08631_));
 sky130_fd_sc_hd__buf_1 _39160_ (.A(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__nand2_4 _39161_ (.A(_05895_),
    .B(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__buf_1 _39162_ (.A(\pcpi_mul.rs2[21] ),
    .X(_08634_));
 sky130_fd_sc_hd__buf_1 _39163_ (.A(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__buf_1 _39164_ (.A(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__nand2_4 _39165_ (.A(_06276_),
    .B(_08636_),
    .Y(_08637_));
 sky130_fd_sc_hd__xnor2_4 _39166_ (.A(_08633_),
    .B(_08637_),
    .Y(_08638_));
 sky130_vsdinv _39167_ (.A(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__buf_1 _39168_ (.A(\pcpi_mul.rs2[18] ),
    .X(_08640_));
 sky130_fd_sc_hd__nand2_4 _39169_ (.A(_06141_),
    .B(_08640_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand2_4 _39170_ (.A(_06380_),
    .B(_08197_),
    .Y(_08642_));
 sky130_fd_sc_hd__buf_1 _39171_ (.A(\pcpi_mul.rs2[19] ),
    .X(_08643_));
 sky130_fd_sc_hd__nand2_4 _39172_ (.A(_05942_),
    .B(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__nand2_4 _39173_ (.A(_08642_),
    .B(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__buf_1 _39174_ (.A(_03551_),
    .X(_08646_));
 sky130_fd_sc_hd__buf_1 _39175_ (.A(_03556_),
    .X(_08647_));
 sky130_fd_sc_hd__nand4_4 _39176_ (.A(_06380_),
    .B(_06226_),
    .C(_08646_),
    .D(_08647_),
    .Y(_08648_));
 sky130_fd_sc_hd__nand2_4 _39177_ (.A(_08645_),
    .B(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__xor2_4 _39178_ (.A(_08641_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__xor2_4 _39179_ (.A(_08639_),
    .B(_08650_),
    .X(_08651_));
 sky130_fd_sc_hd__xor2_4 _39180_ (.A(_08628_),
    .B(_08651_),
    .X(_08652_));
 sky130_vsdinv _39181_ (.A(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__nand2_4 _39182_ (.A(_08626_),
    .B(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__nand3_4 _39183_ (.A(_08622_),
    .B(_08625_),
    .C(_08652_),
    .Y(_08655_));
 sky130_fd_sc_hd__nand2_4 _39184_ (.A(_08654_),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__nand2_4 _39185_ (.A(_08656_),
    .B(_08430_),
    .Y(_08657_));
 sky130_vsdinv _39186_ (.A(_08430_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand3_4 _39187_ (.A(_08654_),
    .B(_08658_),
    .C(_08655_),
    .Y(_08659_));
 sky130_fd_sc_hd__and2_4 _39188_ (.A(_08657_),
    .B(_08659_),
    .X(_08660_));
 sky130_vsdinv _39189_ (.A(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__nand2_4 _39190_ (.A(_08564_),
    .B(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__nand3_4 _39191_ (.A(_08561_),
    .B(_08660_),
    .C(_08563_),
    .Y(_08663_));
 sky130_fd_sc_hd__nand2_4 _39192_ (.A(_08662_),
    .B(_08663_),
    .Y(_08664_));
 sky130_fd_sc_hd__nand2_4 _39193_ (.A(_08469_),
    .B(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__nand3_4 _39194_ (.A(_08468_),
    .B(_08662_),
    .C(_08663_),
    .Y(_08666_));
 sky130_fd_sc_hd__nand2_4 _39195_ (.A(_08665_),
    .B(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__a21boi_4 _39196_ (.A1(_08330_),
    .A2(_08335_),
    .B1_N(_08331_),
    .Y(_08668_));
 sky130_fd_sc_hd__nand2_4 _39197_ (.A(_08349_),
    .B(_08344_),
    .Y(_08669_));
 sky130_fd_sc_hd__xor2_4 _39198_ (.A(_08668_),
    .B(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__nand2_4 _39199_ (.A(_08667_),
    .B(_08670_),
    .Y(_08671_));
 sky130_vsdinv _39200_ (.A(_08670_),
    .Y(_08672_));
 sky130_fd_sc_hd__nand3_4 _39201_ (.A(_08672_),
    .B(_08665_),
    .C(_08666_),
    .Y(_08673_));
 sky130_fd_sc_hd__nand2_4 _39202_ (.A(_08671_),
    .B(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__a21boi_4 _39203_ (.A1(_08440_),
    .A2(_08449_),
    .B1_N(_08441_),
    .Y(_08675_));
 sky130_fd_sc_hd__nand2_4 _39204_ (.A(_08674_),
    .B(_08675_),
    .Y(_08676_));
 sky130_vsdinv _39205_ (.A(_08675_),
    .Y(_08677_));
 sky130_fd_sc_hd__nand3_4 _39206_ (.A(_08677_),
    .B(_08671_),
    .C(_08673_),
    .Y(_08678_));
 sky130_fd_sc_hd__nand2_4 _39207_ (.A(_08676_),
    .B(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__nand2_4 _39208_ (.A(_08679_),
    .B(_08445_),
    .Y(_08680_));
 sky130_fd_sc_hd__nand3_4 _39209_ (.A(_08676_),
    .B(_08678_),
    .C(_08444_),
    .Y(_08681_));
 sky130_fd_sc_hd__nand2_4 _39210_ (.A(_08680_),
    .B(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__a21boi_4 _39211_ (.A1(_08454_),
    .A2(_08457_),
    .B1_N(_08455_),
    .Y(_08683_));
 sky130_fd_sc_hd__nand2_4 _39212_ (.A(_08682_),
    .B(_08683_),
    .Y(_08684_));
 sky130_vsdinv _39213_ (.A(_08683_),
    .Y(_08685_));
 sky130_fd_sc_hd__nand3_4 _39214_ (.A(_08685_),
    .B(_08681_),
    .C(_08680_),
    .Y(_08686_));
 sky130_fd_sc_hd__and2_4 _39215_ (.A(_08684_),
    .B(_08686_),
    .X(_08687_));
 sky130_fd_sc_hd__nand4_4 _39216_ (.A(_08239_),
    .B(_08238_),
    .C(_08463_),
    .D(_08465_),
    .Y(_08688_));
 sky130_fd_sc_hd__nand2_4 _39217_ (.A(_08465_),
    .B(_08239_),
    .Y(_08689_));
 sky130_fd_sc_hd__nand2_4 _39218_ (.A(_08689_),
    .B(_08463_),
    .Y(_08690_));
 sky130_fd_sc_hd__o21ai_4 _39219_ (.A1(_08688_),
    .A2(_08247_),
    .B1(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__xor2_4 _39220_ (.A(_08687_),
    .B(_08691_),
    .X(_01427_));
 sky130_fd_sc_hd__a21boi_4 _39221_ (.A1(_08676_),
    .A2(_08444_),
    .B1_N(_08678_),
    .Y(_08692_));
 sky130_vsdinv _39222_ (.A(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__nand2_4 _39223_ (.A(_08663_),
    .B(_08659_),
    .Y(_08694_));
 sky130_vsdinv _39224_ (.A(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__nand2_4 _39225_ (.A(_07432_),
    .B(_06372_),
    .Y(_08696_));
 sky130_fd_sc_hd__nand2_4 _39226_ (.A(_07435_),
    .B(_06376_),
    .Y(_08697_));
 sky130_fd_sc_hd__nand2_4 _39227_ (.A(_08696_),
    .B(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__nand4_4 _39228_ (.A(_07439_),
    .B(_07294_),
    .C(_03481_),
    .D(_06939_),
    .Y(_08699_));
 sky130_fd_sc_hd__nand2_4 _39229_ (.A(_07444_),
    .B(_06606_),
    .Y(_08700_));
 sky130_vsdinv _39230_ (.A(_08700_),
    .Y(_08701_));
 sky130_fd_sc_hd__a21o_4 _39231_ (.A1(_08698_),
    .A2(_08699_),
    .B1(_08701_),
    .X(_08702_));
 sky130_fd_sc_hd__nand3_4 _39232_ (.A(_08698_),
    .B(_08699_),
    .C(_08701_),
    .Y(_08703_));
 sky130_fd_sc_hd__nand2_4 _39233_ (.A(_08702_),
    .B(_08703_),
    .Y(_08704_));
 sky130_vsdinv _39234_ (.A(_08605_),
    .Y(_08705_));
 sky130_fd_sc_hd__a21boi_4 _39235_ (.A1(_08610_),
    .A2(_08705_),
    .B1_N(_08611_),
    .Y(_08706_));
 sky130_fd_sc_hd__nand2_4 _39236_ (.A(_08704_),
    .B(_08706_),
    .Y(_08707_));
 sky130_vsdinv _39237_ (.A(_08706_),
    .Y(_08708_));
 sky130_fd_sc_hd__nand3_4 _39238_ (.A(_08708_),
    .B(_08703_),
    .C(_08702_),
    .Y(_08709_));
 sky130_fd_sc_hd__nand2_4 _39239_ (.A(_08707_),
    .B(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__a21boi_4 _39240_ (.A1(_08473_),
    .A2(_08476_),
    .B1_N(_08474_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_4 _39241_ (.A(_08710_),
    .B(_08711_),
    .Y(_08712_));
 sky130_vsdinv _39242_ (.A(_08711_),
    .Y(_08713_));
 sky130_fd_sc_hd__nand3_4 _39243_ (.A(_08707_),
    .B(_08709_),
    .C(_08713_),
    .Y(_08714_));
 sky130_fd_sc_hd__nand2_4 _39244_ (.A(_08712_),
    .B(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__a21boi_4 _39245_ (.A1(_08602_),
    .A2(_08613_),
    .B1_N(_08604_),
    .Y(_08716_));
 sky130_fd_sc_hd__nand2_4 _39246_ (.A(_08715_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__nand2_4 _39247_ (.A(_08615_),
    .B(_08604_),
    .Y(_08718_));
 sky130_fd_sc_hd__nand3_4 _39248_ (.A(_08718_),
    .B(_08714_),
    .C(_08712_),
    .Y(_08719_));
 sky130_fd_sc_hd__nand2_4 _39249_ (.A(_08717_),
    .B(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__a21boi_4 _39250_ (.A1(_08482_),
    .A2(_08486_),
    .B1_N(_08484_),
    .Y(_08721_));
 sky130_fd_sc_hd__nand2_4 _39251_ (.A(_08720_),
    .B(_08721_),
    .Y(_08722_));
 sky130_vsdinv _39252_ (.A(_08721_),
    .Y(_08723_));
 sky130_fd_sc_hd__nand3_4 _39253_ (.A(_08717_),
    .B(_08719_),
    .C(_08723_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand2_4 _39254_ (.A(_08722_),
    .B(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__a21boi_4 _39255_ (.A1(_08491_),
    .A2(_08497_),
    .B1_N(_08493_),
    .Y(_08726_));
 sky130_fd_sc_hd__nand2_4 _39256_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__nand2_4 _39257_ (.A(_08498_),
    .B(_08493_),
    .Y(_08728_));
 sky130_fd_sc_hd__nand3_4 _39258_ (.A(_08728_),
    .B(_08724_),
    .C(_08722_),
    .Y(_08729_));
 sky130_fd_sc_hd__nand2_4 _39259_ (.A(_08727_),
    .B(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__buf_1 _39260_ (.A(_06051_),
    .X(_08731_));
 sky130_fd_sc_hd__nand2_4 _39261_ (.A(_08510_),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__buf_1 _39262_ (.A(_03340_),
    .X(_08733_));
 sky130_fd_sc_hd__buf_1 _39263_ (.A(_06134_),
    .X(_08734_));
 sky130_fd_sc_hd__nand2_4 _39264_ (.A(_08733_),
    .B(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__nand2_4 _39265_ (.A(_08732_),
    .B(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__nand4_4 _39266_ (.A(_08510_),
    .B(_08733_),
    .C(_08734_),
    .D(_08731_),
    .Y(_08737_));
 sky130_fd_sc_hd__nand2_4 _39267_ (.A(_08308_),
    .B(_06327_),
    .Y(_08738_));
 sky130_vsdinv _39268_ (.A(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__a21o_4 _39269_ (.A1(_08736_),
    .A2(_08737_),
    .B1(_08739_),
    .X(_08740_));
 sky130_fd_sc_hd__nand3_4 _39270_ (.A(_08736_),
    .B(_08737_),
    .C(_08739_),
    .Y(_08741_));
 sky130_fd_sc_hd__a21boi_4 _39271_ (.A1(_08509_),
    .A2(_08513_),
    .B1_N(_08511_),
    .Y(_08742_));
 sky130_fd_sc_hd__a21boi_4 _39272_ (.A1(_08740_),
    .A2(_08741_),
    .B1_N(_08742_),
    .Y(_08743_));
 sky130_vsdinv _39273_ (.A(_08742_),
    .Y(_08744_));
 sky130_fd_sc_hd__nand3_4 _39274_ (.A(_08744_),
    .B(_08741_),
    .C(_08740_),
    .Y(_08745_));
 sky130_vsdinv _39275_ (.A(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__nor2_4 _39276_ (.A(_08743_),
    .B(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__buf_1 _39277_ (.A(_03353_),
    .X(_08748_));
 sky130_fd_sc_hd__buf_1 _39278_ (.A(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__nand2_4 _39279_ (.A(_08749_),
    .B(_07154_),
    .Y(_08750_));
 sky130_fd_sc_hd__o21ai_4 _39280_ (.A1(_03359_),
    .A2(_07619_),
    .B1(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__buf_1 _39281_ (.A(_08313_),
    .X(_08752_));
 sky130_fd_sc_hd__buf_1 _39282_ (.A(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__buf_1 _39283_ (.A(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__buf_1 _39284_ (.A(_08530_),
    .X(_08755_));
 sky130_fd_sc_hd__buf_1 _39285_ (.A(_08755_),
    .X(_08756_));
 sky130_fd_sc_hd__nand4_4 _39286_ (.A(_08754_),
    .B(_08756_),
    .C(_03436_),
    .D(_05940_),
    .Y(_08757_));
 sky130_fd_sc_hd__buf_1 _39287_ (.A(\pcpi_mul.rs1[23] ),
    .X(_08758_));
 sky130_fd_sc_hd__buf_1 _39288_ (.A(_08758_),
    .X(_08759_));
 sky130_fd_sc_hd__buf_1 _39289_ (.A(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__nand2_4 _39290_ (.A(_08760_),
    .B(_03420_),
    .Y(_08761_));
 sky130_vsdinv _39291_ (.A(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__a21oi_4 _39292_ (.A1(_08751_),
    .A2(_08757_),
    .B1(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__nand3_4 _39293_ (.A(_08751_),
    .B(_08757_),
    .C(_08762_),
    .Y(_08764_));
 sky130_vsdinv _39294_ (.A(_08764_),
    .Y(_08765_));
 sky130_fd_sc_hd__nor2_4 _39295_ (.A(_08763_),
    .B(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__nand2_4 _39296_ (.A(_08747_),
    .B(_08766_),
    .Y(_08767_));
 sky130_vsdinv _39297_ (.A(_08766_),
    .Y(_08768_));
 sky130_fd_sc_hd__o21ai_4 _39298_ (.A1(_08743_),
    .A2(_08746_),
    .B1(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__nand2_4 _39299_ (.A(_08767_),
    .B(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__a21o_4 _39300_ (.A1(_08519_),
    .A2(_08538_),
    .B1(_08770_),
    .X(_08771_));
 sky130_fd_sc_hd__nand3_4 _39301_ (.A(_08770_),
    .B(_08519_),
    .C(_08538_),
    .Y(_08772_));
 sky130_fd_sc_hd__nand2_4 _39302_ (.A(_08771_),
    .B(_08772_),
    .Y(_08773_));
 sky130_fd_sc_hd__a21boi_4 _39303_ (.A1(_08525_),
    .A2(_08533_),
    .B1_N(_08529_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand2_4 _39304_ (.A(_08773_),
    .B(_08774_),
    .Y(_08775_));
 sky130_vsdinv _39305_ (.A(_08774_),
    .Y(_08776_));
 sky130_fd_sc_hd__nand3_4 _39306_ (.A(_08771_),
    .B(_08772_),
    .C(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__nand2_4 _39307_ (.A(_08775_),
    .B(_08777_),
    .Y(_08778_));
 sky130_fd_sc_hd__nand2_4 _39308_ (.A(_08730_),
    .B(_08778_),
    .Y(_08779_));
 sky130_fd_sc_hd__nand4_4 _39309_ (.A(_08777_),
    .B(_08727_),
    .C(_08729_),
    .D(_08775_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand2_4 _39310_ (.A(_08779_),
    .B(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__nand2_4 _39311_ (.A(_08781_),
    .B(_08625_),
    .Y(_08782_));
 sky130_vsdinv _39312_ (.A(_08625_),
    .Y(_08783_));
 sky130_fd_sc_hd__nand3_4 _39313_ (.A(_08779_),
    .B(_08780_),
    .C(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__nand2_4 _39314_ (.A(_08782_),
    .B(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__a21boi_4 _39315_ (.A1(_08553_),
    .A2(_08502_),
    .B1_N(_08503_),
    .Y(_08786_));
 sky130_fd_sc_hd__nand2_4 _39316_ (.A(_08785_),
    .B(_08786_),
    .Y(_08787_));
 sky130_vsdinv _39317_ (.A(_08786_),
    .Y(_08788_));
 sky130_fd_sc_hd__nand3_4 _39318_ (.A(_08782_),
    .B(_08788_),
    .C(_08784_),
    .Y(_08789_));
 sky130_fd_sc_hd__nand2_4 _39319_ (.A(_08787_),
    .B(_08789_),
    .Y(_08790_));
 sky130_vsdinv _39320_ (.A(_08641_),
    .Y(_08791_));
 sky130_fd_sc_hd__a21boi_4 _39321_ (.A1(_08645_),
    .A2(_08791_),
    .B1_N(_08648_),
    .Y(_08792_));
 sky130_vsdinv _39322_ (.A(_08792_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand2_4 _39323_ (.A(_06937_),
    .B(_03540_),
    .Y(_08794_));
 sky130_fd_sc_hd__buf_1 _39324_ (.A(_03534_),
    .X(_08795_));
 sky130_fd_sc_hd__nand2_4 _39325_ (.A(_06941_),
    .B(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__nand2_4 _39326_ (.A(_08794_),
    .B(_08796_),
    .Y(_08797_));
 sky130_fd_sc_hd__nand4_4 _39327_ (.A(_06084_),
    .B(_06339_),
    .C(_07553_),
    .D(_07556_),
    .Y(_08798_));
 sky130_fd_sc_hd__nand2_4 _39328_ (.A(_07761_),
    .B(_03529_),
    .Y(_08799_));
 sky130_vsdinv _39329_ (.A(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__nand3_4 _39330_ (.A(_08797_),
    .B(_08798_),
    .C(_08800_),
    .Y(_08801_));
 sky130_fd_sc_hd__nand2_4 _39331_ (.A(_08797_),
    .B(_08798_),
    .Y(_08802_));
 sky130_fd_sc_hd__nand2_4 _39332_ (.A(_08802_),
    .B(_08799_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand3_4 _39333_ (.A(_08793_),
    .B(_08801_),
    .C(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__nand2_4 _39334_ (.A(_08803_),
    .B(_08801_),
    .Y(_08805_));
 sky130_fd_sc_hd__nand2_4 _39335_ (.A(_08805_),
    .B(_08792_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand2_4 _39336_ (.A(_08804_),
    .B(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__a21boi_4 _39337_ (.A1(_08570_),
    .A2(_08575_),
    .B1_N(_08573_),
    .Y(_08808_));
 sky130_fd_sc_hd__nand2_4 _39338_ (.A(_08807_),
    .B(_08808_),
    .Y(_08809_));
 sky130_vsdinv _39339_ (.A(_08808_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand3_4 _39340_ (.A(_08804_),
    .B(_08806_),
    .C(_08810_),
    .Y(_08811_));
 sky130_fd_sc_hd__nand2_4 _39341_ (.A(_08809_),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__a21boi_4 _39342_ (.A1(_08580_),
    .A2(_08586_),
    .B1_N(_08582_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_4 _39343_ (.A(_08812_),
    .B(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__nand2_4 _39344_ (.A(_08587_),
    .B(_08582_),
    .Y(_08815_));
 sky130_fd_sc_hd__nand3_4 _39345_ (.A(_08815_),
    .B(_08809_),
    .C(_08811_),
    .Y(_08816_));
 sky130_fd_sc_hd__nand2_4 _39346_ (.A(_08814_),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__nand2_4 _39347_ (.A(_07753_),
    .B(_07734_),
    .Y(_08818_));
 sky130_fd_sc_hd__nand2_4 _39348_ (.A(_06455_),
    .B(_07737_),
    .Y(_08819_));
 sky130_fd_sc_hd__nand2_4 _39349_ (.A(_08818_),
    .B(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__nand4_4 _39350_ (.A(_06564_),
    .B(_07654_),
    .C(_07518_),
    .D(_07187_),
    .Y(_08821_));
 sky130_fd_sc_hd__nand2_4 _39351_ (.A(_06571_),
    .B(_03512_),
    .Y(_08822_));
 sky130_vsdinv _39352_ (.A(_08822_),
    .Y(_08823_));
 sky130_fd_sc_hd__nand3_4 _39353_ (.A(_08820_),
    .B(_08821_),
    .C(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__a21o_4 _39354_ (.A1(_08820_),
    .A2(_08821_),
    .B1(_08823_),
    .X(_08825_));
 sky130_fd_sc_hd__nand2_4 _39355_ (.A(_08599_),
    .B(_08593_),
    .Y(_08826_));
 sky130_fd_sc_hd__a21oi_4 _39356_ (.A1(_08824_),
    .A2(_08825_),
    .B1(_08826_),
    .Y(_08827_));
 sky130_vsdinv _39357_ (.A(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__nand3_4 _39358_ (.A(_08826_),
    .B(_08824_),
    .C(_08825_),
    .Y(_08829_));
 sky130_fd_sc_hd__nand2_4 _39359_ (.A(_08470_),
    .B(_06751_),
    .Y(_08830_));
 sky130_vsdinv _39360_ (.A(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__nand2_4 _39361_ (.A(_06995_),
    .B(_07543_),
    .Y(_08832_));
 sky130_fd_sc_hd__nand2_4 _39362_ (.A(_06852_),
    .B(_07541_),
    .Y(_08833_));
 sky130_fd_sc_hd__nand2_4 _39363_ (.A(_08832_),
    .B(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__buf_1 _39364_ (.A(_06711_),
    .X(_08835_));
 sky130_fd_sc_hd__nand4_4 _39365_ (.A(_08835_),
    .B(_07005_),
    .C(_06891_),
    .D(_07668_),
    .Y(_08836_));
 sky130_fd_sc_hd__nand2_4 _39366_ (.A(_08834_),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__xor2_4 _39367_ (.A(_08831_),
    .B(_08837_),
    .X(_08838_));
 sky130_vsdinv _39368_ (.A(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__a21oi_4 _39369_ (.A1(_08828_),
    .A2(_08829_),
    .B1(_08839_),
    .Y(_08840_));
 sky130_vsdinv _39370_ (.A(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__nand3_4 _39371_ (.A(_08828_),
    .B(_08839_),
    .C(_08829_),
    .Y(_08842_));
 sky130_fd_sc_hd__nand2_4 _39372_ (.A(_08841_),
    .B(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__nand2_4 _39373_ (.A(_08817_),
    .B(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__nand4_4 _39374_ (.A(_08842_),
    .B(_08814_),
    .C(_08841_),
    .D(_08816_),
    .Y(_08845_));
 sky130_fd_sc_hd__nand2_4 _39375_ (.A(_08844_),
    .B(_08845_),
    .Y(_08846_));
 sky130_fd_sc_hd__nand2_4 _39376_ (.A(_08651_),
    .B(_08628_),
    .Y(_08847_));
 sky130_fd_sc_hd__nand2_4 _39377_ (.A(_08846_),
    .B(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nand4_4 _39378_ (.A(_08628_),
    .B(_08844_),
    .C(_08845_),
    .D(_08651_),
    .Y(_08849_));
 sky130_fd_sc_hd__nand2_4 _39379_ (.A(_08848_),
    .B(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__a21boi_4 _39380_ (.A1(_08590_),
    .A2(_08617_),
    .B1_N(_08592_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand2_4 _39381_ (.A(_08850_),
    .B(_08851_),
    .Y(_08852_));
 sky130_vsdinv _39382_ (.A(_08851_),
    .Y(_08853_));
 sky130_fd_sc_hd__nand3_4 _39383_ (.A(_08848_),
    .B(_08849_),
    .C(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_4 _39384_ (.A(_08852_),
    .B(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__nand2_4 _39385_ (.A(_08650_),
    .B(_08639_),
    .Y(_08856_));
 sky130_fd_sc_hd__buf_1 _39386_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08857_));
 sky130_fd_sc_hd__nand2_4 _39387_ (.A(_03248_),
    .B(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__buf_1 _39388_ (.A(\pcpi_mul.rs1[0] ),
    .X(_08859_));
 sky130_fd_sc_hd__nand2_4 _39389_ (.A(_08859_),
    .B(_03575_),
    .Y(_08860_));
 sky130_fd_sc_hd__nand2_4 _39390_ (.A(_08858_),
    .B(_08860_),
    .Y(_08861_));
 sky130_fd_sc_hd__buf_1 _39391_ (.A(_03574_),
    .X(_08862_));
 sky130_fd_sc_hd__nand4_4 _39392_ (.A(_08859_),
    .B(_03248_),
    .C(_08857_),
    .D(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__nand2_4 _39393_ (.A(_06054_),
    .B(_03562_),
    .Y(_08864_));
 sky130_vsdinv _39394_ (.A(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__a21o_4 _39395_ (.A1(_08861_),
    .A2(_08863_),
    .B1(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__nand3_4 _39396_ (.A(_08861_),
    .B(_08863_),
    .C(_08865_),
    .Y(_08867_));
 sky130_fd_sc_hd__nor2_4 _39397_ (.A(_08633_),
    .B(_08637_),
    .Y(_08868_));
 sky130_fd_sc_hd__a21oi_4 _39398_ (.A1(_08866_),
    .A2(_08867_),
    .B1(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__nand3_4 _39399_ (.A(_08866_),
    .B(_08868_),
    .C(_08867_),
    .Y(_08870_));
 sky130_vsdinv _39400_ (.A(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__nor2_4 _39401_ (.A(_08869_),
    .B(_08871_),
    .Y(_08872_));
 sky130_fd_sc_hd__buf_1 _39402_ (.A(\pcpi_mul.rs2[18] ),
    .X(_08873_));
 sky130_fd_sc_hd__nand2_4 _39403_ (.A(_06159_),
    .B(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__buf_1 _39404_ (.A(\pcpi_mul.rs2[20] ),
    .X(_08875_));
 sky130_fd_sc_hd__nand2_4 _39405_ (.A(_05942_),
    .B(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__nand2_4 _39406_ (.A(_06222_),
    .B(_08190_),
    .Y(_08877_));
 sky130_fd_sc_hd__nand2_4 _39407_ (.A(_08876_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__nand4_4 _39408_ (.A(_06226_),
    .B(_05951_),
    .C(_08646_),
    .D(_08197_),
    .Y(_08879_));
 sky130_fd_sc_hd__nand2_4 _39409_ (.A(_08878_),
    .B(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__xor2_4 _39410_ (.A(_08874_),
    .B(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__nand2_4 _39411_ (.A(_08872_),
    .B(_08881_),
    .Y(_08882_));
 sky130_vsdinv _39412_ (.A(_08881_),
    .Y(_08883_));
 sky130_fd_sc_hd__o21ai_4 _39413_ (.A1(_08869_),
    .A2(_08871_),
    .B1(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__nand2_4 _39414_ (.A(_08882_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__xor2_4 _39415_ (.A(_08856_),
    .B(_08885_),
    .X(_08886_));
 sky130_vsdinv _39416_ (.A(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__nand2_4 _39417_ (.A(_08855_),
    .B(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__nand3_4 _39418_ (.A(_08852_),
    .B(_08854_),
    .C(_08886_),
    .Y(_08889_));
 sky130_fd_sc_hd__nand2_4 _39419_ (.A(_08888_),
    .B(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__nand2_4 _39420_ (.A(_08890_),
    .B(_08655_),
    .Y(_08891_));
 sky130_vsdinv _39421_ (.A(_08655_),
    .Y(_08892_));
 sky130_fd_sc_hd__nand3_4 _39422_ (.A(_08888_),
    .B(_08892_),
    .C(_08889_),
    .Y(_08893_));
 sky130_fd_sc_hd__nand2_4 _39423_ (.A(_08891_),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__nand2_4 _39424_ (.A(_08790_),
    .B(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__nand4_4 _39425_ (.A(_08789_),
    .B(_08787_),
    .C(_08891_),
    .D(_08893_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand2_4 _39426_ (.A(_08895_),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__nand2_4 _39427_ (.A(_08695_),
    .B(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__nand3_4 _39428_ (.A(_08694_),
    .B(_08896_),
    .C(_08895_),
    .Y(_08899_));
 sky130_fd_sc_hd__nand2_4 _39429_ (.A(_08898_),
    .B(_08899_),
    .Y(_08900_));
 sky130_fd_sc_hd__a21boi_4 _39430_ (.A1(_08543_),
    .A2(_08549_),
    .B1_N(_08545_),
    .Y(_08901_));
 sky130_fd_sc_hd__nand2_4 _39431_ (.A(_08563_),
    .B(_08558_),
    .Y(_08902_));
 sky130_fd_sc_hd__xor2_4 _39432_ (.A(_08901_),
    .B(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__nand2_4 _39433_ (.A(_08900_),
    .B(_08903_),
    .Y(_08904_));
 sky130_vsdinv _39434_ (.A(_08903_),
    .Y(_08905_));
 sky130_fd_sc_hd__nand3_4 _39435_ (.A(_08905_),
    .B(_08898_),
    .C(_08899_),
    .Y(_08906_));
 sky130_fd_sc_hd__nand2_4 _39436_ (.A(_08904_),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__a21oi_4 _39437_ (.A1(_08662_),
    .A2(_08663_),
    .B1(_08468_),
    .Y(_08908_));
 sky130_fd_sc_hd__o21ai_4 _39438_ (.A1(_08670_),
    .A2(_08908_),
    .B1(_08666_),
    .Y(_08909_));
 sky130_vsdinv _39439_ (.A(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__nand2_4 _39440_ (.A(_08907_),
    .B(_08910_),
    .Y(_08911_));
 sky130_fd_sc_hd__nand3_4 _39441_ (.A(_08904_),
    .B(_08909_),
    .C(_08906_),
    .Y(_08912_));
 sky130_fd_sc_hd__nand2_4 _39442_ (.A(_08911_),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__a21oi_4 _39443_ (.A1(_08349_),
    .A2(_08344_),
    .B1(_08668_),
    .Y(_08914_));
 sky130_vsdinv _39444_ (.A(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__nand2_4 _39445_ (.A(_08913_),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand3_4 _39446_ (.A(_08911_),
    .B(_08914_),
    .C(_08912_),
    .Y(_08917_));
 sky130_fd_sc_hd__nand3_4 _39447_ (.A(_08693_),
    .B(_08916_),
    .C(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand2_4 _39448_ (.A(_08916_),
    .B(_08917_),
    .Y(_08919_));
 sky130_fd_sc_hd__nand2_4 _39449_ (.A(_08919_),
    .B(_08692_),
    .Y(_08920_));
 sky130_fd_sc_hd__and2_4 _39450_ (.A(_08918_),
    .B(_08920_),
    .X(_08921_));
 sky130_vsdinv _39451_ (.A(_08686_),
    .Y(_08922_));
 sky130_fd_sc_hd__a21oi_4 _39452_ (.A1(_08691_),
    .A2(_08684_),
    .B1(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__xnor2_4 _39453_ (.A(_08921_),
    .B(_08923_),
    .Y(_01428_));
 sky130_vsdinv _39454_ (.A(_08874_),
    .Y(_08924_));
 sky130_fd_sc_hd__a21boi_4 _39455_ (.A1(_08878_),
    .A2(_08924_),
    .B1_N(_08879_),
    .Y(_08925_));
 sky130_vsdinv _39456_ (.A(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__nand2_4 _39457_ (.A(_06941_),
    .B(_08124_),
    .Y(_08927_));
 sky130_fd_sc_hd__buf_1 _39458_ (.A(\pcpi_mul.rs1[8] ),
    .X(_08928_));
 sky130_fd_sc_hd__nand2_4 _39459_ (.A(_08928_),
    .B(_08127_),
    .Y(_08929_));
 sky130_fd_sc_hd__nand2_4 _39460_ (.A(_08927_),
    .B(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__nand4_4 _39461_ (.A(_06339_),
    .B(_06342_),
    .C(_03535_),
    .D(_07716_),
    .Y(_08931_));
 sky130_fd_sc_hd__nand2_4 _39462_ (.A(_07464_),
    .B(_03529_),
    .Y(_08932_));
 sky130_vsdinv _39463_ (.A(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__nand3_4 _39464_ (.A(_08930_),
    .B(_08931_),
    .C(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand2_4 _39465_ (.A(_08930_),
    .B(_08931_),
    .Y(_08935_));
 sky130_fd_sc_hd__nand2_4 _39466_ (.A(_08935_),
    .B(_08932_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand3_4 _39467_ (.A(_08926_),
    .B(_08934_),
    .C(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__nand2_4 _39468_ (.A(_08936_),
    .B(_08934_),
    .Y(_08938_));
 sky130_fd_sc_hd__nand2_4 _39469_ (.A(_08938_),
    .B(_08925_),
    .Y(_08939_));
 sky130_fd_sc_hd__nand2_4 _39470_ (.A(_08937_),
    .B(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__a21boi_4 _39471_ (.A1(_08797_),
    .A2(_08800_),
    .B1_N(_08798_),
    .Y(_08941_));
 sky130_fd_sc_hd__nand2_4 _39472_ (.A(_08940_),
    .B(_08941_),
    .Y(_08942_));
 sky130_vsdinv _39473_ (.A(_08941_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand3_4 _39474_ (.A(_08937_),
    .B(_08939_),
    .C(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__nand2_4 _39475_ (.A(_08942_),
    .B(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__a21boi_4 _39476_ (.A1(_08806_),
    .A2(_08810_),
    .B1_N(_08804_),
    .Y(_08946_));
 sky130_fd_sc_hd__nand2_4 _39477_ (.A(_08945_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__nand2_4 _39478_ (.A(_08811_),
    .B(_08804_),
    .Y(_08948_));
 sky130_fd_sc_hd__nand3_4 _39479_ (.A(_08948_),
    .B(_08944_),
    .C(_08942_),
    .Y(_08949_));
 sky130_fd_sc_hd__nand2_4 _39480_ (.A(_08947_),
    .B(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__a21boi_4 _39481_ (.A1(_08820_),
    .A2(_08823_),
    .B1_N(_08821_),
    .Y(_08951_));
 sky130_fd_sc_hd__nand2_4 _39482_ (.A(_06454_),
    .B(_07733_),
    .Y(_08952_));
 sky130_fd_sc_hd__buf_1 _39483_ (.A(\pcpi_mul.rs2[13] ),
    .X(_08953_));
 sky130_fd_sc_hd__nand2_4 _39484_ (.A(_08606_),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_4 _39485_ (.A(_08952_),
    .B(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__nand4_4 _39486_ (.A(_06454_),
    .B(_08606_),
    .C(_03516_),
    .D(_07361_),
    .Y(_08956_));
 sky130_fd_sc_hd__nand2_4 _39487_ (.A(_08955_),
    .B(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__nand2_4 _39488_ (.A(_03302_),
    .B(_03511_),
    .Y(_08958_));
 sky130_fd_sc_hd__nand2_4 _39489_ (.A(_08957_),
    .B(_08958_),
    .Y(_08959_));
 sky130_vsdinv _39490_ (.A(_08958_),
    .Y(_08960_));
 sky130_fd_sc_hd__nand3_4 _39491_ (.A(_08955_),
    .B(_08956_),
    .C(_08960_),
    .Y(_08961_));
 sky130_fd_sc_hd__nand2_4 _39492_ (.A(_08959_),
    .B(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__nor2_4 _39493_ (.A(_08951_),
    .B(_08962_),
    .Y(_08963_));
 sky130_vsdinv _39494_ (.A(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand2_4 _39495_ (.A(_08962_),
    .B(_08951_),
    .Y(_08965_));
 sky130_fd_sc_hd__buf_1 _39496_ (.A(_07156_),
    .X(_08966_));
 sky130_fd_sc_hd__nand2_4 _39497_ (.A(_08966_),
    .B(_03495_),
    .Y(_08967_));
 sky130_fd_sc_hd__nand2_4 _39498_ (.A(_06852_),
    .B(_07543_),
    .Y(_08968_));
 sky130_fd_sc_hd__nand2_4 _39499_ (.A(_03314_),
    .B(_07541_),
    .Y(_08969_));
 sky130_fd_sc_hd__nand2_4 _39500_ (.A(_08968_),
    .B(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__buf_1 _39501_ (.A(_03310_),
    .X(_08971_));
 sky130_fd_sc_hd__nand4_4 _39502_ (.A(_08971_),
    .B(_08470_),
    .C(_06891_),
    .D(_07344_),
    .Y(_08972_));
 sky130_fd_sc_hd__nand2_4 _39503_ (.A(_08970_),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__xor2_4 _39504_ (.A(_08967_),
    .B(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__a21o_4 _39505_ (.A1(_08964_),
    .A2(_08965_),
    .B1(_08974_),
    .X(_08975_));
 sky130_fd_sc_hd__nand3_4 _39506_ (.A(_08964_),
    .B(_08974_),
    .C(_08965_),
    .Y(_08976_));
 sky130_fd_sc_hd__nand2_4 _39507_ (.A(_08975_),
    .B(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__nand2_4 _39508_ (.A(_08950_),
    .B(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__nand4_4 _39509_ (.A(_08976_),
    .B(_08947_),
    .C(_08975_),
    .D(_08949_),
    .Y(_08979_));
 sky130_fd_sc_hd__nand2_4 _39510_ (.A(_08978_),
    .B(_08979_),
    .Y(_08980_));
 sky130_vsdinv _39511_ (.A(_08856_),
    .Y(_08981_));
 sky130_fd_sc_hd__nand3_4 _39512_ (.A(_08882_),
    .B(_08884_),
    .C(_08981_),
    .Y(_08982_));
 sky130_fd_sc_hd__nand2_4 _39513_ (.A(_08980_),
    .B(_08982_),
    .Y(_08983_));
 sky130_vsdinv _39514_ (.A(_08982_),
    .Y(_08984_));
 sky130_fd_sc_hd__nand3_4 _39515_ (.A(_08978_),
    .B(_08979_),
    .C(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__nand2_4 _39516_ (.A(_08983_),
    .B(_08985_),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_4 _39517_ (.A(_08845_),
    .B(_08816_),
    .Y(_08987_));
 sky130_vsdinv _39518_ (.A(_08987_),
    .Y(_08988_));
 sky130_fd_sc_hd__nand2_4 _39519_ (.A(_08986_),
    .B(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__nand3_4 _39520_ (.A(_08983_),
    .B(_08987_),
    .C(_08985_),
    .Y(_08990_));
 sky130_fd_sc_hd__buf_1 _39521_ (.A(_05883_),
    .X(_08991_));
 sky130_fd_sc_hd__nand2_4 _39522_ (.A(_08991_),
    .B(_03575_),
    .Y(_08992_));
 sky130_fd_sc_hd__nand2_4 _39523_ (.A(_06054_),
    .B(_08857_),
    .Y(_08993_));
 sky130_fd_sc_hd__nand2_4 _39524_ (.A(_08992_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__buf_1 _39525_ (.A(_08629_),
    .X(_08995_));
 sky130_fd_sc_hd__nand4_4 _39526_ (.A(_08991_),
    .B(_05899_),
    .C(_08995_),
    .D(_08862_),
    .Y(_08996_));
 sky130_fd_sc_hd__nand2_4 _39527_ (.A(_06383_),
    .B(_08634_),
    .Y(_08997_));
 sky130_vsdinv _39528_ (.A(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__a21o_4 _39529_ (.A1(_08994_),
    .A2(_08996_),
    .B1(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__nand3_4 _39530_ (.A(_08994_),
    .B(_08996_),
    .C(_08998_),
    .Y(_09000_));
 sky130_fd_sc_hd__nand2_4 _39531_ (.A(_08999_),
    .B(_09000_),
    .Y(_09001_));
 sky130_fd_sc_hd__a21boi_4 _39532_ (.A1(_08861_),
    .A2(_08865_),
    .B1_N(_08863_),
    .Y(_09002_));
 sky130_fd_sc_hd__nand2_4 _39533_ (.A(_09001_),
    .B(_09002_),
    .Y(_09003_));
 sky130_vsdinv _39534_ (.A(_09002_),
    .Y(_09004_));
 sky130_fd_sc_hd__nand3_4 _39535_ (.A(_09004_),
    .B(_09000_),
    .C(_08999_),
    .Y(_09005_));
 sky130_fd_sc_hd__nand2_4 _39536_ (.A(_06243_),
    .B(_08873_),
    .Y(_09006_));
 sky130_fd_sc_hd__nand2_4 _39537_ (.A(_06222_),
    .B(_08193_),
    .Y(_09007_));
 sky130_fd_sc_hd__buf_1 _39538_ (.A(\pcpi_mul.rs2[19] ),
    .X(_09008_));
 sky130_fd_sc_hd__nand2_4 _39539_ (.A(_07525_),
    .B(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__nand2_4 _39540_ (.A(_09007_),
    .B(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__nand4_4 _39541_ (.A(_05951_),
    .B(_07525_),
    .C(_08190_),
    .D(_08875_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_4 _39542_ (.A(_09010_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__xor2_4 _39543_ (.A(_09006_),
    .B(_09012_),
    .X(_09013_));
 sky130_fd_sc_hd__a21o_4 _39544_ (.A1(_09003_),
    .A2(_09005_),
    .B1(_09013_),
    .X(_09014_));
 sky130_fd_sc_hd__nand3_4 _39545_ (.A(_09003_),
    .B(_09013_),
    .C(_09005_),
    .Y(_09015_));
 sky130_fd_sc_hd__o21ai_4 _39546_ (.A1(_08869_),
    .A2(_08883_),
    .B1(_08870_),
    .Y(_09016_));
 sky130_fd_sc_hd__a21o_4 _39547_ (.A1(_09014_),
    .A2(_09015_),
    .B1(_09016_),
    .X(_09017_));
 sky130_fd_sc_hd__nand3_4 _39548_ (.A(_09016_),
    .B(_09015_),
    .C(_09014_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand2_4 _39549_ (.A(_05587_),
    .B(_03584_),
    .Y(_09019_));
 sky130_vsdinv _39550_ (.A(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__a21oi_4 _39551_ (.A1(_09017_),
    .A2(_09018_),
    .B1(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__nand3_4 _39552_ (.A(_09017_),
    .B(_09020_),
    .C(_09018_),
    .Y(_09022_));
 sky130_vsdinv _39553_ (.A(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__nor2_4 _39554_ (.A(_09021_),
    .B(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__a21oi_4 _39555_ (.A1(_08989_),
    .A2(_08990_),
    .B1(_09024_),
    .Y(_09025_));
 sky130_fd_sc_hd__nand3_4 _39556_ (.A(_08989_),
    .B(_09024_),
    .C(_08990_),
    .Y(_09026_));
 sky130_vsdinv _39557_ (.A(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__o21ai_4 _39558_ (.A1(_09025_),
    .A2(_09027_),
    .B1(_08889_),
    .Y(_09028_));
 sky130_fd_sc_hd__a21o_4 _39559_ (.A1(_08989_),
    .A2(_08990_),
    .B1(_09024_),
    .X(_09029_));
 sky130_vsdinv _39560_ (.A(_08889_),
    .Y(_09030_));
 sky130_fd_sc_hd__nand3_4 _39561_ (.A(_09029_),
    .B(_09030_),
    .C(_09026_),
    .Y(_09031_));
 sky130_fd_sc_hd__nand2_4 _39562_ (.A(_09028_),
    .B(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__a21bo_4 _39563_ (.A1(_08831_),
    .A2(_08834_),
    .B1_N(_08836_),
    .X(_09033_));
 sky130_fd_sc_hd__nand2_4 _39564_ (.A(_03324_),
    .B(_06593_),
    .Y(_09034_));
 sky130_fd_sc_hd__nand2_4 _39565_ (.A(_07874_),
    .B(_06599_),
    .Y(_09035_));
 sky130_fd_sc_hd__nand2_4 _39566_ (.A(_09034_),
    .B(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__buf_1 _39567_ (.A(_03323_),
    .X(_09037_));
 sky130_fd_sc_hd__buf_1 _39568_ (.A(_07442_),
    .X(_09038_));
 sky130_fd_sc_hd__nand4_4 _39569_ (.A(_09037_),
    .B(_09038_),
    .C(_08259_),
    .D(_08257_),
    .Y(_09039_));
 sky130_fd_sc_hd__nand2_4 _39570_ (.A(_03336_),
    .B(_06605_),
    .Y(_09040_));
 sky130_vsdinv _39571_ (.A(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__nand3_4 _39572_ (.A(_09036_),
    .B(_09039_),
    .C(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__nand2_4 _39573_ (.A(_09036_),
    .B(_09039_),
    .Y(_09043_));
 sky130_fd_sc_hd__nand2_4 _39574_ (.A(_09043_),
    .B(_09040_),
    .Y(_09044_));
 sky130_fd_sc_hd__nand3_4 _39575_ (.A(_09033_),
    .B(_09042_),
    .C(_09044_),
    .Y(_09045_));
 sky130_fd_sc_hd__nand2_4 _39576_ (.A(_09044_),
    .B(_09042_),
    .Y(_09046_));
 sky130_fd_sc_hd__a21boi_4 _39577_ (.A1(_08834_),
    .A2(_08831_),
    .B1_N(_08836_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_4 _39578_ (.A(_09046_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__nand2_4 _39579_ (.A(_09045_),
    .B(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__a21boi_4 _39580_ (.A1(_08698_),
    .A2(_08701_),
    .B1_N(_08699_),
    .Y(_09050_));
 sky130_fd_sc_hd__nand2_4 _39581_ (.A(_09049_),
    .B(_09050_),
    .Y(_09051_));
 sky130_vsdinv _39582_ (.A(_09050_),
    .Y(_09052_));
 sky130_fd_sc_hd__nand3_4 _39583_ (.A(_09045_),
    .B(_09048_),
    .C(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__nand2_4 _39584_ (.A(_09051_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__o21a_4 _39585_ (.A1(_08838_),
    .A2(_08827_),
    .B1(_08829_),
    .X(_09055_));
 sky130_fd_sc_hd__nand2_4 _39586_ (.A(_09054_),
    .B(_09055_),
    .Y(_09056_));
 sky130_fd_sc_hd__o21ai_4 _39587_ (.A1(_08838_),
    .A2(_08827_),
    .B1(_08829_),
    .Y(_09057_));
 sky130_fd_sc_hd__nand3_4 _39588_ (.A(_09057_),
    .B(_09053_),
    .C(_09051_),
    .Y(_09058_));
 sky130_fd_sc_hd__nand2_4 _39589_ (.A(_09056_),
    .B(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__a21boi_4 _39590_ (.A1(_08707_),
    .A2(_08713_),
    .B1_N(_08709_),
    .Y(_09060_));
 sky130_fd_sc_hd__nand2_4 _39591_ (.A(_09059_),
    .B(_09060_),
    .Y(_09061_));
 sky130_vsdinv _39592_ (.A(_09060_),
    .Y(_09062_));
 sky130_fd_sc_hd__nand3_4 _39593_ (.A(_09056_),
    .B(_09058_),
    .C(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_4 _39594_ (.A(_09061_),
    .B(_09063_),
    .Y(_09064_));
 sky130_fd_sc_hd__a21boi_4 _39595_ (.A1(_08717_),
    .A2(_08723_),
    .B1_N(_08719_),
    .Y(_09065_));
 sky130_fd_sc_hd__nand2_4 _39596_ (.A(_09064_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__nand2_4 _39597_ (.A(_08724_),
    .B(_08719_),
    .Y(_09067_));
 sky130_fd_sc_hd__nand3_4 _39598_ (.A(_09067_),
    .B(_09063_),
    .C(_09061_),
    .Y(_09068_));
 sky130_fd_sc_hd__nand2_4 _39599_ (.A(_09066_),
    .B(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__buf_1 _39600_ (.A(_08045_),
    .X(_09070_));
 sky130_fd_sc_hd__nand2_4 _39601_ (.A(_09070_),
    .B(_08731_),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_4 _39602_ (.A(_08308_),
    .B(_07131_),
    .Y(_09072_));
 sky130_fd_sc_hd__nand2_4 _39603_ (.A(_09071_),
    .B(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__buf_1 _39604_ (.A(_08054_),
    .X(_09074_));
 sky130_fd_sc_hd__nand4_4 _39605_ (.A(_08046_),
    .B(_09074_),
    .C(_08734_),
    .D(_08731_),
    .Y(_09075_));
 sky130_fd_sc_hd__nand2_4 _39606_ (.A(_08748_),
    .B(_06327_),
    .Y(_09076_));
 sky130_vsdinv _39607_ (.A(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__nand3_4 _39608_ (.A(_09073_),
    .B(_09075_),
    .C(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__a21o_4 _39609_ (.A1(_09073_),
    .A2(_09075_),
    .B1(_09077_),
    .X(_09079_));
 sky130_fd_sc_hd__a21boi_4 _39610_ (.A1(_08736_),
    .A2(_08739_),
    .B1_N(_08737_),
    .Y(_09080_));
 sky130_vsdinv _39611_ (.A(_09080_),
    .Y(_09081_));
 sky130_fd_sc_hd__a21o_4 _39612_ (.A1(_09078_),
    .A2(_09079_),
    .B1(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__nand3_4 _39613_ (.A(_09081_),
    .B(_09078_),
    .C(_09079_),
    .Y(_09083_));
 sky130_fd_sc_hd__nand2_4 _39614_ (.A(_03357_),
    .B(_05909_),
    .Y(_09084_));
 sky130_fd_sc_hd__o21ai_4 _39615_ (.A1(_03362_),
    .A2(_07618_),
    .B1(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__buf_1 _39616_ (.A(\pcpi_mul.rs1[22] ),
    .X(_09086_));
 sky130_fd_sc_hd__buf_1 _39617_ (.A(_09086_),
    .X(_09087_));
 sky130_fd_sc_hd__buf_1 _39618_ (.A(_08758_),
    .X(_09088_));
 sky130_fd_sc_hd__nand4_4 _39619_ (.A(_09087_),
    .B(_09088_),
    .C(_07001_),
    .D(_06705_),
    .Y(_09089_));
 sky130_fd_sc_hd__buf_1 _39620_ (.A(\pcpi_mul.rs1[24] ),
    .X(_09090_));
 sky130_fd_sc_hd__nand2_4 _39621_ (.A(_09090_),
    .B(_06853_),
    .Y(_09091_));
 sky130_vsdinv _39622_ (.A(_09091_),
    .Y(_09092_));
 sky130_fd_sc_hd__a21o_4 _39623_ (.A1(_09085_),
    .A2(_09089_),
    .B1(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__nand3_4 _39624_ (.A(_09085_),
    .B(_09089_),
    .C(_09092_),
    .Y(_09094_));
 sky130_fd_sc_hd__and2_4 _39625_ (.A(_09093_),
    .B(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__buf_1 _39626_ (.A(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__a21o_4 _39627_ (.A1(_09082_),
    .A2(_09083_),
    .B1(_09096_),
    .X(_09097_));
 sky130_fd_sc_hd__nand3_4 _39628_ (.A(_09082_),
    .B(_09096_),
    .C(_09083_),
    .Y(_09098_));
 sky130_fd_sc_hd__nand2_4 _39629_ (.A(_09097_),
    .B(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__a21o_4 _39630_ (.A1(_08745_),
    .A2(_08767_),
    .B1(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__nand3_4 _39631_ (.A(_09099_),
    .B(_08745_),
    .C(_08767_),
    .Y(_09101_));
 sky130_fd_sc_hd__nand2_4 _39632_ (.A(_09100_),
    .B(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__a21boi_4 _39633_ (.A1(_08751_),
    .A2(_08762_),
    .B1_N(_08757_),
    .Y(_09103_));
 sky130_fd_sc_hd__nand2_4 _39634_ (.A(_09102_),
    .B(_09103_),
    .Y(_09104_));
 sky130_vsdinv _39635_ (.A(_09103_),
    .Y(_09105_));
 sky130_fd_sc_hd__nand3_4 _39636_ (.A(_09100_),
    .B(_09101_),
    .C(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__nand2_4 _39637_ (.A(_09104_),
    .B(_09106_),
    .Y(_09107_));
 sky130_fd_sc_hd__nand2_4 _39638_ (.A(_09069_),
    .B(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__nand4_4 _39639_ (.A(_09106_),
    .B(_09104_),
    .C(_09066_),
    .D(_09068_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand2_4 _39640_ (.A(_09108_),
    .B(_09109_),
    .Y(_09110_));
 sky130_fd_sc_hd__a21boi_4 _39641_ (.A1(_08848_),
    .A2(_08853_),
    .B1_N(_08849_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand2_4 _39642_ (.A(_09110_),
    .B(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__nand2_4 _39643_ (.A(_08854_),
    .B(_08849_),
    .Y(_09113_));
 sky130_fd_sc_hd__nand3_4 _39644_ (.A(_09113_),
    .B(_09109_),
    .C(_09108_),
    .Y(_09114_));
 sky130_fd_sc_hd__nand2_4 _39645_ (.A(_09112_),
    .B(_09114_),
    .Y(_09115_));
 sky130_fd_sc_hd__nand2_4 _39646_ (.A(_08780_),
    .B(_08729_),
    .Y(_09116_));
 sky130_vsdinv _39647_ (.A(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__nand2_4 _39648_ (.A(_09115_),
    .B(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__nand3_4 _39649_ (.A(_09112_),
    .B(_09114_),
    .C(_09116_),
    .Y(_09119_));
 sky130_fd_sc_hd__nand2_4 _39650_ (.A(_09118_),
    .B(_09119_),
    .Y(_09120_));
 sky130_fd_sc_hd__nand2_4 _39651_ (.A(_09032_),
    .B(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__nand4_4 _39652_ (.A(_09119_),
    .B(_09028_),
    .C(_09118_),
    .D(_09031_),
    .Y(_09122_));
 sky130_fd_sc_hd__nand2_4 _39653_ (.A(_09121_),
    .B(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__nand3_4 _39654_ (.A(_09123_),
    .B(_08893_),
    .C(_08896_),
    .Y(_09124_));
 sky130_fd_sc_hd__nand2_4 _39655_ (.A(_08896_),
    .B(_08893_),
    .Y(_09125_));
 sky130_fd_sc_hd__nand3_4 _39656_ (.A(_09125_),
    .B(_09122_),
    .C(_09121_),
    .Y(_09126_));
 sky130_fd_sc_hd__nand2_4 _39657_ (.A(_09124_),
    .B(_09126_),
    .Y(_09127_));
 sky130_fd_sc_hd__a21boi_4 _39658_ (.A1(_08776_),
    .A2(_08772_),
    .B1_N(_08771_),
    .Y(_09128_));
 sky130_fd_sc_hd__nand2_4 _39659_ (.A(_08789_),
    .B(_08784_),
    .Y(_09129_));
 sky130_fd_sc_hd__xor2_4 _39660_ (.A(_09128_),
    .B(_09129_),
    .X(_09130_));
 sky130_fd_sc_hd__nand2_4 _39661_ (.A(_09127_),
    .B(_09130_),
    .Y(_09131_));
 sky130_vsdinv _39662_ (.A(_09130_),
    .Y(_09132_));
 sky130_fd_sc_hd__nand3_4 _39663_ (.A(_09124_),
    .B(_09132_),
    .C(_09126_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand2_4 _39664_ (.A(_09131_),
    .B(_09133_),
    .Y(_09134_));
 sky130_fd_sc_hd__a21boi_4 _39665_ (.A1(_08905_),
    .A2(_08898_),
    .B1_N(_08899_),
    .Y(_09135_));
 sky130_fd_sc_hd__nand2_4 _39666_ (.A(_09134_),
    .B(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__nand2_4 _39667_ (.A(_08906_),
    .B(_08899_),
    .Y(_09137_));
 sky130_fd_sc_hd__nand3_4 _39668_ (.A(_09137_),
    .B(_09133_),
    .C(_09131_),
    .Y(_09138_));
 sky130_fd_sc_hd__nand2_4 _39669_ (.A(_09136_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__a21oi_4 _39670_ (.A1(_08563_),
    .A2(_08558_),
    .B1(_08901_),
    .Y(_09140_));
 sky130_vsdinv _39671_ (.A(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__nand2_4 _39672_ (.A(_09139_),
    .B(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__nand3_4 _39673_ (.A(_09136_),
    .B(_09138_),
    .C(_09140_),
    .Y(_09143_));
 sky130_fd_sc_hd__a21oi_4 _39674_ (.A1(_08904_),
    .A2(_08906_),
    .B1(_08909_),
    .Y(_09144_));
 sky130_fd_sc_hd__o21ai_4 _39675_ (.A1(_08915_),
    .A2(_09144_),
    .B1(_08912_),
    .Y(_09145_));
 sky130_fd_sc_hd__a21oi_4 _39676_ (.A1(_09142_),
    .A2(_09143_),
    .B1(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__nand3_4 _39677_ (.A(_09142_),
    .B(_09145_),
    .C(_09143_),
    .Y(_09147_));
 sky130_vsdinv _39678_ (.A(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__nor2_4 _39679_ (.A(_09146_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__nand4_4 _39680_ (.A(_08686_),
    .B(_08918_),
    .C(_08684_),
    .D(_08920_),
    .Y(_09150_));
 sky130_fd_sc_hd__nor2_4 _39681_ (.A(_08688_),
    .B(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__and2_4 _39682_ (.A(_08243_),
    .B(_09151_),
    .X(_09152_));
 sky130_fd_sc_hd__nand2_4 _39683_ (.A(_08246_),
    .B(_09151_),
    .Y(_09153_));
 sky130_fd_sc_hd__a21boi_4 _39684_ (.A1(_08922_),
    .A2(_08920_),
    .B1_N(_08918_),
    .Y(_09154_));
 sky130_fd_sc_hd__o21a_4 _39685_ (.A1(_08690_),
    .A2(_09150_),
    .B1(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__nand2_4 _39686_ (.A(_09153_),
    .B(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__a21oi_4 _39687_ (.A1(_07414_),
    .A2(_09152_),
    .B1(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__xnor2_4 _39688_ (.A(_09149_),
    .B(_09157_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_4 _39689_ (.A(_09122_),
    .B(_09031_),
    .Y(_09158_));
 sky130_vsdinv _39690_ (.A(_08967_),
    .Y(_09159_));
 sky130_fd_sc_hd__a21bo_4 _39691_ (.A1(_09159_),
    .A2(_08970_),
    .B1_N(_08972_),
    .X(_09160_));
 sky130_fd_sc_hd__nand2_4 _39692_ (.A(_07443_),
    .B(_06481_),
    .Y(_09161_));
 sky130_fd_sc_hd__nand2_4 _39693_ (.A(_08050_),
    .B(_03480_),
    .Y(_09162_));
 sky130_fd_sc_hd__nand2_4 _39694_ (.A(_09161_),
    .B(_09162_),
    .Y(_09163_));
 sky130_fd_sc_hd__nand4_4 _39695_ (.A(_09038_),
    .B(_07629_),
    .C(_08259_),
    .D(_08257_),
    .Y(_09164_));
 sky130_fd_sc_hd__nand2_4 _39696_ (.A(_07877_),
    .B(_06605_),
    .Y(_09165_));
 sky130_vsdinv _39697_ (.A(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__nand3_4 _39698_ (.A(_09163_),
    .B(_09164_),
    .C(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__nand2_4 _39699_ (.A(_09163_),
    .B(_09164_),
    .Y(_09168_));
 sky130_fd_sc_hd__nand2_4 _39700_ (.A(_09168_),
    .B(_09165_),
    .Y(_09169_));
 sky130_fd_sc_hd__nand3_4 _39701_ (.A(_09160_),
    .B(_09167_),
    .C(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__nand2_4 _39702_ (.A(_09169_),
    .B(_09167_),
    .Y(_09171_));
 sky130_fd_sc_hd__a21boi_4 _39703_ (.A1(_08970_),
    .A2(_09159_),
    .B1_N(_08972_),
    .Y(_09172_));
 sky130_fd_sc_hd__nand2_4 _39704_ (.A(_09171_),
    .B(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__nand2_4 _39705_ (.A(_09170_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__a21boi_4 _39706_ (.A1(_09036_),
    .A2(_09041_),
    .B1_N(_09039_),
    .Y(_09175_));
 sky130_fd_sc_hd__nand2_4 _39707_ (.A(_09174_),
    .B(_09175_),
    .Y(_09176_));
 sky130_vsdinv _39708_ (.A(_09175_),
    .Y(_09177_));
 sky130_fd_sc_hd__nand3_4 _39709_ (.A(_09170_),
    .B(_09173_),
    .C(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__nand2_4 _39710_ (.A(_09176_),
    .B(_09178_),
    .Y(_09179_));
 sky130_fd_sc_hd__a21oi_4 _39711_ (.A1(_08974_),
    .A2(_08965_),
    .B1(_08963_),
    .Y(_09180_));
 sky130_fd_sc_hd__nand2_4 _39712_ (.A(_09179_),
    .B(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__a21o_4 _39713_ (.A1(_08974_),
    .A2(_08965_),
    .B1(_08963_),
    .X(_09182_));
 sky130_fd_sc_hd__nand3_4 _39714_ (.A(_09182_),
    .B(_09178_),
    .C(_09176_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_4 _39715_ (.A(_09181_),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__a21boi_4 _39716_ (.A1(_09048_),
    .A2(_09052_),
    .B1_N(_09045_),
    .Y(_09185_));
 sky130_fd_sc_hd__nand2_4 _39717_ (.A(_09184_),
    .B(_09185_),
    .Y(_09186_));
 sky130_vsdinv _39718_ (.A(_09185_),
    .Y(_09187_));
 sky130_fd_sc_hd__nand3_4 _39719_ (.A(_09181_),
    .B(_09183_),
    .C(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__nand2_4 _39720_ (.A(_09186_),
    .B(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__a21boi_4 _39721_ (.A1(_09056_),
    .A2(_09062_),
    .B1_N(_09058_),
    .Y(_09190_));
 sky130_fd_sc_hd__nand2_4 _39722_ (.A(_09189_),
    .B(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__nand2_4 _39723_ (.A(_09063_),
    .B(_09058_),
    .Y(_09192_));
 sky130_fd_sc_hd__nand3_4 _39724_ (.A(_09192_),
    .B(_09188_),
    .C(_09186_),
    .Y(_09193_));
 sky130_fd_sc_hd__nand2_4 _39725_ (.A(_09191_),
    .B(_09193_),
    .Y(_09194_));
 sky130_vsdinv _39726_ (.A(_09083_),
    .Y(_09195_));
 sky130_fd_sc_hd__a21oi_4 _39727_ (.A1(_09082_),
    .A2(_09096_),
    .B1(_09195_),
    .Y(_09196_));
 sky130_vsdinv _39728_ (.A(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__nand2_4 _39729_ (.A(_09074_),
    .B(_08505_),
    .Y(_09198_));
 sky130_fd_sc_hd__nand2_4 _39730_ (.A(_08314_),
    .B(_07131_),
    .Y(_09199_));
 sky130_fd_sc_hd__nand2_4 _39731_ (.A(_09198_),
    .B(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__nand4_4 _39732_ (.A(_09074_),
    .B(_08314_),
    .C(_08507_),
    .D(_06314_),
    .Y(_09201_));
 sky130_fd_sc_hd__buf_1 _39733_ (.A(_09086_),
    .X(_09202_));
 sky130_fd_sc_hd__nand2_4 _39734_ (.A(_09202_),
    .B(_05995_),
    .Y(_09203_));
 sky130_vsdinv _39735_ (.A(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__a21o_4 _39736_ (.A1(_09200_),
    .A2(_09201_),
    .B1(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__nand3_4 _39737_ (.A(_09200_),
    .B(_09201_),
    .C(_09204_),
    .Y(_09206_));
 sky130_fd_sc_hd__a21boi_4 _39738_ (.A1(_09073_),
    .A2(_09077_),
    .B1_N(_09075_),
    .Y(_09207_));
 sky130_fd_sc_hd__a21boi_4 _39739_ (.A1(_09205_),
    .A2(_09206_),
    .B1_N(_09207_),
    .Y(_09208_));
 sky130_vsdinv _39740_ (.A(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__nand2_4 _39741_ (.A(_03361_),
    .B(_05938_),
    .Y(_09210_));
 sky130_fd_sc_hd__o21ai_4 _39742_ (.A1(_03366_),
    .A2(_07618_),
    .B1(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__buf_1 _39743_ (.A(\pcpi_mul.rs1[24] ),
    .X(_09212_));
 sky130_fd_sc_hd__nand4_4 _39744_ (.A(_09088_),
    .B(_09212_),
    .C(_08047_),
    .D(_08043_),
    .Y(_09213_));
 sky130_fd_sc_hd__buf_1 _39745_ (.A(\pcpi_mul.rs1[25] ),
    .X(_09214_));
 sky130_fd_sc_hd__nand2_4 _39746_ (.A(_09214_),
    .B(_05954_),
    .Y(_09215_));
 sky130_vsdinv _39747_ (.A(_09215_),
    .Y(_09216_));
 sky130_fd_sc_hd__a21oi_4 _39748_ (.A1(_09211_),
    .A2(_09213_),
    .B1(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__nand3_4 _39749_ (.A(_09211_),
    .B(_09213_),
    .C(_09216_),
    .Y(_09218_));
 sky130_vsdinv _39750_ (.A(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__nor2_4 _39751_ (.A(_09217_),
    .B(_09219_),
    .Y(_09220_));
 sky130_vsdinv _39752_ (.A(_09207_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand3_4 _39753_ (.A(_09221_),
    .B(_09205_),
    .C(_09206_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand3_4 _39754_ (.A(_09209_),
    .B(_09220_),
    .C(_09222_),
    .Y(_09223_));
 sky130_vsdinv _39755_ (.A(_09222_),
    .Y(_09224_));
 sky130_vsdinv _39756_ (.A(_09220_),
    .Y(_09225_));
 sky130_fd_sc_hd__o21ai_4 _39757_ (.A1(_09208_),
    .A2(_09224_),
    .B1(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__nand3_4 _39758_ (.A(_09197_),
    .B(_09223_),
    .C(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__nand2_4 _39759_ (.A(_09226_),
    .B(_09223_),
    .Y(_09228_));
 sky130_fd_sc_hd__nand2_4 _39760_ (.A(_09228_),
    .B(_09196_),
    .Y(_09229_));
 sky130_fd_sc_hd__a21boi_4 _39761_ (.A1(_09085_),
    .A2(_09092_),
    .B1_N(_09089_),
    .Y(_09230_));
 sky130_vsdinv _39762_ (.A(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__a21oi_4 _39763_ (.A1(_09227_),
    .A2(_09229_),
    .B1(_09231_),
    .Y(_09232_));
 sky130_vsdinv _39764_ (.A(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__nand3_4 _39765_ (.A(_09227_),
    .B(_09229_),
    .C(_09231_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_4 _39766_ (.A(_09233_),
    .B(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand2_4 _39767_ (.A(_09194_),
    .B(_09235_),
    .Y(_09236_));
 sky130_fd_sc_hd__nand4_4 _39768_ (.A(_09234_),
    .B(_09191_),
    .C(_09233_),
    .D(_09193_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_4 _39769_ (.A(_09236_),
    .B(_09237_),
    .Y(_09238_));
 sky130_vsdinv _39770_ (.A(_08985_),
    .Y(_09239_));
 sky130_fd_sc_hd__a21oi_4 _39771_ (.A1(_08983_),
    .A2(_08987_),
    .B1(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__nand2_4 _39772_ (.A(_09238_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__a21o_4 _39773_ (.A1(_08983_),
    .A2(_08987_),
    .B1(_09239_),
    .X(_09242_));
 sky130_fd_sc_hd__nand3_4 _39774_ (.A(_09242_),
    .B(_09237_),
    .C(_09236_),
    .Y(_09243_));
 sky130_fd_sc_hd__nand2_4 _39775_ (.A(_09109_),
    .B(_09068_),
    .Y(_09244_));
 sky130_fd_sc_hd__nand3_4 _39776_ (.A(_09241_),
    .B(_09243_),
    .C(_09244_),
    .Y(_09245_));
 sky130_vsdinv _39777_ (.A(_09006_),
    .Y(_09246_));
 sky130_fd_sc_hd__a21boi_4 _39778_ (.A1(_09010_),
    .A2(_09246_),
    .B1_N(_09011_),
    .Y(_09247_));
 sky130_vsdinv _39779_ (.A(_09247_),
    .Y(_09248_));
 sky130_fd_sc_hd__nand2_4 _39780_ (.A(_08928_),
    .B(_07709_),
    .Y(_09249_));
 sky130_fd_sc_hd__nand2_4 _39781_ (.A(_07464_),
    .B(_08571_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand2_4 _39782_ (.A(_09249_),
    .B(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__nand4_4 _39783_ (.A(_06342_),
    .B(_03290_),
    .C(_08795_),
    .D(_03540_),
    .Y(_09252_));
 sky130_fd_sc_hd__nand2_4 _39784_ (.A(_06566_),
    .B(_03529_),
    .Y(_09253_));
 sky130_vsdinv _39785_ (.A(_09253_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand3_4 _39786_ (.A(_09251_),
    .B(_09252_),
    .C(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__nand2_4 _39787_ (.A(_09251_),
    .B(_09252_),
    .Y(_09256_));
 sky130_fd_sc_hd__nand2_4 _39788_ (.A(_09256_),
    .B(_09253_),
    .Y(_09257_));
 sky130_fd_sc_hd__nand3_4 _39789_ (.A(_09248_),
    .B(_09255_),
    .C(_09257_),
    .Y(_09258_));
 sky130_fd_sc_hd__nand2_4 _39790_ (.A(_09257_),
    .B(_09255_),
    .Y(_09259_));
 sky130_fd_sc_hd__nand2_4 _39791_ (.A(_09259_),
    .B(_09247_),
    .Y(_09260_));
 sky130_fd_sc_hd__nand2_4 _39792_ (.A(_09258_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__a21boi_4 _39793_ (.A1(_08930_),
    .A2(_08933_),
    .B1_N(_08931_),
    .Y(_09262_));
 sky130_fd_sc_hd__nand2_4 _39794_ (.A(_09261_),
    .B(_09262_),
    .Y(_09263_));
 sky130_vsdinv _39795_ (.A(_09262_),
    .Y(_09264_));
 sky130_fd_sc_hd__nand3_4 _39796_ (.A(_09258_),
    .B(_09260_),
    .C(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__nand2_4 _39797_ (.A(_09263_),
    .B(_09265_),
    .Y(_09266_));
 sky130_fd_sc_hd__a21boi_4 _39798_ (.A1(_08939_),
    .A2(_08943_),
    .B1_N(_08937_),
    .Y(_09267_));
 sky130_fd_sc_hd__nand2_4 _39799_ (.A(_09266_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__nand2_4 _39800_ (.A(_08944_),
    .B(_08937_),
    .Y(_09269_));
 sky130_fd_sc_hd__nand3_4 _39801_ (.A(_09269_),
    .B(_09265_),
    .C(_09263_),
    .Y(_09270_));
 sky130_fd_sc_hd__nand2_4 _39802_ (.A(_09268_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__nand2_4 _39803_ (.A(_03297_),
    .B(_07053_),
    .Y(_09272_));
 sky130_fd_sc_hd__nand2_4 _39804_ (.A(_06710_),
    .B(_07049_),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2_4 _39805_ (.A(_09272_),
    .B(_09273_),
    .Y(_09274_));
 sky130_fd_sc_hd__nand4_4 _39806_ (.A(_06842_),
    .B(_06710_),
    .C(_07355_),
    .D(_03524_),
    .Y(_09275_));
 sky130_fd_sc_hd__nand2_4 _39807_ (.A(_09274_),
    .B(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__nand2_4 _39808_ (.A(_03309_),
    .B(_07043_),
    .Y(_09277_));
 sky130_fd_sc_hd__nand2_4 _39809_ (.A(_09276_),
    .B(_09277_),
    .Y(_09278_));
 sky130_vsdinv _39810_ (.A(_09277_),
    .Y(_09279_));
 sky130_fd_sc_hd__nand3_4 _39811_ (.A(_09274_),
    .B(_09275_),
    .C(_09279_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_4 _39812_ (.A(_08961_),
    .B(_08956_),
    .Y(_09281_));
 sky130_fd_sc_hd__a21oi_4 _39813_ (.A1(_09278_),
    .A2(_09280_),
    .B1(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__nand3_4 _39814_ (.A(_09281_),
    .B(_09280_),
    .C(_09278_),
    .Y(_09283_));
 sky130_vsdinv _39815_ (.A(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__nand2_4 _39816_ (.A(_03324_),
    .B(_06750_),
    .Y(_09285_));
 sky130_vsdinv _39817_ (.A(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__nand2_4 _39818_ (.A(_07421_),
    .B(_06747_),
    .Y(_09287_));
 sky130_fd_sc_hd__nand2_4 _39819_ (.A(_07438_),
    .B(_03500_),
    .Y(_09288_));
 sky130_fd_sc_hd__nand2_4 _39820_ (.A(_09287_),
    .B(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nand4_4 _39821_ (.A(_07421_),
    .B(_07438_),
    .C(_03500_),
    .D(_06747_),
    .Y(_09290_));
 sky130_fd_sc_hd__nand2_4 _39822_ (.A(_09289_),
    .B(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__xor2_4 _39823_ (.A(_09286_),
    .B(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__o21ai_4 _39824_ (.A1(_09282_),
    .A2(_09284_),
    .B1(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__a21o_4 _39825_ (.A1(_09278_),
    .A2(_09280_),
    .B1(_09281_),
    .X(_09294_));
 sky130_fd_sc_hd__xor2_4 _39826_ (.A(_09285_),
    .B(_09291_),
    .X(_09295_));
 sky130_fd_sc_hd__nand3_4 _39827_ (.A(_09294_),
    .B(_09295_),
    .C(_09283_),
    .Y(_09296_));
 sky130_fd_sc_hd__and2_4 _39828_ (.A(_09293_),
    .B(_09296_),
    .X(_09297_));
 sky130_vsdinv _39829_ (.A(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__nand2_4 _39830_ (.A(_09271_),
    .B(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__nand3_4 _39831_ (.A(_09268_),
    .B(_09297_),
    .C(_09270_),
    .Y(_09300_));
 sky130_fd_sc_hd__nand2_4 _39832_ (.A(_09299_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__nand2_4 _39833_ (.A(_09301_),
    .B(_09018_),
    .Y(_09302_));
 sky130_vsdinv _39834_ (.A(_09018_),
    .Y(_09303_));
 sky130_fd_sc_hd__nand3_4 _39835_ (.A(_09299_),
    .B(_09300_),
    .C(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__nand2_4 _39836_ (.A(_09302_),
    .B(_09304_),
    .Y(_09305_));
 sky130_fd_sc_hd__o21a_4 _39837_ (.A1(_08977_),
    .A2(_08950_),
    .B1(_08949_),
    .X(_09306_));
 sky130_fd_sc_hd__nand2_4 _39838_ (.A(_09305_),
    .B(_09306_),
    .Y(_09307_));
 sky130_vsdinv _39839_ (.A(_09306_),
    .Y(_09308_));
 sky130_fd_sc_hd__nand3_4 _39840_ (.A(_09308_),
    .B(_09302_),
    .C(_09304_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand2_4 _39841_ (.A(_09307_),
    .B(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__a21boi_4 _39842_ (.A1(_09003_),
    .A2(_09013_),
    .B1_N(_09005_),
    .Y(_09311_));
 sky130_vsdinv _39843_ (.A(_09311_),
    .Y(_09312_));
 sky130_fd_sc_hd__buf_1 _39844_ (.A(_03574_),
    .X(_09313_));
 sky130_fd_sc_hd__nand2_4 _39845_ (.A(_06126_),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__nand2_4 _39846_ (.A(_03256_),
    .B(_08995_),
    .Y(_09315_));
 sky130_fd_sc_hd__nand2_4 _39847_ (.A(_09314_),
    .B(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__nand4_4 _39848_ (.A(_05935_),
    .B(_06007_),
    .C(_08630_),
    .D(_09313_),
    .Y(_09317_));
 sky130_fd_sc_hd__nand2_4 _39849_ (.A(_06141_),
    .B(_08634_),
    .Y(_09318_));
 sky130_vsdinv _39850_ (.A(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__a21o_4 _39851_ (.A1(_09316_),
    .A2(_09317_),
    .B1(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__nand3_4 _39852_ (.A(_09316_),
    .B(_09317_),
    .C(_09319_),
    .Y(_09321_));
 sky130_fd_sc_hd__nand2_4 _39853_ (.A(_09320_),
    .B(_09321_),
    .Y(_09322_));
 sky130_fd_sc_hd__a21boi_4 _39854_ (.A1(_08994_),
    .A2(_08998_),
    .B1_N(_08996_),
    .Y(_09323_));
 sky130_fd_sc_hd__nand2_4 _39855_ (.A(_09322_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__nand2_4 _39856_ (.A(_06544_),
    .B(_08640_),
    .Y(_09325_));
 sky130_fd_sc_hd__nand2_4 _39857_ (.A(_07525_),
    .B(_08875_),
    .Y(_09326_));
 sky130_fd_sc_hd__nand2_4 _39858_ (.A(_06937_),
    .B(_08190_),
    .Y(_09327_));
 sky130_fd_sc_hd__nand2_4 _39859_ (.A(_09326_),
    .B(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__nand4_4 _39860_ (.A(_06075_),
    .B(_06937_),
    .C(_08643_),
    .D(_08197_),
    .Y(_09329_));
 sky130_fd_sc_hd__nand2_4 _39861_ (.A(_09328_),
    .B(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__xor2_4 _39862_ (.A(_09325_),
    .B(_09330_),
    .X(_09331_));
 sky130_vsdinv _39863_ (.A(_09323_),
    .Y(_09332_));
 sky130_fd_sc_hd__nand3_4 _39864_ (.A(_09332_),
    .B(_09321_),
    .C(_09320_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand3_4 _39865_ (.A(_09324_),
    .B(_09331_),
    .C(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_4 _39866_ (.A(_09324_),
    .B(_09333_),
    .Y(_09335_));
 sky130_vsdinv _39867_ (.A(_09331_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand2_4 _39868_ (.A(_09335_),
    .B(_09336_),
    .Y(_09337_));
 sky130_fd_sc_hd__nand3_4 _39869_ (.A(_09312_),
    .B(_09334_),
    .C(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__nand2_4 _39870_ (.A(_09337_),
    .B(_09334_),
    .Y(_09339_));
 sky130_fd_sc_hd__nand2_4 _39871_ (.A(_09339_),
    .B(_09311_),
    .Y(_09340_));
 sky130_fd_sc_hd__nand2_4 _39872_ (.A(_09338_),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__buf_1 _39873_ (.A(\pcpi_mul.rs2[25] ),
    .X(_09342_));
 sky130_fd_sc_hd__buf_1 _39874_ (.A(_09342_),
    .X(_09343_));
 sky130_fd_sc_hd__buf_1 _39875_ (.A(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__nand2_4 _39876_ (.A(_05584_),
    .B(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__buf_1 _39877_ (.A(\pcpi_mul.rs2[24] ),
    .X(_09346_));
 sky130_fd_sc_hd__buf_1 _39878_ (.A(_09346_),
    .X(_09347_));
 sky130_fd_sc_hd__nand2_4 _39879_ (.A(_06746_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__nor2_4 _39880_ (.A(_09345_),
    .B(_09348_),
    .Y(_09349_));
 sky130_vsdinv _39881_ (.A(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__nand2_4 _39882_ (.A(_09345_),
    .B(_09348_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand2_4 _39883_ (.A(_09350_),
    .B(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_4 _39884_ (.A(_09341_),
    .B(_09352_),
    .Y(_09353_));
 sky130_vsdinv _39885_ (.A(_09352_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand3_4 _39886_ (.A(_09338_),
    .B(_09340_),
    .C(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__nand2_4 _39887_ (.A(_09353_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__nand2_4 _39888_ (.A(_09356_),
    .B(_09022_),
    .Y(_09357_));
 sky130_fd_sc_hd__nand3_4 _39889_ (.A(_09023_),
    .B(_09353_),
    .C(_09355_),
    .Y(_09358_));
 sky130_fd_sc_hd__and2_4 _39890_ (.A(_09357_),
    .B(_09358_),
    .X(_09359_));
 sky130_vsdinv _39891_ (.A(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__nand2_4 _39892_ (.A(_09310_),
    .B(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__nand3_4 _39893_ (.A(_09359_),
    .B(_09307_),
    .C(_09309_),
    .Y(_09362_));
 sky130_fd_sc_hd__nand2_4 _39894_ (.A(_09361_),
    .B(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__nand2_4 _39895_ (.A(_09363_),
    .B(_09026_),
    .Y(_09364_));
 sky130_fd_sc_hd__nand2_4 _39896_ (.A(_09241_),
    .B(_09243_),
    .Y(_09365_));
 sky130_vsdinv _39897_ (.A(_09244_),
    .Y(_09366_));
 sky130_fd_sc_hd__nand2_4 _39898_ (.A(_09365_),
    .B(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand3_4 _39899_ (.A(_09361_),
    .B(_09027_),
    .C(_09362_),
    .Y(_09368_));
 sky130_fd_sc_hd__nand4_4 _39900_ (.A(_09245_),
    .B(_09364_),
    .C(_09367_),
    .D(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__nand2_4 _39901_ (.A(_09364_),
    .B(_09368_),
    .Y(_09370_));
 sky130_fd_sc_hd__nand2_4 _39902_ (.A(_09367_),
    .B(_09245_),
    .Y(_09371_));
 sky130_fd_sc_hd__nand2_4 _39903_ (.A(_09370_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__nand3_4 _39904_ (.A(_09158_),
    .B(_09369_),
    .C(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand2_4 _39905_ (.A(_09372_),
    .B(_09369_),
    .Y(_09374_));
 sky130_fd_sc_hd__nand3_4 _39906_ (.A(_09374_),
    .B(_09031_),
    .C(_09122_),
    .Y(_09375_));
 sky130_fd_sc_hd__nand2_4 _39907_ (.A(_09373_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__a21boi_4 _39908_ (.A1(_09105_),
    .A2(_09101_),
    .B1_N(_09100_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand2_4 _39909_ (.A(_09119_),
    .B(_09114_),
    .Y(_09378_));
 sky130_fd_sc_hd__xor2_4 _39910_ (.A(_09377_),
    .B(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__nand2_4 _39911_ (.A(_09376_),
    .B(_09379_),
    .Y(_09380_));
 sky130_vsdinv _39912_ (.A(_09379_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand3_4 _39913_ (.A(_09373_),
    .B(_09375_),
    .C(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__nand2_4 _39914_ (.A(_09380_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__a21boi_4 _39915_ (.A1(_09124_),
    .A2(_09132_),
    .B1_N(_09126_),
    .Y(_09384_));
 sky130_fd_sc_hd__nand2_4 _39916_ (.A(_09383_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__nand2_4 _39917_ (.A(_09133_),
    .B(_09126_),
    .Y(_09386_));
 sky130_fd_sc_hd__nand3_4 _39918_ (.A(_09386_),
    .B(_09382_),
    .C(_09380_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand2_4 _39919_ (.A(_09385_),
    .B(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__a21oi_4 _39920_ (.A1(_08789_),
    .A2(_08784_),
    .B1(_09128_),
    .Y(_09389_));
 sky130_vsdinv _39921_ (.A(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__nand2_4 _39922_ (.A(_09388_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__nand3_4 _39923_ (.A(_09385_),
    .B(_09387_),
    .C(_09389_),
    .Y(_09392_));
 sky130_fd_sc_hd__a21oi_4 _39924_ (.A1(_09131_),
    .A2(_09133_),
    .B1(_09137_),
    .Y(_09393_));
 sky130_fd_sc_hd__o21ai_4 _39925_ (.A1(_09141_),
    .A2(_09393_),
    .B1(_09138_),
    .Y(_09394_));
 sky130_fd_sc_hd__a21oi_4 _39926_ (.A1(_09391_),
    .A2(_09392_),
    .B1(_09394_),
    .Y(_09395_));
 sky130_fd_sc_hd__nand3_4 _39927_ (.A(_09394_),
    .B(_09391_),
    .C(_09392_),
    .Y(_09396_));
 sky130_vsdinv _39928_ (.A(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__nor2_4 _39929_ (.A(_09395_),
    .B(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__o21ai_4 _39930_ (.A1(_09146_),
    .A2(_09157_),
    .B1(_09147_),
    .Y(_09399_));
 sky130_fd_sc_hd__xor2_4 _39931_ (.A(_09398_),
    .B(_09399_),
    .X(_01430_));
 sky130_fd_sc_hd__o21a_4 _39932_ (.A1(_09371_),
    .A2(_09370_),
    .B1(_09368_),
    .X(_09400_));
 sky130_fd_sc_hd__nand2_4 _39933_ (.A(_09362_),
    .B(_09358_),
    .Y(_09401_));
 sky130_vsdinv _39934_ (.A(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__nand2_4 _39935_ (.A(_06450_),
    .B(_07921_),
    .Y(_09403_));
 sky130_fd_sc_hd__nand2_4 _39936_ (.A(_03293_),
    .B(_07712_),
    .Y(_09404_));
 sky130_fd_sc_hd__nand2_4 _39937_ (.A(_09403_),
    .B(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__nand4_4 _39938_ (.A(_07464_),
    .B(_06566_),
    .C(_08127_),
    .D(_08124_),
    .Y(_09406_));
 sky130_fd_sc_hd__nand2_4 _39939_ (.A(_09405_),
    .B(_09406_),
    .Y(_09407_));
 sky130_fd_sc_hd__nand2_4 _39940_ (.A(_08606_),
    .B(_07561_),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_4 _39941_ (.A(_09407_),
    .B(_09408_),
    .Y(_09409_));
 sky130_vsdinv _39942_ (.A(_09408_),
    .Y(_09410_));
 sky130_fd_sc_hd__nand3_4 _39943_ (.A(_09405_),
    .B(_09406_),
    .C(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__nand2_4 _39944_ (.A(_09409_),
    .B(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__maj3_4 _39945_ (.A(_09325_),
    .B(_09326_),
    .C(_09327_),
    .X(_09413_));
 sky130_fd_sc_hd__nand2_4 _39946_ (.A(_09412_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__buf_1 _39947_ (.A(_03556_),
    .X(_09415_));
 sky130_fd_sc_hd__buf_1 _39948_ (.A(_09008_),
    .X(_09416_));
 sky130_fd_sc_hd__a22oi_4 _39949_ (.A1(_08565_),
    .A2(_09415_),
    .B1(_07346_),
    .B2(_09416_),
    .Y(_09417_));
 sky130_fd_sc_hd__o21ai_4 _39950_ (.A1(_09325_),
    .A2(_09417_),
    .B1(_09329_),
    .Y(_09418_));
 sky130_fd_sc_hd__nand3_4 _39951_ (.A(_09418_),
    .B(_09411_),
    .C(_09409_),
    .Y(_09419_));
 sky130_fd_sc_hd__nand2_4 _39952_ (.A(_09414_),
    .B(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__a21boi_4 _39953_ (.A1(_09251_),
    .A2(_09254_),
    .B1_N(_09252_),
    .Y(_09421_));
 sky130_fd_sc_hd__nand2_4 _39954_ (.A(_09420_),
    .B(_09421_),
    .Y(_09422_));
 sky130_vsdinv _39955_ (.A(_09421_),
    .Y(_09423_));
 sky130_fd_sc_hd__nand3_4 _39956_ (.A(_09414_),
    .B(_09419_),
    .C(_09423_),
    .Y(_09424_));
 sky130_fd_sc_hd__nand2_4 _39957_ (.A(_09422_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__a21boi_4 _39958_ (.A1(_09260_),
    .A2(_09264_),
    .B1_N(_09258_),
    .Y(_09426_));
 sky130_fd_sc_hd__nand2_4 _39959_ (.A(_09425_),
    .B(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_4 _39960_ (.A(_09265_),
    .B(_09258_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand3_4 _39961_ (.A(_09428_),
    .B(_09424_),
    .C(_09422_),
    .Y(_09429_));
 sky130_fd_sc_hd__nand2_4 _39962_ (.A(_09280_),
    .B(_09275_),
    .Y(_09430_));
 sky130_vsdinv _39963_ (.A(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__nand2_4 _39964_ (.A(_03302_),
    .B(_03524_),
    .Y(_09432_));
 sky130_fd_sc_hd__nand2_4 _39965_ (.A(_07145_),
    .B(_07355_),
    .Y(_09433_));
 sky130_fd_sc_hd__nand2_4 _39966_ (.A(_09432_),
    .B(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__nand4_4 _39967_ (.A(_07818_),
    .B(_06998_),
    .C(_08953_),
    .D(_07733_),
    .Y(_09435_));
 sky130_fd_sc_hd__nand2_4 _39968_ (.A(_09434_),
    .B(_09435_),
    .Y(_09436_));
 sky130_fd_sc_hd__nand2_4 _39969_ (.A(_07297_),
    .B(_07043_),
    .Y(_09437_));
 sky130_fd_sc_hd__nand2_4 _39970_ (.A(_09436_),
    .B(_09437_),
    .Y(_09438_));
 sky130_vsdinv _39971_ (.A(_09437_),
    .Y(_09439_));
 sky130_fd_sc_hd__nand3_4 _39972_ (.A(_09434_),
    .B(_09435_),
    .C(_09439_),
    .Y(_09440_));
 sky130_fd_sc_hd__nand2_4 _39973_ (.A(_09438_),
    .B(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__nand2_4 _39974_ (.A(_09431_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__nand3_4 _39975_ (.A(_09430_),
    .B(_09440_),
    .C(_09438_),
    .Y(_09443_));
 sky130_fd_sc_hd__nand2_4 _39976_ (.A(_07443_),
    .B(_06750_),
    .Y(_09444_));
 sky130_fd_sc_hd__nand2_4 _39977_ (.A(_07301_),
    .B(_08162_),
    .Y(_09445_));
 sky130_fd_sc_hd__nand2_4 _39978_ (.A(_08289_),
    .B(_03500_),
    .Y(_09446_));
 sky130_fd_sc_hd__nand2_4 _39979_ (.A(_09445_),
    .B(_09446_),
    .Y(_09447_));
 sky130_fd_sc_hd__nand4_4 _39980_ (.A(_08966_),
    .B(_08294_),
    .C(_06505_),
    .D(_06636_),
    .Y(_09448_));
 sky130_fd_sc_hd__nand2_4 _39981_ (.A(_09447_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__xor2_4 _39982_ (.A(_09444_),
    .B(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__a21oi_4 _39983_ (.A1(_09442_),
    .A2(_09443_),
    .B1(_09450_),
    .Y(_09451_));
 sky130_fd_sc_hd__nand3_4 _39984_ (.A(_09450_),
    .B(_09442_),
    .C(_09443_),
    .Y(_09452_));
 sky130_vsdinv _39985_ (.A(_09452_),
    .Y(_09453_));
 sky130_fd_sc_hd__nor2_4 _39986_ (.A(_09451_),
    .B(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__a21o_4 _39987_ (.A1(_09427_),
    .A2(_09429_),
    .B1(_09454_),
    .X(_09455_));
 sky130_fd_sc_hd__nand3_4 _39988_ (.A(_09427_),
    .B(_09429_),
    .C(_09454_),
    .Y(_09456_));
 sky130_fd_sc_hd__nand2_4 _39989_ (.A(_09455_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__nand2_4 _39990_ (.A(_09457_),
    .B(_09338_),
    .Y(_09458_));
 sky130_vsdinv _39991_ (.A(_09338_),
    .Y(_09459_));
 sky130_fd_sc_hd__nand3_4 _39992_ (.A(_09455_),
    .B(_09459_),
    .C(_09456_),
    .Y(_09460_));
 sky130_fd_sc_hd__nand2_4 _39993_ (.A(_09458_),
    .B(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__a21boi_4 _39994_ (.A1(_09268_),
    .A2(_09297_),
    .B1_N(_09270_),
    .Y(_09462_));
 sky130_fd_sc_hd__nand2_4 _39995_ (.A(_09461_),
    .B(_09462_),
    .Y(_09463_));
 sky130_vsdinv _39996_ (.A(_09462_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand3_4 _39997_ (.A(_09458_),
    .B(_09464_),
    .C(_09460_),
    .Y(_09465_));
 sky130_fd_sc_hd__nand2_4 _39998_ (.A(_09463_),
    .B(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__buf_1 _39999_ (.A(\pcpi_mul.rs2[23] ),
    .X(_09467_));
 sky130_fd_sc_hd__nand2_4 _40000_ (.A(_06383_),
    .B(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand2_4 _40001_ (.A(_07364_),
    .B(_03568_),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_4 _40002_ (.A(_09468_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__nand4_4 _40003_ (.A(_03256_),
    .B(_07364_),
    .C(_08995_),
    .D(_08862_),
    .Y(_09471_));
 sky130_fd_sc_hd__nand2_4 _40004_ (.A(_06018_),
    .B(_03562_),
    .Y(_09472_));
 sky130_vsdinv _40005_ (.A(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__a21o_4 _40006_ (.A1(_09470_),
    .A2(_09471_),
    .B1(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__nand3_4 _40007_ (.A(_09470_),
    .B(_09471_),
    .C(_09473_),
    .Y(_09475_));
 sky130_fd_sc_hd__nand2_4 _40008_ (.A(_09474_),
    .B(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__a21boi_4 _40009_ (.A1(_09316_),
    .A2(_09319_),
    .B1_N(_09317_),
    .Y(_09477_));
 sky130_fd_sc_hd__nand2_4 _40010_ (.A(_09476_),
    .B(_09477_),
    .Y(_09478_));
 sky130_vsdinv _40011_ (.A(_09477_),
    .Y(_09479_));
 sky130_fd_sc_hd__nand3_4 _40012_ (.A(_09479_),
    .B(_09475_),
    .C(_09474_),
    .Y(_09480_));
 sky130_fd_sc_hd__nand2_4 _40013_ (.A(_09478_),
    .B(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__nand2_4 _40014_ (.A(_08928_),
    .B(_08873_),
    .Y(_09482_));
 sky130_fd_sc_hd__nand2_4 _40015_ (.A(_06169_),
    .B(_08875_),
    .Y(_09483_));
 sky130_fd_sc_hd__nand2_4 _40016_ (.A(_06544_),
    .B(_08643_),
    .Y(_09484_));
 sky130_fd_sc_hd__nand2_4 _40017_ (.A(_09483_),
    .B(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__buf_1 _40018_ (.A(_03556_),
    .X(_09486_));
 sky130_fd_sc_hd__nand4_4 _40019_ (.A(_06244_),
    .B(_06251_),
    .C(_07976_),
    .D(_09486_),
    .Y(_09487_));
 sky130_fd_sc_hd__nand2_4 _40020_ (.A(_09485_),
    .B(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__xor2_4 _40021_ (.A(_09482_),
    .B(_09488_),
    .X(_09489_));
 sky130_vsdinv _40022_ (.A(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__nand2_4 _40023_ (.A(_09481_),
    .B(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__nand3_4 _40024_ (.A(_09478_),
    .B(_09489_),
    .C(_09480_),
    .Y(_09492_));
 sky130_fd_sc_hd__nand2_4 _40025_ (.A(_09491_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__a21boi_4 _40026_ (.A1(_09324_),
    .A2(_09331_),
    .B1_N(_09333_),
    .Y(_09494_));
 sky130_fd_sc_hd__nand2_4 _40027_ (.A(_09493_),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__nand2_4 _40028_ (.A(_09334_),
    .B(_09333_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand3_4 _40029_ (.A(_09496_),
    .B(_09492_),
    .C(_09491_),
    .Y(_09497_));
 sky130_fd_sc_hd__nand2_4 _40030_ (.A(_09495_),
    .B(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_4 _40031_ (.A(_08991_),
    .B(_09342_),
    .Y(_09499_));
 sky130_fd_sc_hd__buf_1 _40032_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09500_));
 sky130_fd_sc_hd__nand2_4 _40033_ (.A(_08859_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__nand2_4 _40034_ (.A(_09499_),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__nand4_4 _40035_ (.A(_08859_),
    .B(_08991_),
    .C(_03586_),
    .D(_09500_),
    .Y(_09503_));
 sky130_fd_sc_hd__nand2_4 _40036_ (.A(_06054_),
    .B(_03580_),
    .Y(_09504_));
 sky130_vsdinv _40037_ (.A(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__a21o_4 _40038_ (.A1(_09502_),
    .A2(_09503_),
    .B1(_09505_),
    .X(_09506_));
 sky130_fd_sc_hd__nand3_4 _40039_ (.A(_09502_),
    .B(_09503_),
    .C(_09505_),
    .Y(_09507_));
 sky130_fd_sc_hd__and2_4 _40040_ (.A(_09506_),
    .B(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__xor2_4 _40041_ (.A(_09349_),
    .B(_09508_),
    .X(_09509_));
 sky130_vsdinv _40042_ (.A(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__nand2_4 _40043_ (.A(_09498_),
    .B(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand3_4 _40044_ (.A(_09495_),
    .B(_09497_),
    .C(_09509_),
    .Y(_09512_));
 sky130_fd_sc_hd__nand2_4 _40045_ (.A(_09511_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__nand2_4 _40046_ (.A(_09513_),
    .B(_09355_),
    .Y(_09514_));
 sky130_vsdinv _40047_ (.A(_09355_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand3_4 _40048_ (.A(_09515_),
    .B(_09511_),
    .C(_09512_),
    .Y(_09516_));
 sky130_fd_sc_hd__and2_4 _40049_ (.A(_09514_),
    .B(_09516_),
    .X(_09517_));
 sky130_vsdinv _40050_ (.A(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__nand2_4 _40051_ (.A(_09466_),
    .B(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__nand3_4 _40052_ (.A(_09463_),
    .B(_09517_),
    .C(_09465_),
    .Y(_09520_));
 sky130_fd_sc_hd__nand2_4 _40053_ (.A(_09519_),
    .B(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand2_4 _40054_ (.A(_09402_),
    .B(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand3_4 _40055_ (.A(_09401_),
    .B(_09520_),
    .C(_09519_),
    .Y(_09523_));
 sky130_fd_sc_hd__nand2_4 _40056_ (.A(_09522_),
    .B(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__nand2_4 _40057_ (.A(_03335_),
    .B(_03490_),
    .Y(_09525_));
 sky130_fd_sc_hd__nand2_4 _40058_ (.A(_08045_),
    .B(_06375_),
    .Y(_09526_));
 sky130_fd_sc_hd__nand2_4 _40059_ (.A(_09525_),
    .B(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__nand4_4 _40060_ (.A(_08050_),
    .B(_07877_),
    .C(_07095_),
    .D(_08081_),
    .Y(_09528_));
 sky130_fd_sc_hd__nand2_4 _40061_ (.A(_09527_),
    .B(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__nand2_4 _40062_ (.A(_03346_),
    .B(_03475_),
    .Y(_09530_));
 sky130_fd_sc_hd__nand2_4 _40063_ (.A(_09529_),
    .B(_09530_),
    .Y(_09531_));
 sky130_vsdinv _40064_ (.A(_09530_),
    .Y(_09532_));
 sky130_fd_sc_hd__nand3_4 _40065_ (.A(_09527_),
    .B(_09528_),
    .C(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__nand2_4 _40066_ (.A(_09531_),
    .B(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__a21boi_4 _40067_ (.A1(_09289_),
    .A2(_09286_),
    .B1_N(_09290_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand2_4 _40068_ (.A(_09534_),
    .B(_09535_),
    .Y(_09536_));
 sky130_vsdinv _40069_ (.A(_09290_),
    .Y(_09537_));
 sky130_fd_sc_hd__a21o_4 _40070_ (.A1(_09289_),
    .A2(_09286_),
    .B1(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__nand3_4 _40071_ (.A(_09538_),
    .B(_09533_),
    .C(_09531_),
    .Y(_09539_));
 sky130_fd_sc_hd__nand2_4 _40072_ (.A(_09536_),
    .B(_09539_),
    .Y(_09540_));
 sky130_fd_sc_hd__a21boi_4 _40073_ (.A1(_09163_),
    .A2(_09166_),
    .B1_N(_09164_),
    .Y(_09541_));
 sky130_fd_sc_hd__nand2_4 _40074_ (.A(_09540_),
    .B(_09541_),
    .Y(_09542_));
 sky130_vsdinv _40075_ (.A(_09541_),
    .Y(_09543_));
 sky130_fd_sc_hd__nand3_4 _40076_ (.A(_09536_),
    .B(_09539_),
    .C(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nand2_4 _40077_ (.A(_09542_),
    .B(_09544_),
    .Y(_09545_));
 sky130_fd_sc_hd__a21oi_4 _40078_ (.A1(_09294_),
    .A2(_09295_),
    .B1(_09284_),
    .Y(_09546_));
 sky130_fd_sc_hd__nand2_4 _40079_ (.A(_09545_),
    .B(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__o21ai_4 _40080_ (.A1(_09282_),
    .A2(_09292_),
    .B1(_09283_),
    .Y(_09548_));
 sky130_fd_sc_hd__nand3_4 _40081_ (.A(_09548_),
    .B(_09542_),
    .C(_09544_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand2_4 _40082_ (.A(_09547_),
    .B(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__a21boi_4 _40083_ (.A1(_09173_),
    .A2(_09177_),
    .B1_N(_09170_),
    .Y(_09551_));
 sky130_fd_sc_hd__nand2_4 _40084_ (.A(_09550_),
    .B(_09551_),
    .Y(_09552_));
 sky130_vsdinv _40085_ (.A(_09551_),
    .Y(_09553_));
 sky130_fd_sc_hd__nand3_4 _40086_ (.A(_09547_),
    .B(_09553_),
    .C(_09549_),
    .Y(_09554_));
 sky130_fd_sc_hd__nand2_4 _40087_ (.A(_09552_),
    .B(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__a21boi_4 _40088_ (.A1(_09181_),
    .A2(_09187_),
    .B1_N(_09183_),
    .Y(_09556_));
 sky130_fd_sc_hd__nand2_4 _40089_ (.A(_09555_),
    .B(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand2_4 _40090_ (.A(_09188_),
    .B(_09183_),
    .Y(_09558_));
 sky130_fd_sc_hd__nand3_4 _40091_ (.A(_09558_),
    .B(_09552_),
    .C(_09554_),
    .Y(_09559_));
 sky130_fd_sc_hd__nand2_4 _40092_ (.A(_09557_),
    .B(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__nand2_4 _40093_ (.A(_08527_),
    .B(_08505_),
    .Y(_09561_));
 sky130_fd_sc_hd__nand2_4 _40094_ (.A(_09202_),
    .B(_08507_),
    .Y(_09562_));
 sky130_fd_sc_hd__nand2_4 _40095_ (.A(_09561_),
    .B(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__nand4_4 _40096_ (.A(_08527_),
    .B(_03357_),
    .C(_07131_),
    .D(_08505_),
    .Y(_09564_));
 sky130_fd_sc_hd__buf_1 _40097_ (.A(\pcpi_mul.rs1[23] ),
    .X(_09565_));
 sky130_fd_sc_hd__nand2_4 _40098_ (.A(_09565_),
    .B(_05995_),
    .Y(_09566_));
 sky130_vsdinv _40099_ (.A(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand3_4 _40100_ (.A(_09563_),
    .B(_09564_),
    .C(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__a21o_4 _40101_ (.A1(_09563_),
    .A2(_09564_),
    .B1(_09567_),
    .X(_09569_));
 sky130_fd_sc_hd__a21boi_4 _40102_ (.A1(_09200_),
    .A2(_09204_),
    .B1_N(_09201_),
    .Y(_09570_));
 sky130_vsdinv _40103_ (.A(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__a21o_4 _40104_ (.A1(_09568_),
    .A2(_09569_),
    .B1(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__nand3_4 _40105_ (.A(_09571_),
    .B(_09568_),
    .C(_09569_),
    .Y(_09573_));
 sky130_fd_sc_hd__buf_1 _40106_ (.A(_03365_),
    .X(_09574_));
 sky130_fd_sc_hd__nand2_4 _40107_ (.A(_09574_),
    .B(_05939_),
    .Y(_09575_));
 sky130_fd_sc_hd__o21ai_4 _40108_ (.A1(_03376_),
    .A2(_07144_),
    .B1(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__buf_1 _40109_ (.A(_09090_),
    .X(_09577_));
 sky130_fd_sc_hd__buf_1 _40110_ (.A(_09214_),
    .X(_09578_));
 sky130_fd_sc_hd__nand4_4 _40111_ (.A(_09577_),
    .B(_09578_),
    .C(_08310_),
    .D(_08311_),
    .Y(_09579_));
 sky130_fd_sc_hd__buf_1 _40112_ (.A(_03379_),
    .X(_09580_));
 sky130_fd_sc_hd__nand2_4 _40113_ (.A(_09580_),
    .B(_05955_),
    .Y(_09581_));
 sky130_vsdinv _40114_ (.A(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__a21oi_4 _40115_ (.A1(_09576_),
    .A2(_09579_),
    .B1(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__nand3_4 _40116_ (.A(_09576_),
    .B(_09579_),
    .C(_09582_),
    .Y(_09584_));
 sky130_vsdinv _40117_ (.A(_09584_),
    .Y(_09585_));
 sky130_fd_sc_hd__nor2_4 _40118_ (.A(_09583_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__a21o_4 _40119_ (.A1(_09572_),
    .A2(_09573_),
    .B1(_09586_),
    .X(_09587_));
 sky130_fd_sc_hd__nand3_4 _40120_ (.A(_09572_),
    .B(_09586_),
    .C(_09573_),
    .Y(_09588_));
 sky130_fd_sc_hd__nand2_4 _40121_ (.A(_09587_),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__o21ai_4 _40122_ (.A1(_09208_),
    .A2(_09225_),
    .B1(_09222_),
    .Y(_09590_));
 sky130_vsdinv _40123_ (.A(_09590_),
    .Y(_09591_));
 sky130_fd_sc_hd__nand2_4 _40124_ (.A(_09589_),
    .B(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__nand3_4 _40125_ (.A(_09587_),
    .B(_09590_),
    .C(_09588_),
    .Y(_09593_));
 sky130_fd_sc_hd__a21boi_4 _40126_ (.A1(_09211_),
    .A2(_09216_),
    .B1_N(_09213_),
    .Y(_09594_));
 sky130_vsdinv _40127_ (.A(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__a21oi_4 _40128_ (.A1(_09592_),
    .A2(_09593_),
    .B1(_09595_),
    .Y(_09596_));
 sky130_vsdinv _40129_ (.A(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__nand3_4 _40130_ (.A(_09592_),
    .B(_09595_),
    .C(_09593_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand2_4 _40131_ (.A(_09597_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__nand2_4 _40132_ (.A(_09560_),
    .B(_09599_),
    .Y(_09600_));
 sky130_vsdinv _40133_ (.A(_09598_),
    .Y(_09601_));
 sky130_fd_sc_hd__nor2_4 _40134_ (.A(_09596_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__nand3_4 _40135_ (.A(_09602_),
    .B(_09559_),
    .C(_09557_),
    .Y(_09603_));
 sky130_fd_sc_hd__nand2_4 _40136_ (.A(_09600_),
    .B(_09603_),
    .Y(_09604_));
 sky130_vsdinv _40137_ (.A(_09304_),
    .Y(_09605_));
 sky130_fd_sc_hd__a21oi_4 _40138_ (.A1(_09308_),
    .A2(_09302_),
    .B1(_09605_),
    .Y(_09606_));
 sky130_fd_sc_hd__nand2_4 _40139_ (.A(_09604_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__a21o_4 _40140_ (.A1(_09308_),
    .A2(_09302_),
    .B1(_09605_),
    .X(_09608_));
 sky130_fd_sc_hd__nand3_4 _40141_ (.A(_09608_),
    .B(_09600_),
    .C(_09603_),
    .Y(_09609_));
 sky130_fd_sc_hd__nand2_4 _40142_ (.A(_09607_),
    .B(_09609_),
    .Y(_09610_));
 sky130_fd_sc_hd__o21a_4 _40143_ (.A1(_09235_),
    .A2(_09194_),
    .B1(_09193_),
    .X(_09611_));
 sky130_fd_sc_hd__nand2_4 _40144_ (.A(_09610_),
    .B(_09611_),
    .Y(_09612_));
 sky130_vsdinv _40145_ (.A(_09611_),
    .Y(_09613_));
 sky130_fd_sc_hd__nand3_4 _40146_ (.A(_09613_),
    .B(_09607_),
    .C(_09609_),
    .Y(_09614_));
 sky130_fd_sc_hd__nand2_4 _40147_ (.A(_09612_),
    .B(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__nand2_4 _40148_ (.A(_09524_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__nand4_4 _40149_ (.A(_09614_),
    .B(_09522_),
    .C(_09612_),
    .D(_09523_),
    .Y(_09617_));
 sky130_fd_sc_hd__nand2_4 _40150_ (.A(_09616_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__nand2_4 _40151_ (.A(_09400_),
    .B(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__nand2_4 _40152_ (.A(_09369_),
    .B(_09368_),
    .Y(_09620_));
 sky130_fd_sc_hd__nand3_4 _40153_ (.A(_09620_),
    .B(_09617_),
    .C(_09616_),
    .Y(_09621_));
 sky130_fd_sc_hd__nand2_4 _40154_ (.A(_09619_),
    .B(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__a21boi_4 _40155_ (.A1(_09229_),
    .A2(_09231_),
    .B1_N(_09227_),
    .Y(_09623_));
 sky130_fd_sc_hd__nand2_4 _40156_ (.A(_09245_),
    .B(_09243_),
    .Y(_09624_));
 sky130_fd_sc_hd__xor2_4 _40157_ (.A(_09623_),
    .B(_09624_),
    .X(_09625_));
 sky130_fd_sc_hd__nand2_4 _40158_ (.A(_09622_),
    .B(_09625_),
    .Y(_09626_));
 sky130_vsdinv _40159_ (.A(_09625_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand3_4 _40160_ (.A(_09619_),
    .B(_09621_),
    .C(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__nand2_4 _40161_ (.A(_09626_),
    .B(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__a21boi_4 _40162_ (.A1(_09375_),
    .A2(_09381_),
    .B1_N(_09373_),
    .Y(_09630_));
 sky130_fd_sc_hd__nand2_4 _40163_ (.A(_09629_),
    .B(_09630_),
    .Y(_09631_));
 sky130_fd_sc_hd__nand2_4 _40164_ (.A(_09382_),
    .B(_09373_),
    .Y(_09632_));
 sky130_fd_sc_hd__nand3_4 _40165_ (.A(_09632_),
    .B(_09628_),
    .C(_09626_),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2_4 _40166_ (.A(_09631_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__a21oi_4 _40167_ (.A1(_09119_),
    .A2(_09114_),
    .B1(_09377_),
    .Y(_09635_));
 sky130_vsdinv _40168_ (.A(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__nand2_4 _40169_ (.A(_09634_),
    .B(_09636_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand3_4 _40170_ (.A(_09631_),
    .B(_09633_),
    .C(_09635_),
    .Y(_09638_));
 sky130_fd_sc_hd__nand2_4 _40171_ (.A(_09637_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__a21boi_4 _40172_ (.A1(_09385_),
    .A2(_09389_),
    .B1_N(_09387_),
    .Y(_09640_));
 sky130_fd_sc_hd__nand2_4 _40173_ (.A(_09639_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__nand2_4 _40174_ (.A(_09392_),
    .B(_09387_),
    .Y(_09642_));
 sky130_fd_sc_hd__nand3_4 _40175_ (.A(_09642_),
    .B(_09637_),
    .C(_09638_),
    .Y(_09643_));
 sky130_fd_sc_hd__and2_4 _40176_ (.A(_09641_),
    .B(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__buf_1 _40177_ (.A(_09644_),
    .X(_09645_));
 sky130_vsdinv _40178_ (.A(_09645_),
    .Y(_09646_));
 sky130_vsdinv _40179_ (.A(_09157_),
    .Y(_09647_));
 sky130_fd_sc_hd__and2_4 _40180_ (.A(_09398_),
    .B(_09149_),
    .X(_09648_));
 sky130_fd_sc_hd__nand2_4 _40181_ (.A(_09396_),
    .B(_09147_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21o_4 _40182_ (.A1(_09391_),
    .A2(_09392_),
    .B1(_09394_),
    .X(_09650_));
 sky130_fd_sc_hd__nand2_4 _40183_ (.A(_09649_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__a21boi_4 _40184_ (.A1(_09647_),
    .A2(_09648_),
    .B1_N(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__xor2_4 _40185_ (.A(_09646_),
    .B(_09652_),
    .X(_01431_));
 sky130_fd_sc_hd__nand2_4 _40186_ (.A(_09520_),
    .B(_09516_),
    .Y(_09653_));
 sky130_vsdinv _40187_ (.A(_09653_),
    .Y(_09654_));
 sky130_vsdinv _40188_ (.A(_09482_),
    .Y(_09655_));
 sky130_fd_sc_hd__a21bo_4 _40189_ (.A1(_09655_),
    .A2(_09485_),
    .B1_N(_09487_),
    .X(_09656_));
 sky130_fd_sc_hd__nand2_4 _40190_ (.A(_06454_),
    .B(_07921_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand2_4 _40191_ (.A(_06842_),
    .B(_07712_),
    .Y(_09658_));
 sky130_fd_sc_hd__nand2_4 _40192_ (.A(_09657_),
    .B(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__nand4_4 _40193_ (.A(_07653_),
    .B(_06570_),
    .C(_08127_),
    .D(_08124_),
    .Y(_09660_));
 sky130_fd_sc_hd__nand2_4 _40194_ (.A(_07818_),
    .B(_07561_),
    .Y(_09661_));
 sky130_vsdinv _40195_ (.A(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__nand3_4 _40196_ (.A(_09659_),
    .B(_09660_),
    .C(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__nand2_4 _40197_ (.A(_09659_),
    .B(_09660_),
    .Y(_09664_));
 sky130_fd_sc_hd__nand2_4 _40198_ (.A(_09664_),
    .B(_09661_),
    .Y(_09665_));
 sky130_fd_sc_hd__nand3_4 _40199_ (.A(_09656_),
    .B(_09663_),
    .C(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__nand2_4 _40200_ (.A(_09665_),
    .B(_09663_),
    .Y(_09667_));
 sky130_fd_sc_hd__a21boi_4 _40201_ (.A1(_09485_),
    .A2(_09655_),
    .B1_N(_09487_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand2_4 _40202_ (.A(_09667_),
    .B(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__nand2_4 _40203_ (.A(_09666_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__a21boi_4 _40204_ (.A1(_09405_),
    .A2(_09410_),
    .B1_N(_09406_),
    .Y(_09671_));
 sky130_fd_sc_hd__nand2_4 _40205_ (.A(_09670_),
    .B(_09671_),
    .Y(_09672_));
 sky130_vsdinv _40206_ (.A(_09671_),
    .Y(_09673_));
 sky130_fd_sc_hd__nand3_4 _40207_ (.A(_09666_),
    .B(_09669_),
    .C(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__nand2_4 _40208_ (.A(_09672_),
    .B(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__a21boi_4 _40209_ (.A1(_09414_),
    .A2(_09423_),
    .B1_N(_09419_),
    .Y(_09676_));
 sky130_fd_sc_hd__nand2_4 _40210_ (.A(_09675_),
    .B(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__nand2_4 _40211_ (.A(_09424_),
    .B(_09419_),
    .Y(_09678_));
 sky130_fd_sc_hd__nand3_4 _40212_ (.A(_09678_),
    .B(_09672_),
    .C(_09674_),
    .Y(_09679_));
 sky130_fd_sc_hd__nand2_4 _40213_ (.A(_09677_),
    .B(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__nand2_4 _40214_ (.A(_07145_),
    .B(_07053_),
    .Y(_09681_));
 sky130_fd_sc_hd__nand2_4 _40215_ (.A(_07297_),
    .B(_07049_),
    .Y(_09682_));
 sky130_fd_sc_hd__nand2_4 _40216_ (.A(_09681_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__nand4_4 _40217_ (.A(_06998_),
    .B(_07297_),
    .C(_08953_),
    .D(_07733_),
    .Y(_09684_));
 sky130_fd_sc_hd__nand2_4 _40218_ (.A(_09683_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__nand2_4 _40219_ (.A(_07301_),
    .B(_07366_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand2_4 _40220_ (.A(_09685_),
    .B(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand4_4 _40221_ (.A(_08026_),
    .B(_09683_),
    .C(_09684_),
    .D(_08383_),
    .Y(_09688_));
 sky130_fd_sc_hd__nand2_4 _40222_ (.A(_09687_),
    .B(_09688_),
    .Y(_09689_));
 sky130_fd_sc_hd__a21boi_4 _40223_ (.A1(_09434_),
    .A2(_09439_),
    .B1_N(_09435_),
    .Y(_09690_));
 sky130_fd_sc_hd__nand2_4 _40224_ (.A(_09689_),
    .B(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__nand2_4 _40225_ (.A(_09440_),
    .B(_09435_),
    .Y(_09692_));
 sky130_fd_sc_hd__nand3_4 _40226_ (.A(_09692_),
    .B(_09688_),
    .C(_09687_),
    .Y(_09693_));
 sky130_fd_sc_hd__nand2_4 _40227_ (.A(_08050_),
    .B(_06750_),
    .Y(_09694_));
 sky130_fd_sc_hd__nand2_4 _40228_ (.A(_08289_),
    .B(_08162_),
    .Y(_09695_));
 sky130_fd_sc_hd__nand2_4 _40229_ (.A(_08291_),
    .B(_08164_),
    .Y(_09696_));
 sky130_fd_sc_hd__nand2_4 _40230_ (.A(_09695_),
    .B(_09696_),
    .Y(_09697_));
 sky130_fd_sc_hd__nand4_4 _40231_ (.A(_08294_),
    .B(_08291_),
    .C(_08164_),
    .D(_08162_),
    .Y(_09698_));
 sky130_fd_sc_hd__nand2_4 _40232_ (.A(_09697_),
    .B(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__xor2_4 _40233_ (.A(_09694_),
    .B(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__a21oi_4 _40234_ (.A1(_09691_),
    .A2(_09693_),
    .B1(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__nand3_4 _40235_ (.A(_09700_),
    .B(_09691_),
    .C(_09693_),
    .Y(_09702_));
 sky130_vsdinv _40236_ (.A(_09702_),
    .Y(_09703_));
 sky130_fd_sc_hd__nor2_4 _40237_ (.A(_09701_),
    .B(_09703_),
    .Y(_09704_));
 sky130_vsdinv _40238_ (.A(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__nand2_4 _40239_ (.A(_09680_),
    .B(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__nand3_4 _40240_ (.A(_09677_),
    .B(_09704_),
    .C(_09679_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand2_4 _40241_ (.A(_09706_),
    .B(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__nand2_4 _40242_ (.A(_09708_),
    .B(_09497_),
    .Y(_09709_));
 sky130_vsdinv _40243_ (.A(_09497_),
    .Y(_09710_));
 sky130_fd_sc_hd__nand3_4 _40244_ (.A(_09706_),
    .B(_09710_),
    .C(_09707_),
    .Y(_09711_));
 sky130_fd_sc_hd__nand2_4 _40245_ (.A(_09709_),
    .B(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__a21boi_4 _40246_ (.A1(_09427_),
    .A2(_09454_),
    .B1_N(_09429_),
    .Y(_09713_));
 sky130_fd_sc_hd__nand2_4 _40247_ (.A(_09712_),
    .B(_09713_),
    .Y(_09714_));
 sky130_vsdinv _40248_ (.A(_09713_),
    .Y(_09715_));
 sky130_fd_sc_hd__nand3_4 _40249_ (.A(_09709_),
    .B(_09715_),
    .C(_09711_),
    .Y(_09716_));
 sky130_fd_sc_hd__nand2_4 _40250_ (.A(_09714_),
    .B(_09716_),
    .Y(_09717_));
 sky130_fd_sc_hd__nand2_4 _40251_ (.A(_05950_),
    .B(_09467_),
    .Y(_09718_));
 sky130_fd_sc_hd__nand2_4 _40252_ (.A(_06018_),
    .B(_08629_),
    .Y(_09719_));
 sky130_fd_sc_hd__nand2_4 _40253_ (.A(_09718_),
    .B(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__nand4_4 _40254_ (.A(_07364_),
    .B(_06018_),
    .C(_03568_),
    .D(_09467_),
    .Y(_09721_));
 sky130_fd_sc_hd__nand2_4 _40255_ (.A(_09720_),
    .B(_09721_),
    .Y(_09722_));
 sky130_fd_sc_hd__nand2_4 _40256_ (.A(_06083_),
    .B(\pcpi_mul.rs2[21] ),
    .Y(_09723_));
 sky130_fd_sc_hd__nand2_4 _40257_ (.A(_09722_),
    .B(_09723_),
    .Y(_09724_));
 sky130_vsdinv _40258_ (.A(_09723_),
    .Y(_09725_));
 sky130_fd_sc_hd__nand3_4 _40259_ (.A(_09720_),
    .B(_09721_),
    .C(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand2_4 _40260_ (.A(_09724_),
    .B(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__a21boi_4 _40261_ (.A1(_09470_),
    .A2(_09473_),
    .B1_N(_09471_),
    .Y(_09728_));
 sky130_fd_sc_hd__nand2_4 _40262_ (.A(_09727_),
    .B(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__nand2_4 _40263_ (.A(_09475_),
    .B(_09471_),
    .Y(_09730_));
 sky130_fd_sc_hd__nand3_4 _40264_ (.A(_09730_),
    .B(_09726_),
    .C(_09724_),
    .Y(_09731_));
 sky130_fd_sc_hd__nand2_4 _40265_ (.A(_09729_),
    .B(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__nand2_4 _40266_ (.A(_06450_),
    .B(_08873_),
    .Y(_09733_));
 sky130_vsdinv _40267_ (.A(_09733_),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_4 _40268_ (.A(_06941_),
    .B(_08193_),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_4 _40269_ (.A(_08928_),
    .B(_09008_),
    .Y(_09736_));
 sky130_fd_sc_hd__nand2_4 _40270_ (.A(_09735_),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__nand4_4 _40271_ (.A(_06154_),
    .B(_06254_),
    .C(_09008_),
    .D(_08193_),
    .Y(_09738_));
 sky130_fd_sc_hd__nand2_4 _40272_ (.A(_09737_),
    .B(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__xor2_4 _40273_ (.A(_09734_),
    .B(_09739_),
    .X(_09740_));
 sky130_fd_sc_hd__nand2_4 _40274_ (.A(_09732_),
    .B(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__xor2_4 _40275_ (.A(_09733_),
    .B(_09739_),
    .X(_09742_));
 sky130_fd_sc_hd__nand3_4 _40276_ (.A(_09742_),
    .B(_09729_),
    .C(_09731_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand2_4 _40277_ (.A(_09741_),
    .B(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__nand3_4 _40278_ (.A(_09506_),
    .B(_09349_),
    .C(_09507_),
    .Y(_09745_));
 sky130_fd_sc_hd__nand2_4 _40279_ (.A(_09744_),
    .B(_09745_),
    .Y(_09746_));
 sky130_vsdinv _40280_ (.A(_09745_),
    .Y(_09747_));
 sky130_fd_sc_hd__nand3_4 _40281_ (.A(_09741_),
    .B(_09747_),
    .C(_09743_),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_4 _40282_ (.A(_09746_),
    .B(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__a21boi_4 _40283_ (.A1(_09478_),
    .A2(_09489_),
    .B1_N(_09480_),
    .Y(_09750_));
 sky130_fd_sc_hd__nand2_4 _40284_ (.A(_09749_),
    .B(_09750_),
    .Y(_09751_));
 sky130_vsdinv _40285_ (.A(_09750_),
    .Y(_09752_));
 sky130_fd_sc_hd__nand3_4 _40286_ (.A(_09746_),
    .B(_09752_),
    .C(_09748_),
    .Y(_09753_));
 sky130_fd_sc_hd__nand2_4 _40287_ (.A(_09751_),
    .B(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_4 _40288_ (.A(_05585_),
    .B(_03601_),
    .Y(_09755_));
 sky130_fd_sc_hd__buf_1 _40289_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09756_));
 sky130_fd_sc_hd__nand2_4 _40290_ (.A(_05965_),
    .B(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__nand2_4 _40291_ (.A(_05899_),
    .B(_03586_),
    .Y(_09758_));
 sky130_fd_sc_hd__nand2_4 _40292_ (.A(_09757_),
    .B(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__buf_1 _40293_ (.A(\pcpi_mul.rs2[25] ),
    .X(_09760_));
 sky130_fd_sc_hd__nand4_4 _40294_ (.A(_05884_),
    .B(_06126_),
    .C(_09760_),
    .D(_03595_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_4 _40295_ (.A(_06007_),
    .B(_09346_),
    .Y(_09762_));
 sky130_vsdinv _40296_ (.A(_09762_),
    .Y(_09763_));
 sky130_fd_sc_hd__a21o_4 _40297_ (.A1(_09759_),
    .A2(_09761_),
    .B1(_09763_),
    .X(_09764_));
 sky130_fd_sc_hd__nand3_4 _40298_ (.A(_09759_),
    .B(_09761_),
    .C(_09763_),
    .Y(_09765_));
 sky130_fd_sc_hd__nand2_4 _40299_ (.A(_09764_),
    .B(_09765_),
    .Y(_09766_));
 sky130_fd_sc_hd__a21boi_4 _40300_ (.A1(_09502_),
    .A2(_09505_),
    .B1_N(_09503_),
    .Y(_09767_));
 sky130_fd_sc_hd__nand2_4 _40301_ (.A(_09766_),
    .B(_09767_),
    .Y(_09768_));
 sky130_vsdinv _40302_ (.A(_09767_),
    .Y(_09769_));
 sky130_fd_sc_hd__nand3_4 _40303_ (.A(_09769_),
    .B(_09765_),
    .C(_09764_),
    .Y(_09770_));
 sky130_fd_sc_hd__nand2_4 _40304_ (.A(_09768_),
    .B(_09770_),
    .Y(_09771_));
 sky130_fd_sc_hd__xor2_4 _40305_ (.A(_09755_),
    .B(_09771_),
    .X(_09772_));
 sky130_vsdinv _40306_ (.A(_09772_),
    .Y(_09773_));
 sky130_fd_sc_hd__nand2_4 _40307_ (.A(_09754_),
    .B(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand3_4 _40308_ (.A(_09751_),
    .B(_09753_),
    .C(_09772_),
    .Y(_09775_));
 sky130_fd_sc_hd__nand2_4 _40309_ (.A(_09774_),
    .B(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__nand2_4 _40310_ (.A(_09776_),
    .B(_09512_),
    .Y(_09777_));
 sky130_vsdinv _40311_ (.A(_09512_),
    .Y(_09778_));
 sky130_fd_sc_hd__nand3_4 _40312_ (.A(_09774_),
    .B(_09778_),
    .C(_09775_),
    .Y(_09779_));
 sky130_fd_sc_hd__nand2_4 _40313_ (.A(_09777_),
    .B(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__nand2_4 _40314_ (.A(_09717_),
    .B(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand4_4 _40315_ (.A(_09716_),
    .B(_09714_),
    .C(_09777_),
    .D(_09779_),
    .Y(_09782_));
 sky130_fd_sc_hd__nand2_4 _40316_ (.A(_09781_),
    .B(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__nand2_4 _40317_ (.A(_09654_),
    .B(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__nand3_4 _40318_ (.A(_09653_),
    .B(_09782_),
    .C(_09781_),
    .Y(_09785_));
 sky130_fd_sc_hd__nand2_4 _40319_ (.A(_09784_),
    .B(_09785_),
    .Y(_09786_));
 sky130_fd_sc_hd__nand2_4 _40320_ (.A(_09554_),
    .B(_09549_),
    .Y(_09787_));
 sky130_vsdinv _40321_ (.A(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__nand2_4 _40322_ (.A(_03340_),
    .B(_06592_),
    .Y(_09789_));
 sky130_fd_sc_hd__nand2_4 _40323_ (.A(_08054_),
    .B(_06598_),
    .Y(_09790_));
 sky130_fd_sc_hd__nand2_4 _40324_ (.A(_09789_),
    .B(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand4_4 _40325_ (.A(_08045_),
    .B(_03346_),
    .C(_07095_),
    .D(_03490_),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_4 _40326_ (.A(_09791_),
    .B(_09792_),
    .Y(_09793_));
 sky130_fd_sc_hd__nand2_4 _40327_ (.A(_08313_),
    .B(_03475_),
    .Y(_09794_));
 sky130_fd_sc_hd__nand2_4 _40328_ (.A(_09793_),
    .B(_09794_),
    .Y(_09795_));
 sky130_vsdinv _40329_ (.A(_09794_),
    .Y(_09796_));
 sky130_fd_sc_hd__nand3_4 _40330_ (.A(_09791_),
    .B(_09792_),
    .C(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__nand2_4 _40331_ (.A(_09795_),
    .B(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__maj3_4 _40332_ (.A(_09444_),
    .B(_09445_),
    .C(_09446_),
    .X(_09799_));
 sky130_fd_sc_hd__nand2_4 _40333_ (.A(_09798_),
    .B(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__a22oi_4 _40334_ (.A1(_07305_),
    .A2(_07214_),
    .B1(_07435_),
    .B2(_07956_),
    .Y(_09801_));
 sky130_fd_sc_hd__o21ai_4 _40335_ (.A1(_09444_),
    .A2(_09801_),
    .B1(_09448_),
    .Y(_09802_));
 sky130_fd_sc_hd__nand3_4 _40336_ (.A(_09802_),
    .B(_09797_),
    .C(_09795_),
    .Y(_09803_));
 sky130_fd_sc_hd__nand2_4 _40337_ (.A(_09800_),
    .B(_09803_),
    .Y(_09804_));
 sky130_fd_sc_hd__a21boi_4 _40338_ (.A1(_09527_),
    .A2(_09532_),
    .B1_N(_09528_),
    .Y(_09805_));
 sky130_fd_sc_hd__nand2_4 _40339_ (.A(_09804_),
    .B(_09805_),
    .Y(_09806_));
 sky130_vsdinv _40340_ (.A(_09805_),
    .Y(_09807_));
 sky130_fd_sc_hd__nand3_4 _40341_ (.A(_09800_),
    .B(_09803_),
    .C(_09807_),
    .Y(_09808_));
 sky130_fd_sc_hd__nand2_4 _40342_ (.A(_09806_),
    .B(_09808_),
    .Y(_09809_));
 sky130_vsdinv _40343_ (.A(_09443_),
    .Y(_09810_));
 sky130_fd_sc_hd__a21oi_4 _40344_ (.A1(_09450_),
    .A2(_09442_),
    .B1(_09810_),
    .Y(_09811_));
 sky130_fd_sc_hd__nand2_4 _40345_ (.A(_09809_),
    .B(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__a21o_4 _40346_ (.A1(_09450_),
    .A2(_09442_),
    .B1(_09810_),
    .X(_09813_));
 sky130_fd_sc_hd__nand3_4 _40347_ (.A(_09813_),
    .B(_09808_),
    .C(_09806_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2_4 _40348_ (.A(_09812_),
    .B(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__a21boi_4 _40349_ (.A1(_09536_),
    .A2(_09543_),
    .B1_N(_09539_),
    .Y(_09816_));
 sky130_fd_sc_hd__nand2_4 _40350_ (.A(_09815_),
    .B(_09816_),
    .Y(_09817_));
 sky130_vsdinv _40351_ (.A(_09816_),
    .Y(_09818_));
 sky130_fd_sc_hd__nand3_4 _40352_ (.A(_09812_),
    .B(_09814_),
    .C(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__nand2_4 _40353_ (.A(_09817_),
    .B(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__nand2_4 _40354_ (.A(_09788_),
    .B(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__nand3_4 _40355_ (.A(_09787_),
    .B(_09817_),
    .C(_09819_),
    .Y(_09822_));
 sky130_fd_sc_hd__nand2_4 _40356_ (.A(_09821_),
    .B(_09822_),
    .Y(_09823_));
 sky130_vsdinv _40357_ (.A(_09573_),
    .Y(_09824_));
 sky130_fd_sc_hd__a21oi_4 _40358_ (.A1(_09572_),
    .A2(_09586_),
    .B1(_09824_),
    .Y(_09825_));
 sky130_vsdinv _40359_ (.A(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__nand2_4 _40360_ (.A(_09202_),
    .B(_06052_),
    .Y(_09827_));
 sky130_fd_sc_hd__nand2_4 _40361_ (.A(_09565_),
    .B(_06056_),
    .Y(_09828_));
 sky130_fd_sc_hd__nand2_4 _40362_ (.A(_09827_),
    .B(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__buf_1 _40363_ (.A(_09086_),
    .X(_09830_));
 sky130_fd_sc_hd__buf_1 _40364_ (.A(_08758_),
    .X(_09831_));
 sky130_fd_sc_hd__nand4_4 _40365_ (.A(_09830_),
    .B(_09831_),
    .C(_05963_),
    .D(_05989_),
    .Y(_09832_));
 sky130_fd_sc_hd__buf_1 _40366_ (.A(\pcpi_mul.rs1[24] ),
    .X(_09833_));
 sky130_fd_sc_hd__nand2_4 _40367_ (.A(_09833_),
    .B(_05967_),
    .Y(_09834_));
 sky130_vsdinv _40368_ (.A(_09834_),
    .Y(_09835_));
 sky130_fd_sc_hd__a21o_4 _40369_ (.A1(_09829_),
    .A2(_09832_),
    .B1(_09835_),
    .X(_09836_));
 sky130_fd_sc_hd__nand3_4 _40370_ (.A(_09829_),
    .B(_09832_),
    .C(_09835_),
    .Y(_09837_));
 sky130_fd_sc_hd__a21boi_4 _40371_ (.A1(_09563_),
    .A2(_09567_),
    .B1_N(_09564_),
    .Y(_09838_));
 sky130_fd_sc_hd__a21boi_4 _40372_ (.A1(_09836_),
    .A2(_09837_),
    .B1_N(_09838_),
    .Y(_09839_));
 sky130_vsdinv _40373_ (.A(_09838_),
    .Y(_09840_));
 sky130_fd_sc_hd__nand3_4 _40374_ (.A(_09840_),
    .B(_09837_),
    .C(_09836_),
    .Y(_09841_));
 sky130_vsdinv _40375_ (.A(_09841_),
    .Y(_09842_));
 sky130_fd_sc_hd__buf_1 _40376_ (.A(_03374_),
    .X(_09843_));
 sky130_fd_sc_hd__nand2_4 _40377_ (.A(_09843_),
    .B(_08043_),
    .Y(_09844_));
 sky130_fd_sc_hd__o21ai_4 _40378_ (.A1(_03380_),
    .A2(_05892_),
    .B1(_09844_),
    .Y(_09845_));
 sky130_fd_sc_hd__buf_1 _40379_ (.A(_03374_),
    .X(_09846_));
 sky130_fd_sc_hd__buf_1 _40380_ (.A(_03379_),
    .X(_09847_));
 sky130_fd_sc_hd__nand4_4 _40381_ (.A(_09846_),
    .B(_09847_),
    .C(_07440_),
    .D(_03443_),
    .Y(_09848_));
 sky130_fd_sc_hd__buf_1 _40382_ (.A(\pcpi_mul.rs1[27] ),
    .X(_09849_));
 sky130_fd_sc_hd__nand2_4 _40383_ (.A(_09849_),
    .B(_06853_),
    .Y(_09850_));
 sky130_vsdinv _40384_ (.A(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__a21oi_4 _40385_ (.A1(_09845_),
    .A2(_09848_),
    .B1(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__nand3_4 _40386_ (.A(_09845_),
    .B(_09848_),
    .C(_09851_),
    .Y(_09853_));
 sky130_vsdinv _40387_ (.A(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__nor2_4 _40388_ (.A(_09852_),
    .B(_09854_),
    .Y(_09855_));
 sky130_vsdinv _40389_ (.A(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__o21ai_4 _40390_ (.A1(_09839_),
    .A2(_09842_),
    .B1(_09856_),
    .Y(_09857_));
 sky130_vsdinv _40391_ (.A(_09839_),
    .Y(_09858_));
 sky130_fd_sc_hd__nand3_4 _40392_ (.A(_09858_),
    .B(_09855_),
    .C(_09841_),
    .Y(_09859_));
 sky130_fd_sc_hd__nand3_4 _40393_ (.A(_09826_),
    .B(_09857_),
    .C(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__nand2_4 _40394_ (.A(_09857_),
    .B(_09859_),
    .Y(_09861_));
 sky130_fd_sc_hd__nand2_4 _40395_ (.A(_09861_),
    .B(_09825_),
    .Y(_09862_));
 sky130_fd_sc_hd__a21boi_4 _40396_ (.A1(_09576_),
    .A2(_09582_),
    .B1_N(_09579_),
    .Y(_09863_));
 sky130_vsdinv _40397_ (.A(_09863_),
    .Y(_09864_));
 sky130_fd_sc_hd__a21oi_4 _40398_ (.A1(_09860_),
    .A2(_09862_),
    .B1(_09864_),
    .Y(_09865_));
 sky130_vsdinv _40399_ (.A(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__nand3_4 _40400_ (.A(_09860_),
    .B(_09862_),
    .C(_09864_),
    .Y(_09867_));
 sky130_fd_sc_hd__nand2_4 _40401_ (.A(_09866_),
    .B(_09867_),
    .Y(_09868_));
 sky130_fd_sc_hd__nand2_4 _40402_ (.A(_09823_),
    .B(_09868_),
    .Y(_09869_));
 sky130_vsdinv _40403_ (.A(_09867_),
    .Y(_09870_));
 sky130_fd_sc_hd__nor2_4 _40404_ (.A(_09865_),
    .B(_09870_),
    .Y(_09871_));
 sky130_fd_sc_hd__nand3_4 _40405_ (.A(_09871_),
    .B(_09822_),
    .C(_09821_),
    .Y(_09872_));
 sky130_fd_sc_hd__nand2_4 _40406_ (.A(_09869_),
    .B(_09872_),
    .Y(_09873_));
 sky130_vsdinv _40407_ (.A(_09460_),
    .Y(_09874_));
 sky130_fd_sc_hd__a21oi_4 _40408_ (.A1(_09458_),
    .A2(_09464_),
    .B1(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__nand2_4 _40409_ (.A(_09873_),
    .B(_09875_),
    .Y(_09876_));
 sky130_fd_sc_hd__a21o_4 _40410_ (.A1(_09458_),
    .A2(_09464_),
    .B1(_09874_),
    .X(_09877_));
 sky130_fd_sc_hd__nand3_4 _40411_ (.A(_09877_),
    .B(_09872_),
    .C(_09869_),
    .Y(_09878_));
 sky130_fd_sc_hd__nand2_4 _40412_ (.A(_09876_),
    .B(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__a21boi_4 _40413_ (.A1(_09602_),
    .A2(_09557_),
    .B1_N(_09559_),
    .Y(_09880_));
 sky130_fd_sc_hd__nand2_4 _40414_ (.A(_09879_),
    .B(_09880_),
    .Y(_09881_));
 sky130_vsdinv _40415_ (.A(_09880_),
    .Y(_09882_));
 sky130_fd_sc_hd__nand3_4 _40416_ (.A(_09876_),
    .B(_09878_),
    .C(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__nand2_4 _40417_ (.A(_09881_),
    .B(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__nand2_4 _40418_ (.A(_09786_),
    .B(_09884_),
    .Y(_09885_));
 sky130_fd_sc_hd__nand4_4 _40419_ (.A(_09883_),
    .B(_09784_),
    .C(_09881_),
    .D(_09785_),
    .Y(_09886_));
 sky130_fd_sc_hd__nand2_4 _40420_ (.A(_09885_),
    .B(_09886_),
    .Y(_09887_));
 sky130_fd_sc_hd__a21oi_4 _40421_ (.A1(_09519_),
    .A2(_09520_),
    .B1(_09401_),
    .Y(_09888_));
 sky130_fd_sc_hd__o21a_4 _40422_ (.A1(_09888_),
    .A2(_09615_),
    .B1(_09523_),
    .X(_09889_));
 sky130_fd_sc_hd__nand2_4 _40423_ (.A(_09887_),
    .B(_09889_),
    .Y(_09890_));
 sky130_fd_sc_hd__o21ai_4 _40424_ (.A1(_09888_),
    .A2(_09615_),
    .B1(_09523_),
    .Y(_09891_));
 sky130_fd_sc_hd__nand3_4 _40425_ (.A(_09891_),
    .B(_09886_),
    .C(_09885_),
    .Y(_09892_));
 sky130_fd_sc_hd__nand2_4 _40426_ (.A(_09890_),
    .B(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__a21boi_4 _40427_ (.A1(_09592_),
    .A2(_09595_),
    .B1_N(_09593_),
    .Y(_09894_));
 sky130_fd_sc_hd__nand2_4 _40428_ (.A(_09614_),
    .B(_09609_),
    .Y(_09895_));
 sky130_fd_sc_hd__xor2_4 _40429_ (.A(_09894_),
    .B(_09895_),
    .X(_09896_));
 sky130_fd_sc_hd__nand2_4 _40430_ (.A(_09893_),
    .B(_09896_),
    .Y(_09897_));
 sky130_vsdinv _40431_ (.A(_09896_),
    .Y(_09898_));
 sky130_fd_sc_hd__nand3_4 _40432_ (.A(_09898_),
    .B(_09890_),
    .C(_09892_),
    .Y(_09899_));
 sky130_fd_sc_hd__nand2_4 _40433_ (.A(_09897_),
    .B(_09899_),
    .Y(_09900_));
 sky130_fd_sc_hd__a21boi_4 _40434_ (.A1(_09619_),
    .A2(_09627_),
    .B1_N(_09621_),
    .Y(_09901_));
 sky130_fd_sc_hd__nand2_4 _40435_ (.A(_09900_),
    .B(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__nand2_4 _40436_ (.A(_09628_),
    .B(_09621_),
    .Y(_09903_));
 sky130_fd_sc_hd__nand3_4 _40437_ (.A(_09903_),
    .B(_09899_),
    .C(_09897_),
    .Y(_09904_));
 sky130_fd_sc_hd__nand2_4 _40438_ (.A(_09902_),
    .B(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__a21oi_4 _40439_ (.A1(_09245_),
    .A2(_09243_),
    .B1(_09623_),
    .Y(_09906_));
 sky130_vsdinv _40440_ (.A(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__nand2_4 _40441_ (.A(_09905_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__nand3_4 _40442_ (.A(_09902_),
    .B(_09904_),
    .C(_09906_),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_4 _40443_ (.A(_09908_),
    .B(_09909_),
    .Y(_09910_));
 sky130_fd_sc_hd__a21boi_4 _40444_ (.A1(_09631_),
    .A2(_09635_),
    .B1_N(_09633_),
    .Y(_09911_));
 sky130_fd_sc_hd__nand2_4 _40445_ (.A(_09910_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__nand2_4 _40446_ (.A(_09638_),
    .B(_09633_),
    .Y(_09913_));
 sky130_fd_sc_hd__nand3_4 _40447_ (.A(_09913_),
    .B(_09908_),
    .C(_09909_),
    .Y(_09914_));
 sky130_fd_sc_hd__and2_4 _40448_ (.A(_09912_),
    .B(_09914_),
    .X(_09915_));
 sky130_fd_sc_hd__buf_1 _40449_ (.A(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__o21ai_4 _40450_ (.A1(_09646_),
    .A2(_09652_),
    .B1(_09643_),
    .Y(_09917_));
 sky130_fd_sc_hd__xor2_4 _40451_ (.A(_09916_),
    .B(_09917_),
    .X(_01432_));
 sky130_fd_sc_hd__o21a_4 _40452_ (.A1(_09884_),
    .A2(_09786_),
    .B1(_09785_),
    .X(_09918_));
 sky130_fd_sc_hd__nand2_4 _40453_ (.A(_06842_),
    .B(_03539_),
    .Y(_09919_));
 sky130_fd_sc_hd__nand2_4 _40454_ (.A(_03302_),
    .B(_03534_),
    .Y(_09920_));
 sky130_fd_sc_hd__nand2_4 _40455_ (.A(_09919_),
    .B(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__nand4_4 _40456_ (.A(_06570_),
    .B(_07818_),
    .C(_08571_),
    .D(_07709_),
    .Y(_09922_));
 sky130_fd_sc_hd__nand2_4 _40457_ (.A(_09921_),
    .B(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_4 _40458_ (.A(_07145_),
    .B(\pcpi_mul.rs2[15] ),
    .Y(_09924_));
 sky130_fd_sc_hd__nand2_4 _40459_ (.A(_09923_),
    .B(_09924_),
    .Y(_09925_));
 sky130_vsdinv _40460_ (.A(_09924_),
    .Y(_09926_));
 sky130_fd_sc_hd__nand3_4 _40461_ (.A(_09921_),
    .B(_09922_),
    .C(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__nand2_4 _40462_ (.A(_09925_),
    .B(_09927_),
    .Y(_09928_));
 sky130_fd_sc_hd__a21boi_4 _40463_ (.A1(_09737_),
    .A2(_09734_),
    .B1_N(_09738_),
    .Y(_09929_));
 sky130_fd_sc_hd__nand2_4 _40464_ (.A(_09928_),
    .B(_09929_),
    .Y(_09930_));
 sky130_vsdinv _40465_ (.A(_09738_),
    .Y(_09931_));
 sky130_fd_sc_hd__a21o_4 _40466_ (.A1(_09737_),
    .A2(_09734_),
    .B1(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__nand3_4 _40467_ (.A(_09932_),
    .B(_09927_),
    .C(_09925_),
    .Y(_09933_));
 sky130_fd_sc_hd__nand2_4 _40468_ (.A(_09930_),
    .B(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__a21boi_4 _40469_ (.A1(_09659_),
    .A2(_09662_),
    .B1_N(_09660_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_4 _40470_ (.A(_09934_),
    .B(_09935_),
    .Y(_09936_));
 sky130_vsdinv _40471_ (.A(_09935_),
    .Y(_09937_));
 sky130_fd_sc_hd__nand3_4 _40472_ (.A(_09930_),
    .B(_09933_),
    .C(_09937_),
    .Y(_09938_));
 sky130_fd_sc_hd__nand2_4 _40473_ (.A(_09936_),
    .B(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__a21boi_4 _40474_ (.A1(_09669_),
    .A2(_09673_),
    .B1_N(_09666_),
    .Y(_09940_));
 sky130_fd_sc_hd__nand2_4 _40475_ (.A(_09939_),
    .B(_09940_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_4 _40476_ (.A(_09674_),
    .B(_09666_),
    .Y(_09942_));
 sky130_fd_sc_hd__nand3_4 _40477_ (.A(_09942_),
    .B(_09938_),
    .C(_09936_),
    .Y(_09943_));
 sky130_fd_sc_hd__nand2_4 _40478_ (.A(_09941_),
    .B(_09943_),
    .Y(_09944_));
 sky130_fd_sc_hd__nand2_4 _40479_ (.A(_03313_),
    .B(_07361_),
    .Y(_09945_));
 sky130_fd_sc_hd__nand2_4 _40480_ (.A(_07156_),
    .B(_08953_),
    .Y(_09946_));
 sky130_fd_sc_hd__nand2_4 _40481_ (.A(_09945_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__nand4_4 _40482_ (.A(_06991_),
    .B(_07438_),
    .C(_07058_),
    .D(_07054_),
    .Y(_09948_));
 sky130_fd_sc_hd__nand2_4 _40483_ (.A(_08294_),
    .B(_07366_),
    .Y(_09949_));
 sky130_fd_sc_hd__a21bo_4 _40484_ (.A1(_09947_),
    .A2(_09948_),
    .B1_N(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__nand4_4 _40485_ (.A(_03325_),
    .B(_09947_),
    .C(_09948_),
    .D(_07045_),
    .Y(_09951_));
 sky130_fd_sc_hd__nand2_4 _40486_ (.A(_09950_),
    .B(_09951_),
    .Y(_09952_));
 sky130_fd_sc_hd__maj3_4 _40487_ (.A(_09686_),
    .B(_09681_),
    .C(_09682_),
    .X(_09953_));
 sky130_fd_sc_hd__nand2_4 _40488_ (.A(_09952_),
    .B(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__nand2_4 _40489_ (.A(_09688_),
    .B(_09684_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand3_4 _40490_ (.A(_09955_),
    .B(_09951_),
    .C(_09950_),
    .Y(_09956_));
 sky130_fd_sc_hd__nand2_4 _40491_ (.A(_03341_),
    .B(_07204_),
    .Y(_09957_));
 sky130_fd_sc_hd__nand2_4 _40492_ (.A(_03331_),
    .B(_07343_),
    .Y(_09958_));
 sky130_fd_sc_hd__nand2_4 _40493_ (.A(_07870_),
    .B(_07211_),
    .Y(_09959_));
 sky130_fd_sc_hd__nand2_4 _40494_ (.A(_09958_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__nand4_4 _40495_ (.A(_08291_),
    .B(_03336_),
    .C(_08164_),
    .D(_06747_),
    .Y(_09961_));
 sky130_fd_sc_hd__nand2_4 _40496_ (.A(_09960_),
    .B(_09961_),
    .Y(_09962_));
 sky130_fd_sc_hd__xor2_4 _40497_ (.A(_09957_),
    .B(_09962_),
    .X(_09963_));
 sky130_fd_sc_hd__a21oi_4 _40498_ (.A1(_09954_),
    .A2(_09956_),
    .B1(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__nand3_4 _40499_ (.A(_09954_),
    .B(_09963_),
    .C(_09956_),
    .Y(_09965_));
 sky130_vsdinv _40500_ (.A(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__nor2_4 _40501_ (.A(_09964_),
    .B(_09966_),
    .Y(_09967_));
 sky130_vsdinv _40502_ (.A(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__nand2_4 _40503_ (.A(_09944_),
    .B(_09968_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand3_4 _40504_ (.A(_09941_),
    .B(_09967_),
    .C(_09943_),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_4 _40505_ (.A(_09969_),
    .B(_09970_),
    .Y(_09971_));
 sky130_vsdinv _40506_ (.A(_09748_),
    .Y(_09972_));
 sky130_fd_sc_hd__a21oi_4 _40507_ (.A1(_09746_),
    .A2(_09752_),
    .B1(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__nand2_4 _40508_ (.A(_09971_),
    .B(_09973_),
    .Y(_09974_));
 sky130_vsdinv _40509_ (.A(_09973_),
    .Y(_09975_));
 sky130_fd_sc_hd__nand3_4 _40510_ (.A(_09975_),
    .B(_09970_),
    .C(_09969_),
    .Y(_09976_));
 sky130_fd_sc_hd__nand2_4 _40511_ (.A(_09974_),
    .B(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__a21boi_4 _40512_ (.A1(_09677_),
    .A2(_09704_),
    .B1_N(_09679_),
    .Y(_09978_));
 sky130_fd_sc_hd__nand2_4 _40513_ (.A(_09977_),
    .B(_09978_),
    .Y(_09979_));
 sky130_vsdinv _40514_ (.A(_09978_),
    .Y(_09980_));
 sky130_fd_sc_hd__nand3_4 _40515_ (.A(_09974_),
    .B(_09976_),
    .C(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__nand2_4 _40516_ (.A(_09979_),
    .B(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__nand2_4 _40517_ (.A(_03268_),
    .B(_03575_),
    .Y(_09983_));
 sky130_fd_sc_hd__nand2_4 _40518_ (.A(_06243_),
    .B(_03568_),
    .Y(_09984_));
 sky130_fd_sc_hd__nand2_4 _40519_ (.A(_09983_),
    .B(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__nand4_4 _40520_ (.A(_06159_),
    .B(_06243_),
    .C(_08995_),
    .D(_08862_),
    .Y(_09986_));
 sky130_fd_sc_hd__nand2_4 _40521_ (.A(_09985_),
    .B(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_4 _40522_ (.A(_03274_),
    .B(_03562_),
    .Y(_09988_));
 sky130_fd_sc_hd__nand2_4 _40523_ (.A(_09987_),
    .B(_09988_),
    .Y(_09989_));
 sky130_vsdinv _40524_ (.A(_09988_),
    .Y(_09990_));
 sky130_fd_sc_hd__nand3_4 _40525_ (.A(_09985_),
    .B(_09986_),
    .C(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__nand2_4 _40526_ (.A(_09989_),
    .B(_09991_),
    .Y(_09992_));
 sky130_fd_sc_hd__a21boi_4 _40527_ (.A1(_09720_),
    .A2(_09725_),
    .B1_N(_09721_),
    .Y(_09993_));
 sky130_fd_sc_hd__nand2_4 _40528_ (.A(_09992_),
    .B(_09993_),
    .Y(_09994_));
 sky130_fd_sc_hd__nand2_4 _40529_ (.A(_09726_),
    .B(_09721_),
    .Y(_09995_));
 sky130_fd_sc_hd__nand3_4 _40530_ (.A(_09995_),
    .B(_09991_),
    .C(_09989_),
    .Y(_09996_));
 sky130_fd_sc_hd__nand2_4 _40531_ (.A(_09994_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_4 _40532_ (.A(_07653_),
    .B(_08640_),
    .Y(_09998_));
 sky130_vsdinv _40533_ (.A(_09998_),
    .Y(_09999_));
 sky130_fd_sc_hd__nand2_4 _40534_ (.A(_06549_),
    .B(_08647_),
    .Y(_10000_));
 sky130_fd_sc_hd__nand2_4 _40535_ (.A(_08167_),
    .B(_08646_),
    .Y(_10001_));
 sky130_fd_sc_hd__nand2_4 _40536_ (.A(_10000_),
    .B(_10001_),
    .Y(_10002_));
 sky130_fd_sc_hd__nand4_4 _40537_ (.A(_03280_),
    .B(_08167_),
    .C(_08646_),
    .D(_08647_),
    .Y(_10003_));
 sky130_fd_sc_hd__nand2_4 _40538_ (.A(_10002_),
    .B(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__xor2_4 _40539_ (.A(_09999_),
    .B(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__nand2_4 _40540_ (.A(_09997_),
    .B(_10005_),
    .Y(_10006_));
 sky130_fd_sc_hd__xor2_4 _40541_ (.A(_09998_),
    .B(_10004_),
    .X(_10007_));
 sky130_fd_sc_hd__nand3_4 _40542_ (.A(_10007_),
    .B(_09994_),
    .C(_09996_),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_4 _40543_ (.A(_10006_),
    .B(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__nand2_4 _40544_ (.A(_10009_),
    .B(_09770_),
    .Y(_10010_));
 sky130_vsdinv _40545_ (.A(_09770_),
    .Y(_10011_));
 sky130_fd_sc_hd__nand3_4 _40546_ (.A(_10006_),
    .B(_10011_),
    .C(_10008_),
    .Y(_10012_));
 sky130_fd_sc_hd__nand2_4 _40547_ (.A(_10010_),
    .B(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__a21boi_4 _40548_ (.A1(_09742_),
    .A2(_09729_),
    .B1_N(_09731_),
    .Y(_10014_));
 sky130_fd_sc_hd__nand2_4 _40549_ (.A(_10013_),
    .B(_10014_),
    .Y(_10015_));
 sky130_vsdinv _40550_ (.A(_10014_),
    .Y(_10016_));
 sky130_fd_sc_hd__nand3_4 _40551_ (.A(_10010_),
    .B(_10016_),
    .C(_10012_),
    .Y(_10017_));
 sky130_fd_sc_hd__nand2_4 _40552_ (.A(_10015_),
    .B(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__nand2_4 _40553_ (.A(_06126_),
    .B(_09756_),
    .Y(_10019_));
 sky130_fd_sc_hd__nand2_4 _40554_ (.A(_03256_),
    .B(_03586_),
    .Y(_10020_));
 sky130_fd_sc_hd__nand2_4 _40555_ (.A(_10019_),
    .B(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__nand4_4 _40556_ (.A(_05935_),
    .B(_05942_),
    .C(_09343_),
    .D(_03595_),
    .Y(_10022_));
 sky130_fd_sc_hd__nand2_4 _40557_ (.A(_10021_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__nand2_4 _40558_ (.A(_03261_),
    .B(_03580_),
    .Y(_10024_));
 sky130_fd_sc_hd__nand2_4 _40559_ (.A(_10023_),
    .B(_10024_),
    .Y(_10025_));
 sky130_vsdinv _40560_ (.A(_10024_),
    .Y(_10026_));
 sky130_fd_sc_hd__nand3_4 _40561_ (.A(_10021_),
    .B(_10022_),
    .C(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__nand2_4 _40562_ (.A(_10025_),
    .B(_10027_),
    .Y(_10028_));
 sky130_fd_sc_hd__a21boi_4 _40563_ (.A1(_09759_),
    .A2(_09763_),
    .B1_N(_09761_),
    .Y(_10029_));
 sky130_fd_sc_hd__nand2_4 _40564_ (.A(_10028_),
    .B(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__nand2_4 _40565_ (.A(_09765_),
    .B(_09761_),
    .Y(_10031_));
 sky130_fd_sc_hd__nand3_4 _40566_ (.A(_10031_),
    .B(_10027_),
    .C(_10025_),
    .Y(_10032_));
 sky130_fd_sc_hd__nand2_4 _40567_ (.A(_10030_),
    .B(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__nand2_4 _40568_ (.A(_05583_),
    .B(_03605_),
    .Y(_10034_));
 sky130_fd_sc_hd__buf_1 _40569_ (.A(\pcpi_mul.rs2[27] ),
    .X(_10035_));
 sky130_fd_sc_hd__nand2_4 _40570_ (.A(_05965_),
    .B(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__nor2_4 _40571_ (.A(_10034_),
    .B(_10036_),
    .Y(_10037_));
 sky130_vsdinv _40572_ (.A(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__nand2_4 _40573_ (.A(_10034_),
    .B(_10036_),
    .Y(_10039_));
 sky130_fd_sc_hd__nand2_4 _40574_ (.A(_10038_),
    .B(_10039_),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_4 _40575_ (.A(_10033_),
    .B(_10040_),
    .Y(_10041_));
 sky130_vsdinv _40576_ (.A(_10040_),
    .Y(_10042_));
 sky130_fd_sc_hd__nand3_4 _40577_ (.A(_10030_),
    .B(_10042_),
    .C(_10032_),
    .Y(_10043_));
 sky130_fd_sc_hd__nand2_4 _40578_ (.A(_10041_),
    .B(_10043_),
    .Y(_10044_));
 sky130_vsdinv _40579_ (.A(_09755_),
    .Y(_10045_));
 sky130_fd_sc_hd__nand3_4 _40580_ (.A(_09768_),
    .B(_09770_),
    .C(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__nand2_4 _40581_ (.A(_10044_),
    .B(_10046_),
    .Y(_10047_));
 sky130_vsdinv _40582_ (.A(_10046_),
    .Y(_10048_));
 sky130_fd_sc_hd__nand3_4 _40583_ (.A(_10048_),
    .B(_10041_),
    .C(_10043_),
    .Y(_10049_));
 sky130_fd_sc_hd__and2_4 _40584_ (.A(_10047_),
    .B(_10049_),
    .X(_10050_));
 sky130_vsdinv _40585_ (.A(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__nand2_4 _40586_ (.A(_10018_),
    .B(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__nand3_4 _40587_ (.A(_10015_),
    .B(_10050_),
    .C(_10017_),
    .Y(_10053_));
 sky130_fd_sc_hd__nand2_4 _40588_ (.A(_10052_),
    .B(_10053_),
    .Y(_10054_));
 sky130_fd_sc_hd__nand2_4 _40589_ (.A(_10054_),
    .B(_09775_),
    .Y(_10055_));
 sky130_vsdinv _40590_ (.A(_09775_),
    .Y(_10056_));
 sky130_fd_sc_hd__nand3_4 _40591_ (.A(_10056_),
    .B(_10052_),
    .C(_10053_),
    .Y(_10057_));
 sky130_fd_sc_hd__nand2_4 _40592_ (.A(_10055_),
    .B(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__nand2_4 _40593_ (.A(_09982_),
    .B(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__nand4_4 _40594_ (.A(_09981_),
    .B(_09979_),
    .C(_10055_),
    .D(_10057_),
    .Y(_10060_));
 sky130_fd_sc_hd__nand2_4 _40595_ (.A(_10059_),
    .B(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__nand3_4 _40596_ (.A(_10061_),
    .B(_09779_),
    .C(_09782_),
    .Y(_10062_));
 sky130_fd_sc_hd__nand2_4 _40597_ (.A(_09782_),
    .B(_09779_),
    .Y(_10063_));
 sky130_fd_sc_hd__buf_1 _40598_ (.A(_10060_),
    .X(_10064_));
 sky130_fd_sc_hd__nand3_4 _40599_ (.A(_10063_),
    .B(_10064_),
    .C(_10059_),
    .Y(_10065_));
 sky130_fd_sc_hd__nand2_4 _40600_ (.A(_10062_),
    .B(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__nand2_4 _40601_ (.A(_08759_),
    .B(_06322_),
    .Y(_10067_));
 sky130_fd_sc_hd__nand2_4 _40602_ (.A(_09833_),
    .B(_08028_),
    .Y(_10068_));
 sky130_fd_sc_hd__nand2_4 _40603_ (.A(_10067_),
    .B(_10068_),
    .Y(_10069_));
 sky130_fd_sc_hd__nand4_4 _40604_ (.A(_08759_),
    .B(_09212_),
    .C(_06059_),
    .D(_06431_),
    .Y(_10070_));
 sky130_fd_sc_hd__nand2_4 _40605_ (.A(_03375_),
    .B(_03453_),
    .Y(_10071_));
 sky130_vsdinv _40606_ (.A(_10071_),
    .Y(_10072_));
 sky130_fd_sc_hd__a21o_4 _40607_ (.A1(_10069_),
    .A2(_10070_),
    .B1(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__nand3_4 _40608_ (.A(_10069_),
    .B(_10070_),
    .C(_10072_),
    .Y(_10074_));
 sky130_fd_sc_hd__nand2_4 _40609_ (.A(_10073_),
    .B(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__a21boi_4 _40610_ (.A1(_09829_),
    .A2(_09835_),
    .B1_N(_09832_),
    .Y(_10076_));
 sky130_fd_sc_hd__nand2_4 _40611_ (.A(_10075_),
    .B(_10076_),
    .Y(_10077_));
 sky130_vsdinv _40612_ (.A(_10076_),
    .Y(_10078_));
 sky130_fd_sc_hd__nand3_4 _40613_ (.A(_10078_),
    .B(_10074_),
    .C(_10073_),
    .Y(_10079_));
 sky130_fd_sc_hd__buf_1 _40614_ (.A(_03379_),
    .X(_10080_));
 sky130_fd_sc_hd__nand2_4 _40615_ (.A(_10080_),
    .B(_05910_),
    .Y(_10081_));
 sky130_fd_sc_hd__o21ai_4 _40616_ (.A1(_03384_),
    .A2(_07144_),
    .B1(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__buf_1 _40617_ (.A(\pcpi_mul.rs1[26] ),
    .X(_10083_));
 sky130_fd_sc_hd__buf_1 _40618_ (.A(_10083_),
    .X(_10084_));
 sky130_fd_sc_hd__buf_1 _40619_ (.A(_09849_),
    .X(_10085_));
 sky130_fd_sc_hd__nand4_4 _40620_ (.A(_10084_),
    .B(_10085_),
    .C(_08310_),
    .D(_08311_),
    .Y(_10086_));
 sky130_fd_sc_hd__buf_1 _40621_ (.A(_03387_),
    .X(_10087_));
 sky130_fd_sc_hd__nand2_4 _40622_ (.A(_10087_),
    .B(_06086_),
    .Y(_10088_));
 sky130_vsdinv _40623_ (.A(_10088_),
    .Y(_10089_));
 sky130_fd_sc_hd__a21oi_4 _40624_ (.A1(_10082_),
    .A2(_10086_),
    .B1(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__nand3_4 _40625_ (.A(_10082_),
    .B(_10086_),
    .C(_10089_),
    .Y(_10091_));
 sky130_vsdinv _40626_ (.A(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__nor2_4 _40627_ (.A(_10090_),
    .B(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__a21o_4 _40628_ (.A1(_10077_),
    .A2(_10079_),
    .B1(_10093_),
    .X(_10094_));
 sky130_fd_sc_hd__nand3_4 _40629_ (.A(_10077_),
    .B(_10093_),
    .C(_10079_),
    .Y(_10095_));
 sky130_fd_sc_hd__o21ai_4 _40630_ (.A1(_09839_),
    .A2(_09856_),
    .B1(_09841_),
    .Y(_10096_));
 sky130_fd_sc_hd__a21o_4 _40631_ (.A1(_10094_),
    .A2(_10095_),
    .B1(_10096_),
    .X(_10097_));
 sky130_fd_sc_hd__nand3_4 _40632_ (.A(_10096_),
    .B(_10095_),
    .C(_10094_),
    .Y(_10098_));
 sky130_fd_sc_hd__a21boi_4 _40633_ (.A1(_09845_),
    .A2(_09851_),
    .B1_N(_09848_),
    .Y(_10099_));
 sky130_vsdinv _40634_ (.A(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__nand3_4 _40635_ (.A(_10097_),
    .B(_10098_),
    .C(_10100_),
    .Y(_10101_));
 sky130_vsdinv _40636_ (.A(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__nand2_4 _40637_ (.A(_10097_),
    .B(_10098_),
    .Y(_10103_));
 sky130_fd_sc_hd__nand2_4 _40638_ (.A(_10103_),
    .B(_10099_),
    .Y(_10104_));
 sky130_vsdinv _40639_ (.A(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__nand2_4 _40640_ (.A(_09819_),
    .B(_09814_),
    .Y(_10106_));
 sky130_vsdinv _40641_ (.A(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__nand2_4 _40642_ (.A(_08055_),
    .B(_08081_),
    .Y(_10108_));
 sky130_fd_sc_hd__nand2_4 _40643_ (.A(_03353_),
    .B(_06375_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand2_4 _40644_ (.A(_10108_),
    .B(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__nand4_4 _40645_ (.A(_08522_),
    .B(_08752_),
    .C(_03480_),
    .D(_06481_),
    .Y(_10111_));
 sky130_fd_sc_hd__nand2_4 _40646_ (.A(_10110_),
    .B(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__nand2_4 _40647_ (.A(_09086_),
    .B(_03475_),
    .Y(_10113_));
 sky130_fd_sc_hd__nand2_4 _40648_ (.A(_10112_),
    .B(_10113_),
    .Y(_10114_));
 sky130_vsdinv _40649_ (.A(_10113_),
    .Y(_10115_));
 sky130_fd_sc_hd__nand3_4 _40650_ (.A(_10110_),
    .B(_10111_),
    .C(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__nand2_4 _40651_ (.A(_10114_),
    .B(_10116_),
    .Y(_10117_));
 sky130_vsdinv _40652_ (.A(_09694_),
    .Y(_10118_));
 sky130_fd_sc_hd__a21boi_4 _40653_ (.A1(_09697_),
    .A2(_10118_),
    .B1_N(_09698_),
    .Y(_10119_));
 sky130_fd_sc_hd__nand2_4 _40654_ (.A(_10117_),
    .B(_10119_),
    .Y(_10120_));
 sky130_vsdinv _40655_ (.A(_09698_),
    .Y(_10121_));
 sky130_fd_sc_hd__a21o_4 _40656_ (.A1(_09697_),
    .A2(_10118_),
    .B1(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__nand3_4 _40657_ (.A(_10122_),
    .B(_10116_),
    .C(_10114_),
    .Y(_10123_));
 sky130_fd_sc_hd__nand2_4 _40658_ (.A(_10120_),
    .B(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__a21boi_4 _40659_ (.A1(_09791_),
    .A2(_09796_),
    .B1_N(_09792_),
    .Y(_10125_));
 sky130_fd_sc_hd__nand2_4 _40660_ (.A(_10124_),
    .B(_10125_),
    .Y(_10126_));
 sky130_vsdinv _40661_ (.A(_10125_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand3_4 _40662_ (.A(_10120_),
    .B(_10123_),
    .C(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__nand2_4 _40663_ (.A(_10126_),
    .B(_10128_),
    .Y(_10129_));
 sky130_vsdinv _40664_ (.A(_09693_),
    .Y(_10130_));
 sky130_fd_sc_hd__a21oi_4 _40665_ (.A1(_09700_),
    .A2(_09691_),
    .B1(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__nand2_4 _40666_ (.A(_10129_),
    .B(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__a21o_4 _40667_ (.A1(_09700_),
    .A2(_09691_),
    .B1(_10130_),
    .X(_10133_));
 sky130_fd_sc_hd__nand3_4 _40668_ (.A(_10133_),
    .B(_10128_),
    .C(_10126_),
    .Y(_10134_));
 sky130_fd_sc_hd__nand2_4 _40669_ (.A(_10132_),
    .B(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__a21boi_4 _40670_ (.A1(_09800_),
    .A2(_09807_),
    .B1_N(_09803_),
    .Y(_10136_));
 sky130_fd_sc_hd__nand2_4 _40671_ (.A(_10135_),
    .B(_10136_),
    .Y(_10137_));
 sky130_vsdinv _40672_ (.A(_10136_),
    .Y(_10138_));
 sky130_fd_sc_hd__nand3_4 _40673_ (.A(_10132_),
    .B(_10134_),
    .C(_10138_),
    .Y(_10139_));
 sky130_fd_sc_hd__nand2_4 _40674_ (.A(_10137_),
    .B(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__nand2_4 _40675_ (.A(_10107_),
    .B(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__nand3_4 _40676_ (.A(_10106_),
    .B(_10139_),
    .C(_10137_),
    .Y(_10142_));
 sky130_fd_sc_hd__nand2_4 _40677_ (.A(_10141_),
    .B(_10142_),
    .Y(_10143_));
 sky130_fd_sc_hd__o21ai_4 _40678_ (.A1(_10102_),
    .A2(_10105_),
    .B1(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__and2_4 _40679_ (.A(_10104_),
    .B(_10101_),
    .X(_10145_));
 sky130_fd_sc_hd__nand3_4 _40680_ (.A(_10145_),
    .B(_10142_),
    .C(_10141_),
    .Y(_10146_));
 sky130_fd_sc_hd__nand2_4 _40681_ (.A(_10144_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__a21boi_4 _40682_ (.A1(_09709_),
    .A2(_09715_),
    .B1_N(_09711_),
    .Y(_10148_));
 sky130_fd_sc_hd__nand2_4 _40683_ (.A(_10147_),
    .B(_10148_),
    .Y(_10149_));
 sky130_vsdinv _40684_ (.A(_10148_),
    .Y(_10150_));
 sky130_fd_sc_hd__nand3_4 _40685_ (.A(_10150_),
    .B(_10146_),
    .C(_10144_),
    .Y(_10151_));
 sky130_fd_sc_hd__nand2_4 _40686_ (.A(_10149_),
    .B(_10151_),
    .Y(_10152_));
 sky130_fd_sc_hd__a21boi_4 _40687_ (.A1(_09871_),
    .A2(_09821_),
    .B1_N(_09822_),
    .Y(_10153_));
 sky130_fd_sc_hd__nand2_4 _40688_ (.A(_10152_),
    .B(_10153_),
    .Y(_10154_));
 sky130_vsdinv _40689_ (.A(_10153_),
    .Y(_10155_));
 sky130_fd_sc_hd__nand3_4 _40690_ (.A(_10149_),
    .B(_10151_),
    .C(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__nand2_4 _40691_ (.A(_10154_),
    .B(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__nand2_4 _40692_ (.A(_10066_),
    .B(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__nand4_4 _40693_ (.A(_10156_),
    .B(_10062_),
    .C(_10154_),
    .D(_10065_),
    .Y(_10159_));
 sky130_fd_sc_hd__nand2_4 _40694_ (.A(_10158_),
    .B(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand2_4 _40695_ (.A(_09918_),
    .B(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__nand2_4 _40696_ (.A(_09886_),
    .B(_09785_),
    .Y(_10162_));
 sky130_fd_sc_hd__nand3_4 _40697_ (.A(_10162_),
    .B(_10159_),
    .C(_10158_),
    .Y(_10163_));
 sky130_fd_sc_hd__nand2_4 _40698_ (.A(_10161_),
    .B(_10163_),
    .Y(_10164_));
 sky130_fd_sc_hd__a21boi_4 _40699_ (.A1(_09862_),
    .A2(_09864_),
    .B1_N(_09860_),
    .Y(_10165_));
 sky130_fd_sc_hd__a21boi_4 _40700_ (.A1(_09876_),
    .A2(_09882_),
    .B1_N(_09878_),
    .Y(_10166_));
 sky130_fd_sc_hd__xnor2_4 _40701_ (.A(_10165_),
    .B(_10166_),
    .Y(_10167_));
 sky130_fd_sc_hd__nand2_4 _40702_ (.A(_10164_),
    .B(_10167_),
    .Y(_10168_));
 sky130_vsdinv _40703_ (.A(_10167_),
    .Y(_10169_));
 sky130_fd_sc_hd__nand3_4 _40704_ (.A(_10161_),
    .B(_10163_),
    .C(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__nand2_4 _40705_ (.A(_10168_),
    .B(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__a21boi_4 _40706_ (.A1(_09898_),
    .A2(_09890_),
    .B1_N(_09892_),
    .Y(_10172_));
 sky130_fd_sc_hd__nand2_4 _40707_ (.A(_10171_),
    .B(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__nand2_4 _40708_ (.A(_09899_),
    .B(_09892_),
    .Y(_10174_));
 sky130_fd_sc_hd__nand3_4 _40709_ (.A(_10174_),
    .B(_10168_),
    .C(_10170_),
    .Y(_10175_));
 sky130_fd_sc_hd__nand2_4 _40710_ (.A(_10173_),
    .B(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__a21oi_4 _40711_ (.A1(_09614_),
    .A2(_09609_),
    .B1(_09894_),
    .Y(_10177_));
 sky130_vsdinv _40712_ (.A(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand2_4 _40713_ (.A(_10176_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__nand3_4 _40714_ (.A(_10173_),
    .B(_10177_),
    .C(_10175_),
    .Y(_10180_));
 sky130_fd_sc_hd__nand2_4 _40715_ (.A(_10179_),
    .B(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__a21boi_4 _40716_ (.A1(_09902_),
    .A2(_09906_),
    .B1_N(_09904_),
    .Y(_10182_));
 sky130_fd_sc_hd__nand2_4 _40717_ (.A(_10181_),
    .B(_10182_),
    .Y(_10183_));
 sky130_vsdinv _40718_ (.A(_10182_),
    .Y(_10184_));
 sky130_fd_sc_hd__nand3_4 _40719_ (.A(_10184_),
    .B(_10180_),
    .C(_10179_),
    .Y(_10185_));
 sky130_fd_sc_hd__and2_4 _40720_ (.A(_10183_),
    .B(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__buf_1 _40721_ (.A(_10186_),
    .X(_10187_));
 sky130_fd_sc_hd__nand4_4 _40722_ (.A(_09643_),
    .B(_09641_),
    .C(_09912_),
    .D(_09914_),
    .Y(_10188_));
 sky130_vsdinv _40723_ (.A(_09643_),
    .Y(_10189_));
 sky130_fd_sc_hd__a21boi_4 _40724_ (.A1(_10189_),
    .A2(_09912_),
    .B1_N(_09914_),
    .Y(_10190_));
 sky130_fd_sc_hd__o21ai_4 _40725_ (.A1(_09651_),
    .A2(_10188_),
    .B1(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__a41o_4 _40726_ (.A1(_09647_),
    .A2(_09645_),
    .A3(_09648_),
    .A4(_09916_),
    .B1(_10191_),
    .X(_10192_));
 sky130_fd_sc_hd__xor2_4 _40727_ (.A(_10187_),
    .B(_10192_),
    .X(_01433_));
 sky130_fd_sc_hd__maj3_4 _40728_ (.A(_09949_),
    .B(_09945_),
    .C(_09946_),
    .X(_10193_));
 sky130_vsdinv _40729_ (.A(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__nand2_4 _40730_ (.A(_08966_),
    .B(_07353_),
    .Y(_10195_));
 sky130_fd_sc_hd__nand2_4 _40731_ (.A(_09037_),
    .B(_07521_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand2_4 _40732_ (.A(_10195_),
    .B(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__buf_1 _40733_ (.A(_03317_),
    .X(_10198_));
 sky130_fd_sc_hd__nand4_4 _40734_ (.A(_10198_),
    .B(_07624_),
    .C(_07940_),
    .D(_07941_),
    .Y(_10199_));
 sky130_fd_sc_hd__nand2_4 _40735_ (.A(_03332_),
    .B(_08383_),
    .Y(_10200_));
 sky130_vsdinv _40736_ (.A(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand3_4 _40737_ (.A(_10197_),
    .B(_10199_),
    .C(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__a21o_4 _40738_ (.A1(_10197_),
    .A2(_10199_),
    .B1(_10201_),
    .X(_10203_));
 sky130_fd_sc_hd__nand3_4 _40739_ (.A(_10194_),
    .B(_10202_),
    .C(_10203_),
    .Y(_10204_));
 sky130_fd_sc_hd__nand2_4 _40740_ (.A(_10203_),
    .B(_10202_),
    .Y(_10205_));
 sky130_fd_sc_hd__nand2_4 _40741_ (.A(_10205_),
    .B(_10193_),
    .Y(_10206_));
 sky130_fd_sc_hd__nand2_4 _40742_ (.A(_10204_),
    .B(_10206_),
    .Y(_10207_));
 sky130_fd_sc_hd__nand2_4 _40743_ (.A(_08522_),
    .B(_03495_),
    .Y(_10208_));
 sky130_fd_sc_hd__nand2_4 _40744_ (.A(_08042_),
    .B(_07214_),
    .Y(_10209_));
 sky130_fd_sc_hd__nand2_4 _40745_ (.A(_09070_),
    .B(_07212_),
    .Y(_10210_));
 sky130_fd_sc_hd__nand2_4 _40746_ (.A(_10209_),
    .B(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__buf_1 _40747_ (.A(_07870_),
    .X(_10212_));
 sky130_fd_sc_hd__nand4_4 _40748_ (.A(_10212_),
    .B(_07878_),
    .C(_07956_),
    .D(_06893_),
    .Y(_10213_));
 sky130_fd_sc_hd__nand2_4 _40749_ (.A(_10211_),
    .B(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__xor2_4 _40750_ (.A(_10208_),
    .B(_10214_),
    .X(_10215_));
 sky130_vsdinv _40751_ (.A(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__nand2_4 _40752_ (.A(_10207_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__nand3_4 _40753_ (.A(_10204_),
    .B(_10215_),
    .C(_10206_),
    .Y(_10218_));
 sky130_fd_sc_hd__and2_4 _40754_ (.A(_10217_),
    .B(_10218_),
    .X(_10219_));
 sky130_vsdinv _40755_ (.A(_10219_),
    .Y(_10220_));
 sky130_fd_sc_hd__a21boi_4 _40756_ (.A1(_10002_),
    .A2(_09999_),
    .B1_N(_10003_),
    .Y(_10221_));
 sky130_vsdinv _40757_ (.A(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__nand2_4 _40758_ (.A(_06711_),
    .B(_03540_),
    .Y(_10223_));
 sky130_fd_sc_hd__nand2_4 _40759_ (.A(_06851_),
    .B(_08795_),
    .Y(_10224_));
 sky130_fd_sc_hd__nand2_4 _40760_ (.A(_10223_),
    .B(_10224_),
    .Y(_10225_));
 sky130_fd_sc_hd__nand4_4 _40761_ (.A(_03303_),
    .B(_07146_),
    .C(_07553_),
    .D(_07556_),
    .Y(_10226_));
 sky130_fd_sc_hd__nand2_4 _40762_ (.A(_06991_),
    .B(_07719_),
    .Y(_10227_));
 sky130_vsdinv _40763_ (.A(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__nand3_4 _40764_ (.A(_10225_),
    .B(_10226_),
    .C(_10228_),
    .Y(_10229_));
 sky130_fd_sc_hd__nand2_4 _40765_ (.A(_10225_),
    .B(_10226_),
    .Y(_10230_));
 sky130_fd_sc_hd__nand2_4 _40766_ (.A(_10230_),
    .B(_10227_),
    .Y(_10231_));
 sky130_fd_sc_hd__nand3_4 _40767_ (.A(_10222_),
    .B(_10229_),
    .C(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__nand2_4 _40768_ (.A(_10231_),
    .B(_10229_),
    .Y(_10233_));
 sky130_fd_sc_hd__nand2_4 _40769_ (.A(_10233_),
    .B(_10221_),
    .Y(_10234_));
 sky130_fd_sc_hd__nand2_4 _40770_ (.A(_10232_),
    .B(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__a21boi_4 _40771_ (.A1(_09921_),
    .A2(_09926_),
    .B1_N(_09922_),
    .Y(_10236_));
 sky130_fd_sc_hd__nand2_4 _40772_ (.A(_10235_),
    .B(_10236_),
    .Y(_10237_));
 sky130_vsdinv _40773_ (.A(_10236_),
    .Y(_10238_));
 sky130_fd_sc_hd__nand3_4 _40774_ (.A(_10232_),
    .B(_10234_),
    .C(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__nand2_4 _40775_ (.A(_10237_),
    .B(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__a21boi_4 _40776_ (.A1(_09930_),
    .A2(_09937_),
    .B1_N(_09933_),
    .Y(_10241_));
 sky130_fd_sc_hd__nand2_4 _40777_ (.A(_10240_),
    .B(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__nand2_4 _40778_ (.A(_09938_),
    .B(_09933_),
    .Y(_10243_));
 sky130_fd_sc_hd__nand3_4 _40779_ (.A(_10243_),
    .B(_10237_),
    .C(_10239_),
    .Y(_10244_));
 sky130_fd_sc_hd__nand2_4 _40780_ (.A(_10242_),
    .B(_10244_),
    .Y(_10245_));
 sky130_fd_sc_hd__nand2_4 _40781_ (.A(_10220_),
    .B(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__nand3_4 _40782_ (.A(_10219_),
    .B(_10244_),
    .C(_10242_),
    .Y(_10247_));
 sky130_fd_sc_hd__nand2_4 _40783_ (.A(_10246_),
    .B(_10247_),
    .Y(_10248_));
 sky130_vsdinv _40784_ (.A(_10012_),
    .Y(_10249_));
 sky130_fd_sc_hd__a21oi_4 _40785_ (.A1(_10010_),
    .A2(_10016_),
    .B1(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__nand2_4 _40786_ (.A(_10248_),
    .B(_10250_),
    .Y(_10251_));
 sky130_vsdinv _40787_ (.A(_10250_),
    .Y(_10252_));
 sky130_fd_sc_hd__nand3_4 _40788_ (.A(_10252_),
    .B(_10247_),
    .C(_10246_),
    .Y(_10253_));
 sky130_fd_sc_hd__nand2_4 _40789_ (.A(_10251_),
    .B(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__a21boi_4 _40790_ (.A1(_09941_),
    .A2(_09967_),
    .B1_N(_09943_),
    .Y(_10255_));
 sky130_fd_sc_hd__nand2_4 _40791_ (.A(_10254_),
    .B(_10255_),
    .Y(_10256_));
 sky130_vsdinv _40792_ (.A(_10255_),
    .Y(_10257_));
 sky130_fd_sc_hd__nand3_4 _40793_ (.A(_10251_),
    .B(_10253_),
    .C(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__nand2_4 _40794_ (.A(_10256_),
    .B(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__nand2_4 _40795_ (.A(_03298_),
    .B(_03544_),
    .Y(_10260_));
 sky130_fd_sc_hd__nand2_4 _40796_ (.A(_07753_),
    .B(_09486_),
    .Y(_10261_));
 sky130_fd_sc_hd__buf_1 _40797_ (.A(_03551_),
    .X(_10262_));
 sky130_fd_sc_hd__nand2_4 _40798_ (.A(_06455_),
    .B(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__nand2_4 _40799_ (.A(_10261_),
    .B(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__buf_1 _40800_ (.A(_03290_),
    .X(_10265_));
 sky130_fd_sc_hd__nand4_4 _40801_ (.A(_10265_),
    .B(_07952_),
    .C(_09416_),
    .D(_09415_),
    .Y(_10266_));
 sky130_fd_sc_hd__nand2_4 _40802_ (.A(_10264_),
    .B(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__xor2_4 _40803_ (.A(_10260_),
    .B(_10267_),
    .X(_10268_));
 sky130_vsdinv _40804_ (.A(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__buf_1 _40805_ (.A(_03574_),
    .X(_10270_));
 sky130_fd_sc_hd__nand2_4 _40806_ (.A(_06169_),
    .B(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__buf_1 _40807_ (.A(_08629_),
    .X(_10272_));
 sky130_fd_sc_hd__nand2_4 _40808_ (.A(_06339_),
    .B(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__nand2_4 _40809_ (.A(_10271_),
    .B(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__buf_1 _40810_ (.A(_09467_),
    .X(_10275_));
 sky130_fd_sc_hd__nand4_4 _40811_ (.A(_06325_),
    .B(_03275_),
    .C(_10272_),
    .D(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__nand2_4 _40812_ (.A(_10274_),
    .B(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__nand2_4 _40813_ (.A(_07761_),
    .B(_03563_),
    .Y(_10278_));
 sky130_fd_sc_hd__nand2_4 _40814_ (.A(_10277_),
    .B(_10278_),
    .Y(_10279_));
 sky130_vsdinv _40815_ (.A(_10278_),
    .Y(_10280_));
 sky130_fd_sc_hd__nand3_4 _40816_ (.A(_10274_),
    .B(_10276_),
    .C(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__nand2_4 _40817_ (.A(_10279_),
    .B(_10281_),
    .Y(_10282_));
 sky130_fd_sc_hd__a21boi_4 _40818_ (.A1(_09985_),
    .A2(_09990_),
    .B1_N(_09986_),
    .Y(_10283_));
 sky130_fd_sc_hd__nand2_4 _40819_ (.A(_10282_),
    .B(_10283_),
    .Y(_10284_));
 sky130_fd_sc_hd__nand2_4 _40820_ (.A(_09991_),
    .B(_09986_),
    .Y(_10285_));
 sky130_fd_sc_hd__nand3_4 _40821_ (.A(_10285_),
    .B(_10281_),
    .C(_10279_),
    .Y(_10286_));
 sky130_fd_sc_hd__nand2_4 _40822_ (.A(_10284_),
    .B(_10286_),
    .Y(_10287_));
 sky130_fd_sc_hd__nand2_4 _40823_ (.A(_10269_),
    .B(_10287_),
    .Y(_10288_));
 sky130_fd_sc_hd__nand3_4 _40824_ (.A(_10268_),
    .B(_10284_),
    .C(_10286_),
    .Y(_10289_));
 sky130_fd_sc_hd__nand2_4 _40825_ (.A(_10288_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__nand2_4 _40826_ (.A(_10290_),
    .B(_10032_),
    .Y(_10291_));
 sky130_vsdinv _40827_ (.A(_10032_),
    .Y(_10292_));
 sky130_fd_sc_hd__nand3_4 _40828_ (.A(_10288_),
    .B(_10292_),
    .C(_10289_),
    .Y(_10293_));
 sky130_fd_sc_hd__nand2_4 _40829_ (.A(_10291_),
    .B(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__a21boi_4 _40830_ (.A1(_10007_),
    .A2(_09994_),
    .B1_N(_09996_),
    .Y(_10295_));
 sky130_fd_sc_hd__nand2_4 _40831_ (.A(_10294_),
    .B(_10295_),
    .Y(_10296_));
 sky130_vsdinv _40832_ (.A(_10295_),
    .Y(_10297_));
 sky130_fd_sc_hd__nand3_4 _40833_ (.A(_10291_),
    .B(_10297_),
    .C(_10293_),
    .Y(_10298_));
 sky130_fd_sc_hd__nand2_4 _40834_ (.A(_10296_),
    .B(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__buf_1 _40835_ (.A(_09500_),
    .X(_10300_));
 sky130_fd_sc_hd__nand2_4 _40836_ (.A(_05915_),
    .B(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__buf_1 _40837_ (.A(_09342_),
    .X(_10302_));
 sky130_fd_sc_hd__nand2_4 _40838_ (.A(_07365_),
    .B(_10302_),
    .Y(_10303_));
 sky130_fd_sc_hd__nand2_4 _40839_ (.A(_10301_),
    .B(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__buf_1 _40840_ (.A(_09500_),
    .X(_10305_));
 sky130_fd_sc_hd__nand4_4 _40841_ (.A(_06384_),
    .B(_06010_),
    .C(_03587_),
    .D(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__nand2_4 _40842_ (.A(_10304_),
    .B(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__nand2_4 _40843_ (.A(_06019_),
    .B(_03581_),
    .Y(_10308_));
 sky130_fd_sc_hd__nand2_4 _40844_ (.A(_10307_),
    .B(_10308_),
    .Y(_10309_));
 sky130_vsdinv _40845_ (.A(_10308_),
    .Y(_10310_));
 sky130_fd_sc_hd__nand3_4 _40846_ (.A(_10304_),
    .B(_10306_),
    .C(_10310_),
    .Y(_10311_));
 sky130_fd_sc_hd__nand2_4 _40847_ (.A(_10309_),
    .B(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__nand2_4 _40848_ (.A(_10312_),
    .B(_10038_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand3_4 _40849_ (.A(_10309_),
    .B(_10037_),
    .C(_10311_),
    .Y(_10314_));
 sky130_fd_sc_hd__nand2_4 _40850_ (.A(_10313_),
    .B(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__a21boi_4 _40851_ (.A1(_10021_),
    .A2(_10026_),
    .B1_N(_10022_),
    .Y(_10316_));
 sky130_fd_sc_hd__nand2_4 _40852_ (.A(_10315_),
    .B(_10316_),
    .Y(_10317_));
 sky130_vsdinv _40853_ (.A(_10316_),
    .Y(_10318_));
 sky130_fd_sc_hd__nand3_4 _40854_ (.A(_10313_),
    .B(_10318_),
    .C(_10314_),
    .Y(_10319_));
 sky130_fd_sc_hd__nand2_4 _40855_ (.A(_10317_),
    .B(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__nand2_4 _40856_ (.A(_07359_),
    .B(_03600_),
    .Y(_10321_));
 sky130_fd_sc_hd__buf_1 _40857_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10322_));
 sky130_fd_sc_hd__nand2_4 _40858_ (.A(_06370_),
    .B(_10322_),
    .Y(_10323_));
 sky130_fd_sc_hd__buf_1 _40859_ (.A(\pcpi_mul.rs2[29] ),
    .X(_10324_));
 sky130_fd_sc_hd__nand2_4 _40860_ (.A(_03228_),
    .B(_10324_),
    .Y(_10325_));
 sky130_fd_sc_hd__nand2_4 _40861_ (.A(_10323_),
    .B(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__nand4_4 _40862_ (.A(_03228_),
    .B(_06370_),
    .C(_10322_),
    .D(_10324_),
    .Y(_10327_));
 sky130_fd_sc_hd__nand2_4 _40863_ (.A(_10326_),
    .B(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__xor2_4 _40864_ (.A(_10321_),
    .B(_10328_),
    .X(_10329_));
 sky130_vsdinv _40865_ (.A(_10329_),
    .Y(_10330_));
 sky130_fd_sc_hd__nand2_4 _40866_ (.A(_10320_),
    .B(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__nand3_4 _40867_ (.A(_10317_),
    .B(_10329_),
    .C(_10319_),
    .Y(_10332_));
 sky130_fd_sc_hd__nand2_4 _40868_ (.A(_10331_),
    .B(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__nand2_4 _40869_ (.A(_10333_),
    .B(_10043_),
    .Y(_10334_));
 sky130_vsdinv _40870_ (.A(_10043_),
    .Y(_10335_));
 sky130_fd_sc_hd__nand3_4 _40871_ (.A(_10331_),
    .B(_10335_),
    .C(_10332_),
    .Y(_10336_));
 sky130_fd_sc_hd__nand2_4 _40872_ (.A(_10334_),
    .B(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__nand2_4 _40873_ (.A(_10299_),
    .B(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__nand4_4 _40874_ (.A(_10298_),
    .B(_10296_),
    .C(_10334_),
    .D(_10336_),
    .Y(_10339_));
 sky130_fd_sc_hd__nand2_4 _40875_ (.A(_10338_),
    .B(_10339_),
    .Y(_10340_));
 sky130_fd_sc_hd__nand2_4 _40876_ (.A(_10053_),
    .B(_10049_),
    .Y(_10341_));
 sky130_vsdinv _40877_ (.A(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__nand2_4 _40878_ (.A(_10340_),
    .B(_10342_),
    .Y(_10343_));
 sky130_fd_sc_hd__nand3_4 _40879_ (.A(_10341_),
    .B(_10338_),
    .C(_10339_),
    .Y(_10344_));
 sky130_fd_sc_hd__nand2_4 _40880_ (.A(_10343_),
    .B(_10344_),
    .Y(_10345_));
 sky130_fd_sc_hd__nand2_4 _40881_ (.A(_10259_),
    .B(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__nand4_4 _40882_ (.A(_10258_),
    .B(_10256_),
    .C(_10343_),
    .D(_10344_),
    .Y(_10347_));
 sky130_fd_sc_hd__nand2_4 _40883_ (.A(_10346_),
    .B(_10347_),
    .Y(_10348_));
 sky130_fd_sc_hd__nand3_4 _40884_ (.A(_10348_),
    .B(_10057_),
    .C(_10064_),
    .Y(_10349_));
 sky130_fd_sc_hd__nand2_4 _40885_ (.A(_10064_),
    .B(_10057_),
    .Y(_10350_));
 sky130_fd_sc_hd__nand3_4 _40886_ (.A(_10350_),
    .B(_10347_),
    .C(_10346_),
    .Y(_10351_));
 sky130_fd_sc_hd__nand2_4 _40887_ (.A(_10349_),
    .B(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__nand2_4 _40888_ (.A(_09965_),
    .B(_09956_),
    .Y(_10353_));
 sky130_vsdinv _40889_ (.A(_09957_),
    .Y(_10354_));
 sky130_fd_sc_hd__a21boi_4 _40890_ (.A1(_09960_),
    .A2(_10354_),
    .B1_N(_09961_),
    .Y(_10355_));
 sky130_vsdinv _40891_ (.A(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__nand2_4 _40892_ (.A(_08752_),
    .B(_06593_),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_4 _40893_ (.A(_08530_),
    .B(_06599_),
    .Y(_10358_));
 sky130_fd_sc_hd__nand2_4 _40894_ (.A(_10357_),
    .B(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__nand4_4 _40895_ (.A(_08527_),
    .B(_03357_),
    .C(_06946_),
    .D(_06788_),
    .Y(_10360_));
 sky130_fd_sc_hd__nand2_4 _40896_ (.A(_10359_),
    .B(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__nand2_4 _40897_ (.A(_03361_),
    .B(_06796_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand2_4 _40898_ (.A(_10361_),
    .B(_10362_),
    .Y(_10363_));
 sky130_vsdinv _40899_ (.A(_10362_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand3_4 _40900_ (.A(_10359_),
    .B(_10360_),
    .C(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__nand3_4 _40901_ (.A(_10356_),
    .B(_10363_),
    .C(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__nand2_4 _40902_ (.A(_10363_),
    .B(_10365_),
    .Y(_10367_));
 sky130_fd_sc_hd__nand2_4 _40903_ (.A(_10367_),
    .B(_10355_),
    .Y(_10368_));
 sky130_fd_sc_hd__a21boi_4 _40904_ (.A1(_10110_),
    .A2(_10115_),
    .B1_N(_10111_),
    .Y(_10369_));
 sky130_vsdinv _40905_ (.A(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__nand3_4 _40906_ (.A(_10366_),
    .B(_10368_),
    .C(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__nand2_4 _40907_ (.A(_10366_),
    .B(_10368_),
    .Y(_10372_));
 sky130_fd_sc_hd__nand2_4 _40908_ (.A(_10372_),
    .B(_10369_),
    .Y(_10373_));
 sky130_fd_sc_hd__nand3_4 _40909_ (.A(_10353_),
    .B(_10371_),
    .C(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__nand2_4 _40910_ (.A(_10373_),
    .B(_10371_),
    .Y(_10375_));
 sky130_fd_sc_hd__a21boi_4 _40911_ (.A1(_09954_),
    .A2(_09963_),
    .B1_N(_09956_),
    .Y(_10376_));
 sky130_fd_sc_hd__nand2_4 _40912_ (.A(_10375_),
    .B(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__nand2_4 _40913_ (.A(_10374_),
    .B(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__a21boi_4 _40914_ (.A1(_10120_),
    .A2(_10127_),
    .B1_N(_10123_),
    .Y(_10379_));
 sky130_fd_sc_hd__nand2_4 _40915_ (.A(_10378_),
    .B(_10379_),
    .Y(_10380_));
 sky130_vsdinv _40916_ (.A(_10379_),
    .Y(_10381_));
 sky130_fd_sc_hd__nand3_4 _40917_ (.A(_10374_),
    .B(_10377_),
    .C(_10381_),
    .Y(_10382_));
 sky130_fd_sc_hd__nand2_4 _40918_ (.A(_10380_),
    .B(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__a21boi_4 _40919_ (.A1(_10132_),
    .A2(_10138_),
    .B1_N(_10134_),
    .Y(_10384_));
 sky130_fd_sc_hd__nand2_4 _40920_ (.A(_10383_),
    .B(_10384_),
    .Y(_10385_));
 sky130_vsdinv _40921_ (.A(_10384_),
    .Y(_10386_));
 sky130_fd_sc_hd__nand3_4 _40922_ (.A(_10386_),
    .B(_10382_),
    .C(_10380_),
    .Y(_10387_));
 sky130_fd_sc_hd__nand2_4 _40923_ (.A(_10385_),
    .B(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__nand2_4 _40924_ (.A(_09212_),
    .B(_06052_),
    .Y(_10389_));
 sky130_fd_sc_hd__nand2_4 _40925_ (.A(_09843_),
    .B(_08734_),
    .Y(_10390_));
 sky130_fd_sc_hd__nand2_4 _40926_ (.A(_10389_),
    .B(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__nand4_4 _40927_ (.A(_09833_),
    .B(_09843_),
    .C(_08028_),
    .D(_06322_),
    .Y(_10392_));
 sky130_fd_sc_hd__buf_1 _40928_ (.A(\pcpi_mul.rs1[26] ),
    .X(_10393_));
 sky130_fd_sc_hd__nand2_4 _40929_ (.A(_10393_),
    .B(_03453_),
    .Y(_10394_));
 sky130_vsdinv _40930_ (.A(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__a21o_4 _40931_ (.A1(_10391_),
    .A2(_10392_),
    .B1(_10395_),
    .X(_10396_));
 sky130_fd_sc_hd__nand3_4 _40932_ (.A(_10391_),
    .B(_10392_),
    .C(_10395_),
    .Y(_10397_));
 sky130_fd_sc_hd__a21boi_4 _40933_ (.A1(_10069_),
    .A2(_10072_),
    .B1_N(_10070_),
    .Y(_10398_));
 sky130_fd_sc_hd__a21boi_4 _40934_ (.A1(_10396_),
    .A2(_10397_),
    .B1_N(_10398_),
    .Y(_10399_));
 sky130_vsdinv _40935_ (.A(_10399_),
    .Y(_10400_));
 sky130_vsdinv _40936_ (.A(_10398_),
    .Y(_10401_));
 sky130_fd_sc_hd__nand3_4 _40937_ (.A(_10401_),
    .B(_10396_),
    .C(_10397_),
    .Y(_10402_));
 sky130_fd_sc_hd__nand2_4 _40938_ (.A(_03382_),
    .B(_05909_),
    .Y(_10403_));
 sky130_fd_sc_hd__o21ai_4 _40939_ (.A1(_03388_),
    .A2(_07618_),
    .B1(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__buf_1 _40940_ (.A(\pcpi_mul.rs1[27] ),
    .X(_10405_));
 sky130_fd_sc_hd__buf_1 _40941_ (.A(\pcpi_mul.rs1[28] ),
    .X(_10406_));
 sky130_fd_sc_hd__nand4_4 _40942_ (.A(_10405_),
    .B(_10406_),
    .C(_07001_),
    .D(_06015_),
    .Y(_10407_));
 sky130_fd_sc_hd__buf_1 _40943_ (.A(\pcpi_mul.rs1[29] ),
    .X(_10408_));
 sky130_fd_sc_hd__buf_1 _40944_ (.A(_10408_),
    .X(_10409_));
 sky130_fd_sc_hd__nand2_4 _40945_ (.A(_10409_),
    .B(_06853_),
    .Y(_10410_));
 sky130_vsdinv _40946_ (.A(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__a21o_4 _40947_ (.A1(_10404_),
    .A2(_10407_),
    .B1(_10411_),
    .X(_10412_));
 sky130_fd_sc_hd__nand3_4 _40948_ (.A(_10404_),
    .B(_10407_),
    .C(_10411_),
    .Y(_10413_));
 sky130_fd_sc_hd__and2_4 _40949_ (.A(_10412_),
    .B(_10413_),
    .X(_10414_));
 sky130_fd_sc_hd__buf_1 _40950_ (.A(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__a21o_4 _40951_ (.A1(_10400_),
    .A2(_10402_),
    .B1(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__nand3_4 _40952_ (.A(_10400_),
    .B(_10415_),
    .C(_10402_),
    .Y(_10417_));
 sky130_fd_sc_hd__a21boi_4 _40953_ (.A1(_10077_),
    .A2(_10093_),
    .B1_N(_10079_),
    .Y(_10418_));
 sky130_vsdinv _40954_ (.A(_10418_),
    .Y(_10419_));
 sky130_fd_sc_hd__a21oi_4 _40955_ (.A1(_10416_),
    .A2(_10417_),
    .B1(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__nand3_4 _40956_ (.A(_10416_),
    .B(_10419_),
    .C(_10417_),
    .Y(_10421_));
 sky130_vsdinv _40957_ (.A(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__a21boi_4 _40958_ (.A1(_10082_),
    .A2(_10089_),
    .B1_N(_10086_),
    .Y(_10423_));
 sky130_fd_sc_hd__o21ai_4 _40959_ (.A1(_10420_),
    .A2(_10422_),
    .B1(_10423_),
    .Y(_10424_));
 sky130_vsdinv _40960_ (.A(_10420_),
    .Y(_10425_));
 sky130_vsdinv _40961_ (.A(_10423_),
    .Y(_10426_));
 sky130_fd_sc_hd__nand3_4 _40962_ (.A(_10425_),
    .B(_10426_),
    .C(_10421_),
    .Y(_10427_));
 sky130_fd_sc_hd__nand2_4 _40963_ (.A(_10424_),
    .B(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__nand2_4 _40964_ (.A(_10388_),
    .B(_10428_),
    .Y(_10429_));
 sky130_fd_sc_hd__nand4_4 _40965_ (.A(_10427_),
    .B(_10385_),
    .C(_10387_),
    .D(_10424_),
    .Y(_10430_));
 sky130_fd_sc_hd__nand2_4 _40966_ (.A(_10429_),
    .B(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__a21boi_4 _40967_ (.A1(_09974_),
    .A2(_09980_),
    .B1_N(_09976_),
    .Y(_10432_));
 sky130_fd_sc_hd__nand2_4 _40968_ (.A(_10431_),
    .B(_10432_),
    .Y(_10433_));
 sky130_vsdinv _40969_ (.A(_10432_),
    .Y(_10434_));
 sky130_fd_sc_hd__nand3_4 _40970_ (.A(_10434_),
    .B(_10430_),
    .C(_10429_),
    .Y(_10435_));
 sky130_fd_sc_hd__nand2_4 _40971_ (.A(_10433_),
    .B(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__a21boi_4 _40972_ (.A1(_10145_),
    .A2(_10141_),
    .B1_N(_10142_),
    .Y(_10437_));
 sky130_fd_sc_hd__nand2_4 _40973_ (.A(_10436_),
    .B(_10437_),
    .Y(_10438_));
 sky130_vsdinv _40974_ (.A(_10437_),
    .Y(_10439_));
 sky130_fd_sc_hd__nand3_4 _40975_ (.A(_10433_),
    .B(_10435_),
    .C(_10439_),
    .Y(_10440_));
 sky130_fd_sc_hd__nand2_4 _40976_ (.A(_10438_),
    .B(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__nand2_4 _40977_ (.A(_10352_),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__nand4_4 _40978_ (.A(_10440_),
    .B(_10349_),
    .C(_10438_),
    .D(_10351_),
    .Y(_10443_));
 sky130_fd_sc_hd__nand2_4 _40979_ (.A(_10442_),
    .B(_10443_),
    .Y(_10444_));
 sky130_fd_sc_hd__a21oi_4 _40980_ (.A1(_10064_),
    .A2(_10059_),
    .B1(_10063_),
    .Y(_10445_));
 sky130_fd_sc_hd__o21a_4 _40981_ (.A1(_10445_),
    .A2(_10157_),
    .B1(_10065_),
    .X(_10446_));
 sky130_fd_sc_hd__nand2_4 _40982_ (.A(_10444_),
    .B(_10446_),
    .Y(_10447_));
 sky130_fd_sc_hd__o21ai_4 _40983_ (.A1(_10445_),
    .A2(_10157_),
    .B1(_10065_),
    .Y(_10448_));
 sky130_fd_sc_hd__nand3_4 _40984_ (.A(_10448_),
    .B(_10443_),
    .C(_10442_),
    .Y(_10449_));
 sky130_fd_sc_hd__nand2_4 _40985_ (.A(_10447_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__a21boi_4 _40986_ (.A1(_10097_),
    .A2(_10100_),
    .B1_N(_10098_),
    .Y(_10451_));
 sky130_fd_sc_hd__a21boi_4 _40987_ (.A1(_10149_),
    .A2(_10155_),
    .B1_N(_10151_),
    .Y(_10452_));
 sky130_fd_sc_hd__xnor2_4 _40988_ (.A(_10451_),
    .B(_10452_),
    .Y(_10453_));
 sky130_fd_sc_hd__nand2_4 _40989_ (.A(_10450_),
    .B(_10453_),
    .Y(_10454_));
 sky130_vsdinv _40990_ (.A(_10453_),
    .Y(_10455_));
 sky130_fd_sc_hd__nand3_4 _40991_ (.A(_10447_),
    .B(_10449_),
    .C(_10455_),
    .Y(_10456_));
 sky130_fd_sc_hd__nand2_4 _40992_ (.A(_10454_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__a21boi_4 _40993_ (.A1(_10161_),
    .A2(_10169_),
    .B1_N(_10163_),
    .Y(_10458_));
 sky130_fd_sc_hd__nand2_4 _40994_ (.A(_10457_),
    .B(_10458_),
    .Y(_10459_));
 sky130_fd_sc_hd__nand2_4 _40995_ (.A(_10170_),
    .B(_10163_),
    .Y(_10460_));
 sky130_fd_sc_hd__nand3_4 _40996_ (.A(_10460_),
    .B(_10454_),
    .C(_10456_),
    .Y(_10461_));
 sky130_fd_sc_hd__nand2_4 _40997_ (.A(_10459_),
    .B(_10461_),
    .Y(_10462_));
 sky130_fd_sc_hd__a21oi_4 _40998_ (.A1(_09883_),
    .A2(_09878_),
    .B1(_10165_),
    .Y(_10463_));
 sky130_vsdinv _40999_ (.A(_10463_),
    .Y(_10464_));
 sky130_fd_sc_hd__nand2_4 _41000_ (.A(_10462_),
    .B(_10464_),
    .Y(_10465_));
 sky130_fd_sc_hd__nand3_4 _41001_ (.A(_10459_),
    .B(_10461_),
    .C(_10463_),
    .Y(_10466_));
 sky130_fd_sc_hd__nand2_4 _41002_ (.A(_10465_),
    .B(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__nand2_4 _41003_ (.A(_10180_),
    .B(_10175_),
    .Y(_10468_));
 sky130_vsdinv _41004_ (.A(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__nand2_4 _41005_ (.A(_10467_),
    .B(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__nand3_4 _41006_ (.A(_10468_),
    .B(_10465_),
    .C(_10466_),
    .Y(_10471_));
 sky130_fd_sc_hd__and2_4 _41007_ (.A(_10470_),
    .B(_10471_),
    .X(_10472_));
 sky130_fd_sc_hd__buf_1 _41008_ (.A(_10472_),
    .X(_10473_));
 sky130_fd_sc_hd__a21boi_4 _41009_ (.A1(_10192_),
    .A2(_10183_),
    .B1_N(_10185_),
    .Y(_10474_));
 sky130_fd_sc_hd__xnor2_4 _41010_ (.A(_10473_),
    .B(_10474_),
    .Y(_01434_));
 sky130_fd_sc_hd__o21a_4 _41011_ (.A1(_10441_),
    .A2(_10352_),
    .B1(_10351_),
    .X(_10475_));
 sky130_fd_sc_hd__buf_1 _41012_ (.A(\pcpi_mul.rs2[26] ),
    .X(_10476_));
 sky130_fd_sc_hd__nand2_4 _41013_ (.A(_07365_),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__nand2_4 _41014_ (.A(_06019_),
    .B(_10302_),
    .Y(_10478_));
 sky130_fd_sc_hd__nand2_4 _41015_ (.A(_10477_),
    .B(_10478_),
    .Y(_10479_));
 sky130_fd_sc_hd__buf_1 _41016_ (.A(_03261_),
    .X(_10480_));
 sky130_fd_sc_hd__buf_1 _41017_ (.A(_09342_),
    .X(_10481_));
 sky130_fd_sc_hd__nand4_4 _41018_ (.A(_10480_),
    .B(_08565_),
    .C(_10481_),
    .D(_10305_),
    .Y(_10482_));
 sky130_fd_sc_hd__nand2_4 _41019_ (.A(_06244_),
    .B(_03581_),
    .Y(_10483_));
 sky130_vsdinv _41020_ (.A(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__a21o_4 _41021_ (.A1(_10479_),
    .A2(_10482_),
    .B1(_10484_),
    .X(_10485_));
 sky130_fd_sc_hd__nand3_4 _41022_ (.A(_10479_),
    .B(_10482_),
    .C(_10484_),
    .Y(_10486_));
 sky130_fd_sc_hd__nand2_4 _41023_ (.A(_10485_),
    .B(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__maj3_4 _41024_ (.A(_10321_),
    .B(_10323_),
    .C(_10325_),
    .X(_10488_));
 sky130_fd_sc_hd__nand2_4 _41025_ (.A(_10487_),
    .B(_10488_),
    .Y(_10489_));
 sky130_fd_sc_hd__o21ai_4 _41026_ (.A1(_10321_),
    .A2(_10328_),
    .B1(_10327_),
    .Y(_10490_));
 sky130_fd_sc_hd__nand3_4 _41027_ (.A(_10490_),
    .B(_10486_),
    .C(_10485_),
    .Y(_10491_));
 sky130_fd_sc_hd__nand2_4 _41028_ (.A(_10489_),
    .B(_10491_),
    .Y(_10492_));
 sky130_fd_sc_hd__a21boi_4 _41029_ (.A1(_10304_),
    .A2(_10310_),
    .B1_N(_10306_),
    .Y(_10493_));
 sky130_fd_sc_hd__nand2_4 _41030_ (.A(_10492_),
    .B(_10493_),
    .Y(_10494_));
 sky130_vsdinv _41031_ (.A(_10493_),
    .Y(_10495_));
 sky130_fd_sc_hd__nand3_4 _41032_ (.A(_10489_),
    .B(_10491_),
    .C(_10495_),
    .Y(_10496_));
 sky130_fd_sc_hd__nand2_4 _41033_ (.A(_10494_),
    .B(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__buf_1 _41034_ (.A(\pcpi_mul.rs2[29] ),
    .X(_10498_));
 sky130_fd_sc_hd__buf_1 _41035_ (.A(_10498_),
    .X(_10499_));
 sky130_fd_sc_hd__nand2_4 _41036_ (.A(_05966_),
    .B(_10499_),
    .Y(_10500_));
 sky130_fd_sc_hd__buf_1 _41037_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10501_));
 sky130_fd_sc_hd__buf_1 _41038_ (.A(_10501_),
    .X(_10502_));
 sky130_fd_sc_hd__nand2_4 _41039_ (.A(_07359_),
    .B(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__nand2_4 _41040_ (.A(_10500_),
    .B(_10503_),
    .Y(_10504_));
 sky130_fd_sc_hd__buf_1 _41041_ (.A(_03605_),
    .X(_10505_));
 sky130_fd_sc_hd__buf_1 _41042_ (.A(_03612_),
    .X(_10506_));
 sky130_fd_sc_hd__nand4_4 _41043_ (.A(_06746_),
    .B(_05936_),
    .C(_10505_),
    .D(_10506_),
    .Y(_10507_));
 sky130_fd_sc_hd__buf_1 _41044_ (.A(\pcpi_mul.rs2[27] ),
    .X(_10508_));
 sky130_fd_sc_hd__buf_1 _41045_ (.A(_10508_),
    .X(_10509_));
 sky130_fd_sc_hd__nand2_4 _41046_ (.A(_06385_),
    .B(_10509_),
    .Y(_10510_));
 sky130_fd_sc_hd__a21bo_4 _41047_ (.A1(_10504_),
    .A2(_10507_),
    .B1_N(_10510_),
    .X(_10511_));
 sky130_fd_sc_hd__buf_1 _41048_ (.A(_10508_),
    .X(_10512_));
 sky130_fd_sc_hd__buf_1 _41049_ (.A(_10512_),
    .X(_10513_));
 sky130_fd_sc_hd__nand4_4 _41050_ (.A(_05944_),
    .B(_10504_),
    .C(_10507_),
    .D(_10513_),
    .Y(_10514_));
 sky130_fd_sc_hd__buf_1 _41051_ (.A(\pcpi_mul.rs2[30] ),
    .X(_10515_));
 sky130_fd_sc_hd__buf_1 _41052_ (.A(_10515_),
    .X(_10516_));
 sky130_fd_sc_hd__buf_1 _41053_ (.A(_10516_),
    .X(_10517_));
 sky130_fd_sc_hd__nand2_4 _41054_ (.A(_05585_),
    .B(_10517_),
    .Y(_10518_));
 sky130_vsdinv _41055_ (.A(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__a21o_4 _41056_ (.A1(_10511_),
    .A2(_10514_),
    .B1(_10519_),
    .X(_10520_));
 sky130_fd_sc_hd__nand3_4 _41057_ (.A(_10511_),
    .B(_10519_),
    .C(_10514_),
    .Y(_10521_));
 sky130_fd_sc_hd__and2_4 _41058_ (.A(_10520_),
    .B(_10521_),
    .X(_10522_));
 sky130_vsdinv _41059_ (.A(_10522_),
    .Y(_10523_));
 sky130_fd_sc_hd__nand2_4 _41060_ (.A(_10497_),
    .B(_10523_),
    .Y(_10524_));
 sky130_fd_sc_hd__nand3_4 _41061_ (.A(_10522_),
    .B(_10494_),
    .C(_10496_),
    .Y(_10525_));
 sky130_fd_sc_hd__nand2_4 _41062_ (.A(_10524_),
    .B(_10525_),
    .Y(_10526_));
 sky130_fd_sc_hd__nand2_4 _41063_ (.A(_10526_),
    .B(_10332_),
    .Y(_10527_));
 sky130_vsdinv _41064_ (.A(_10332_),
    .Y(_10528_));
 sky130_fd_sc_hd__nand3_4 _41065_ (.A(_10524_),
    .B(_10528_),
    .C(_10525_),
    .Y(_10529_));
 sky130_fd_sc_hd__nand2_4 _41066_ (.A(_10527_),
    .B(_10529_),
    .Y(_10530_));
 sky130_fd_sc_hd__a21boi_4 _41067_ (.A1(_10313_),
    .A2(_10318_),
    .B1_N(_10314_),
    .Y(_10531_));
 sky130_vsdinv _41068_ (.A(_10531_),
    .Y(_10532_));
 sky130_fd_sc_hd__nand2_4 _41069_ (.A(_06251_),
    .B(_10275_),
    .Y(_10533_));
 sky130_fd_sc_hd__nand2_4 _41070_ (.A(_06346_),
    .B(_03569_),
    .Y(_10534_));
 sky130_fd_sc_hd__nand2_4 _41071_ (.A(_10533_),
    .B(_10534_),
    .Y(_10535_));
 sky130_fd_sc_hd__buf_1 _41072_ (.A(_08857_),
    .X(_10536_));
 sky130_fd_sc_hd__buf_1 _41073_ (.A(_09313_),
    .X(_10537_));
 sky130_fd_sc_hd__nand4_4 _41074_ (.A(_06155_),
    .B(_06255_),
    .C(_10536_),
    .D(_10537_),
    .Y(_10538_));
 sky130_fd_sc_hd__nand2_4 _41075_ (.A(_10535_),
    .B(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__buf_1 _41076_ (.A(_03563_),
    .X(_10540_));
 sky130_fd_sc_hd__nand2_4 _41077_ (.A(_06447_),
    .B(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__nand2_4 _41078_ (.A(_10539_),
    .B(_10541_),
    .Y(_10542_));
 sky130_fd_sc_hd__nand4_4 _41079_ (.A(_06565_),
    .B(_10535_),
    .C(_10538_),
    .D(_08636_),
    .Y(_10543_));
 sky130_fd_sc_hd__nand2_4 _41080_ (.A(_10542_),
    .B(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__a21boi_4 _41081_ (.A1(_10274_),
    .A2(_10280_),
    .B1_N(_10276_),
    .Y(_10545_));
 sky130_fd_sc_hd__nand2_4 _41082_ (.A(_10544_),
    .B(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__nand2_4 _41083_ (.A(_10281_),
    .B(_10276_),
    .Y(_10547_));
 sky130_fd_sc_hd__nand3_4 _41084_ (.A(_10547_),
    .B(_10543_),
    .C(_10542_),
    .Y(_10548_));
 sky130_fd_sc_hd__nand2_4 _41085_ (.A(_10546_),
    .B(_10548_),
    .Y(_10549_));
 sky130_fd_sc_hd__nand2_4 _41086_ (.A(_06455_),
    .B(_09486_),
    .Y(_10550_));
 sky130_fd_sc_hd__nand2_4 _41087_ (.A(_06843_),
    .B(_07976_),
    .Y(_10551_));
 sky130_fd_sc_hd__nand2_4 _41088_ (.A(_10550_),
    .B(_10551_),
    .Y(_10552_));
 sky130_fd_sc_hd__nand4_4 _41089_ (.A(_07952_),
    .B(_08607_),
    .C(_10262_),
    .D(_09415_),
    .Y(_10553_));
 sky130_fd_sc_hd__nand2_4 _41090_ (.A(_07819_),
    .B(_07979_),
    .Y(_10554_));
 sky130_vsdinv _41091_ (.A(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__a21o_4 _41092_ (.A1(_10552_),
    .A2(_10553_),
    .B1(_10555_),
    .X(_10556_));
 sky130_fd_sc_hd__nand3_4 _41093_ (.A(_10552_),
    .B(_10553_),
    .C(_10555_),
    .Y(_10557_));
 sky130_fd_sc_hd__and2_4 _41094_ (.A(_10556_),
    .B(_10557_),
    .X(_10558_));
 sky130_vsdinv _41095_ (.A(_10558_),
    .Y(_10559_));
 sky130_fd_sc_hd__nand2_4 _41096_ (.A(_10549_),
    .B(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__nand3_4 _41097_ (.A(_10558_),
    .B(_10546_),
    .C(_10548_),
    .Y(_10561_));
 sky130_fd_sc_hd__nand3_4 _41098_ (.A(_10532_),
    .B(_10560_),
    .C(_10561_),
    .Y(_10562_));
 sky130_fd_sc_hd__nand2_4 _41099_ (.A(_10560_),
    .B(_10561_),
    .Y(_10563_));
 sky130_fd_sc_hd__nand2_4 _41100_ (.A(_10563_),
    .B(_10531_),
    .Y(_10564_));
 sky130_fd_sc_hd__nand2_4 _41101_ (.A(_10562_),
    .B(_10564_),
    .Y(_10565_));
 sky130_fd_sc_hd__a21boi_4 _41102_ (.A1(_10268_),
    .A2(_10284_),
    .B1_N(_10286_),
    .Y(_10566_));
 sky130_fd_sc_hd__nand2_4 _41103_ (.A(_10565_),
    .B(_10566_),
    .Y(_10567_));
 sky130_vsdinv _41104_ (.A(_10566_),
    .Y(_10568_));
 sky130_fd_sc_hd__nand3_4 _41105_ (.A(_10562_),
    .B(_10564_),
    .C(_10568_),
    .Y(_10569_));
 sky130_fd_sc_hd__nand2_4 _41106_ (.A(_10567_),
    .B(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__nand2_4 _41107_ (.A(_10530_),
    .B(_10570_),
    .Y(_10571_));
 sky130_fd_sc_hd__nand4_4 _41108_ (.A(_10569_),
    .B(_10527_),
    .C(_10567_),
    .D(_10529_),
    .Y(_10572_));
 sky130_fd_sc_hd__nand2_4 _41109_ (.A(_10571_),
    .B(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__nand3_4 _41110_ (.A(_10573_),
    .B(_10336_),
    .C(_10339_),
    .Y(_10574_));
 sky130_fd_sc_hd__nand2_4 _41111_ (.A(_10339_),
    .B(_10336_),
    .Y(_10575_));
 sky130_fd_sc_hd__nand3_4 _41112_ (.A(_10575_),
    .B(_10572_),
    .C(_10571_),
    .Y(_10576_));
 sky130_fd_sc_hd__nand2_4 _41113_ (.A(_10574_),
    .B(_10576_),
    .Y(_10577_));
 sky130_vsdinv _41114_ (.A(_10260_),
    .Y(_10578_));
 sky130_fd_sc_hd__a21boi_4 _41115_ (.A1(_10264_),
    .A2(_10578_),
    .B1_N(_10266_),
    .Y(_10579_));
 sky130_vsdinv _41116_ (.A(_10579_),
    .Y(_10580_));
 sky130_fd_sc_hd__nand2_4 _41117_ (.A(_06999_),
    .B(_08566_),
    .Y(_10581_));
 sky130_fd_sc_hd__nand2_4 _41118_ (.A(_07152_),
    .B(_08568_),
    .Y(_10582_));
 sky130_fd_sc_hd__nand2_4 _41119_ (.A(_10581_),
    .B(_10582_),
    .Y(_10583_));
 sky130_fd_sc_hd__buf_1 _41120_ (.A(_06851_),
    .X(_10584_));
 sky130_fd_sc_hd__nand4_4 _41121_ (.A(_10584_),
    .B(_06992_),
    .C(_08128_),
    .D(_07710_),
    .Y(_10585_));
 sky130_fd_sc_hd__nand2_4 _41122_ (.A(_07157_),
    .B(_07719_),
    .Y(_10586_));
 sky130_vsdinv _41123_ (.A(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__nand3_4 _41124_ (.A(_10583_),
    .B(_10585_),
    .C(_10587_),
    .Y(_10588_));
 sky130_fd_sc_hd__nand2_4 _41125_ (.A(_10583_),
    .B(_10585_),
    .Y(_10589_));
 sky130_fd_sc_hd__nand2_4 _41126_ (.A(_10589_),
    .B(_10586_),
    .Y(_10590_));
 sky130_fd_sc_hd__nand3_4 _41127_ (.A(_10580_),
    .B(_10588_),
    .C(_10590_),
    .Y(_10591_));
 sky130_fd_sc_hd__nand2_4 _41128_ (.A(_10590_),
    .B(_10588_),
    .Y(_10592_));
 sky130_fd_sc_hd__nand2_4 _41129_ (.A(_10592_),
    .B(_10579_),
    .Y(_10593_));
 sky130_fd_sc_hd__nand2_4 _41130_ (.A(_10591_),
    .B(_10593_),
    .Y(_10594_));
 sky130_fd_sc_hd__a21boi_4 _41131_ (.A1(_10225_),
    .A2(_10228_),
    .B1_N(_10226_),
    .Y(_10595_));
 sky130_fd_sc_hd__nand2_4 _41132_ (.A(_10594_),
    .B(_10595_),
    .Y(_10596_));
 sky130_vsdinv _41133_ (.A(_10595_),
    .Y(_10597_));
 sky130_fd_sc_hd__nand3_4 _41134_ (.A(_10591_),
    .B(_10593_),
    .C(_10597_),
    .Y(_10598_));
 sky130_fd_sc_hd__nand2_4 _41135_ (.A(_10596_),
    .B(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__a21boi_4 _41136_ (.A1(_10234_),
    .A2(_10238_),
    .B1_N(_10232_),
    .Y(_10600_));
 sky130_fd_sc_hd__nand2_4 _41137_ (.A(_10599_),
    .B(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__nand2_4 _41138_ (.A(_10239_),
    .B(_10232_),
    .Y(_10602_));
 sky130_fd_sc_hd__nand3_4 _41139_ (.A(_10602_),
    .B(_10598_),
    .C(_10596_),
    .Y(_10603_));
 sky130_fd_sc_hd__nand2_4 _41140_ (.A(_10601_),
    .B(_10603_),
    .Y(_10604_));
 sky130_fd_sc_hd__buf_1 _41141_ (.A(_07434_),
    .X(_10605_));
 sky130_fd_sc_hd__nand2_4 _41142_ (.A(_10605_),
    .B(_07741_),
    .Y(_10606_));
 sky130_fd_sc_hd__nand2_4 _41143_ (.A(_08032_),
    .B(_07940_),
    .Y(_10607_));
 sky130_fd_sc_hd__nand2_4 _41144_ (.A(_10606_),
    .B(_10607_),
    .Y(_10608_));
 sky130_fd_sc_hd__nand4_4 _41145_ (.A(_10605_),
    .B(_07626_),
    .C(_07940_),
    .D(_07941_),
    .Y(_10609_));
 sky130_fd_sc_hd__nand2_4 _41146_ (.A(_10212_),
    .B(_03512_),
    .Y(_10610_));
 sky130_vsdinv _41147_ (.A(_10610_),
    .Y(_10611_));
 sky130_fd_sc_hd__a21o_4 _41148_ (.A1(_10608_),
    .A2(_10609_),
    .B1(_10611_),
    .X(_10612_));
 sky130_fd_sc_hd__nand3_4 _41149_ (.A(_10608_),
    .B(_10609_),
    .C(_10611_),
    .Y(_10613_));
 sky130_fd_sc_hd__nand2_4 _41150_ (.A(_10612_),
    .B(_10613_),
    .Y(_10614_));
 sky130_fd_sc_hd__a21boi_4 _41151_ (.A1(_10197_),
    .A2(_10201_),
    .B1_N(_10199_),
    .Y(_10615_));
 sky130_fd_sc_hd__nand2_4 _41152_ (.A(_10614_),
    .B(_10615_),
    .Y(_10616_));
 sky130_vsdinv _41153_ (.A(_10615_),
    .Y(_10617_));
 sky130_fd_sc_hd__nand3_4 _41154_ (.A(_10617_),
    .B(_10613_),
    .C(_10612_),
    .Y(_10618_));
 sky130_fd_sc_hd__buf_1 _41155_ (.A(_03341_),
    .X(_10619_));
 sky130_fd_sc_hd__nand2_4 _41156_ (.A(_10619_),
    .B(_07344_),
    .Y(_10620_));
 sky130_fd_sc_hd__buf_1 _41157_ (.A(_08055_),
    .X(_10621_));
 sky130_fd_sc_hd__nand2_4 _41158_ (.A(_10621_),
    .B(_07347_),
    .Y(_10622_));
 sky130_fd_sc_hd__nand2_4 _41159_ (.A(_10620_),
    .B(_10622_),
    .Y(_10623_));
 sky130_fd_sc_hd__buf_1 _41160_ (.A(_08733_),
    .X(_10624_));
 sky130_fd_sc_hd__buf_1 _41161_ (.A(_08522_),
    .X(_10625_));
 sky130_fd_sc_hd__nand4_4 _41162_ (.A(_10624_),
    .B(_10625_),
    .C(_06506_),
    .D(_06637_),
    .Y(_10626_));
 sky130_fd_sc_hd__nand2_4 _41163_ (.A(_08753_),
    .B(_07205_),
    .Y(_10627_));
 sky130_vsdinv _41164_ (.A(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__a21o_4 _41165_ (.A1(_10623_),
    .A2(_10626_),
    .B1(_10628_),
    .X(_10629_));
 sky130_fd_sc_hd__nand3_4 _41166_ (.A(_10623_),
    .B(_10626_),
    .C(_10628_),
    .Y(_10630_));
 sky130_fd_sc_hd__nand2_4 _41167_ (.A(_10629_),
    .B(_10630_),
    .Y(_10631_));
 sky130_vsdinv _41168_ (.A(_10631_),
    .Y(_10632_));
 sky130_fd_sc_hd__a21o_4 _41169_ (.A1(_10616_),
    .A2(_10618_),
    .B1(_10632_),
    .X(_10633_));
 sky130_fd_sc_hd__nand3_4 _41170_ (.A(_10616_),
    .B(_10618_),
    .C(_10632_),
    .Y(_10634_));
 sky130_fd_sc_hd__and2_4 _41171_ (.A(_10633_),
    .B(_10634_),
    .X(_10635_));
 sky130_vsdinv _41172_ (.A(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__nand2_4 _41173_ (.A(_10604_),
    .B(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__nand3_4 _41174_ (.A(_10635_),
    .B(_10601_),
    .C(_10603_),
    .Y(_10638_));
 sky130_fd_sc_hd__nand2_4 _41175_ (.A(_10637_),
    .B(_10638_),
    .Y(_10639_));
 sky130_vsdinv _41176_ (.A(_10293_),
    .Y(_10640_));
 sky130_fd_sc_hd__a21oi_4 _41177_ (.A1(_10291_),
    .A2(_10297_),
    .B1(_10640_),
    .Y(_10641_));
 sky130_fd_sc_hd__nand2_4 _41178_ (.A(_10639_),
    .B(_10641_),
    .Y(_10642_));
 sky130_vsdinv _41179_ (.A(_10641_),
    .Y(_10643_));
 sky130_fd_sc_hd__nand3_4 _41180_ (.A(_10643_),
    .B(_10638_),
    .C(_10637_),
    .Y(_10644_));
 sky130_fd_sc_hd__nand2_4 _41181_ (.A(_10642_),
    .B(_10644_),
    .Y(_10645_));
 sky130_fd_sc_hd__a21boi_4 _41182_ (.A1(_10219_),
    .A2(_10242_),
    .B1_N(_10244_),
    .Y(_10646_));
 sky130_fd_sc_hd__nand2_4 _41183_ (.A(_10645_),
    .B(_10646_),
    .Y(_10647_));
 sky130_vsdinv _41184_ (.A(_10646_),
    .Y(_10648_));
 sky130_fd_sc_hd__nand3_4 _41185_ (.A(_10642_),
    .B(_10644_),
    .C(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__nand2_4 _41186_ (.A(_10647_),
    .B(_10649_),
    .Y(_10650_));
 sky130_fd_sc_hd__nand2_4 _41187_ (.A(_10577_),
    .B(_10650_),
    .Y(_10651_));
 sky130_fd_sc_hd__nand4_4 _41188_ (.A(_10649_),
    .B(_10574_),
    .C(_10647_),
    .D(_10576_),
    .Y(_10652_));
 sky130_fd_sc_hd__nand2_4 _41189_ (.A(_10651_),
    .B(_10652_),
    .Y(_10653_));
 sky130_vsdinv _41190_ (.A(_10343_),
    .Y(_10654_));
 sky130_fd_sc_hd__o21a_4 _41191_ (.A1(_10654_),
    .A2(_10259_),
    .B1(_10344_),
    .X(_10655_));
 sky130_fd_sc_hd__nand2_4 _41192_ (.A(_10653_),
    .B(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__o21ai_4 _41193_ (.A1(_10654_),
    .A2(_10259_),
    .B1(_10344_),
    .Y(_10657_));
 sky130_fd_sc_hd__nand3_4 _41194_ (.A(_10657_),
    .B(_10652_),
    .C(_10651_),
    .Y(_10658_));
 sky130_fd_sc_hd__nand2_4 _41195_ (.A(_10656_),
    .B(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__nand2_4 _41196_ (.A(_10218_),
    .B(_10204_),
    .Y(_10660_));
 sky130_fd_sc_hd__nand2_4 _41197_ (.A(_09087_),
    .B(_06372_),
    .Y(_10661_));
 sky130_fd_sc_hd__nand2_4 _41198_ (.A(_09088_),
    .B(_06477_),
    .Y(_10662_));
 sky130_fd_sc_hd__nand2_4 _41199_ (.A(_10661_),
    .B(_10662_),
    .Y(_10663_));
 sky130_fd_sc_hd__buf_1 _41200_ (.A(_08530_),
    .X(_10664_));
 sky130_fd_sc_hd__nand4_4 _41201_ (.A(_10664_),
    .B(_09831_),
    .C(_03481_),
    .D(_06939_),
    .Y(_10665_));
 sky130_fd_sc_hd__buf_1 _41202_ (.A(_03365_),
    .X(_10666_));
 sky130_fd_sc_hd__nand2_4 _41203_ (.A(_10666_),
    .B(_06606_),
    .Y(_10667_));
 sky130_vsdinv _41204_ (.A(_10667_),
    .Y(_10668_));
 sky130_fd_sc_hd__a21o_4 _41205_ (.A1(_10663_),
    .A2(_10665_),
    .B1(_10668_),
    .X(_10669_));
 sky130_fd_sc_hd__nand3_4 _41206_ (.A(_10663_),
    .B(_10665_),
    .C(_10668_),
    .Y(_10670_));
 sky130_fd_sc_hd__nand2_4 _41207_ (.A(_10669_),
    .B(_10670_),
    .Y(_10671_));
 sky130_vsdinv _41208_ (.A(_10208_),
    .Y(_10672_));
 sky130_fd_sc_hd__a21boi_4 _41209_ (.A1(_10211_),
    .A2(_10672_),
    .B1_N(_10213_),
    .Y(_10673_));
 sky130_fd_sc_hd__nand2_4 _41210_ (.A(_10671_),
    .B(_10673_),
    .Y(_10674_));
 sky130_vsdinv _41211_ (.A(_10673_),
    .Y(_10675_));
 sky130_fd_sc_hd__nand3_4 _41212_ (.A(_10675_),
    .B(_10669_),
    .C(_10670_),
    .Y(_10676_));
 sky130_fd_sc_hd__a21boi_4 _41213_ (.A1(_10359_),
    .A2(_10364_),
    .B1_N(_10360_),
    .Y(_10677_));
 sky130_vsdinv _41214_ (.A(_10677_),
    .Y(_10678_));
 sky130_fd_sc_hd__nand3_4 _41215_ (.A(_10674_),
    .B(_10676_),
    .C(_10678_),
    .Y(_10679_));
 sky130_fd_sc_hd__nand2_4 _41216_ (.A(_10674_),
    .B(_10676_),
    .Y(_10680_));
 sky130_fd_sc_hd__nand2_4 _41217_ (.A(_10680_),
    .B(_10677_),
    .Y(_10681_));
 sky130_fd_sc_hd__nand3_4 _41218_ (.A(_10660_),
    .B(_10679_),
    .C(_10681_),
    .Y(_10682_));
 sky130_fd_sc_hd__nand2_4 _41219_ (.A(_10681_),
    .B(_10679_),
    .Y(_10683_));
 sky130_fd_sc_hd__a21boi_4 _41220_ (.A1(_10215_),
    .A2(_10206_),
    .B1_N(_10204_),
    .Y(_10684_));
 sky130_fd_sc_hd__nand2_4 _41221_ (.A(_10683_),
    .B(_10684_),
    .Y(_10685_));
 sky130_fd_sc_hd__nand2_4 _41222_ (.A(_10682_),
    .B(_10685_),
    .Y(_10686_));
 sky130_fd_sc_hd__a21boi_4 _41223_ (.A1(_10368_),
    .A2(_10370_),
    .B1_N(_10366_),
    .Y(_10687_));
 sky130_fd_sc_hd__nand2_4 _41224_ (.A(_10686_),
    .B(_10687_),
    .Y(_10688_));
 sky130_vsdinv _41225_ (.A(_10687_),
    .Y(_10689_));
 sky130_fd_sc_hd__nand3_4 _41226_ (.A(_10682_),
    .B(_10685_),
    .C(_10689_),
    .Y(_10690_));
 sky130_fd_sc_hd__nand2_4 _41227_ (.A(_10688_),
    .B(_10690_),
    .Y(_10691_));
 sky130_fd_sc_hd__a21boi_4 _41228_ (.A1(_10377_),
    .A2(_10381_),
    .B1_N(_10374_),
    .Y(_10692_));
 sky130_fd_sc_hd__nand2_4 _41229_ (.A(_10691_),
    .B(_10692_),
    .Y(_10693_));
 sky130_vsdinv _41230_ (.A(_10692_),
    .Y(_10694_));
 sky130_fd_sc_hd__nand3_4 _41231_ (.A(_10694_),
    .B(_10690_),
    .C(_10688_),
    .Y(_10695_));
 sky130_fd_sc_hd__nand2_4 _41232_ (.A(_10693_),
    .B(_10695_),
    .Y(_10696_));
 sky130_vsdinv _41233_ (.A(_10402_),
    .Y(_10697_));
 sky130_fd_sc_hd__a21oi_4 _41234_ (.A1(_10400_),
    .A2(_10415_),
    .B1(_10697_),
    .Y(_10698_));
 sky130_vsdinv _41235_ (.A(_10698_),
    .Y(_10699_));
 sky130_fd_sc_hd__nand2_4 _41236_ (.A(_09214_),
    .B(_06314_),
    .Y(_10700_));
 sky130_fd_sc_hd__nand2_4 _41237_ (.A(_10393_),
    .B(_08507_),
    .Y(_10701_));
 sky130_fd_sc_hd__nand2_4 _41238_ (.A(_10700_),
    .B(_10701_),
    .Y(_10702_));
 sky130_fd_sc_hd__buf_1 _41239_ (.A(_03374_),
    .X(_10703_));
 sky130_fd_sc_hd__nand4_4 _41240_ (.A(_10703_),
    .B(_10083_),
    .C(_05963_),
    .D(_05989_),
    .Y(_10704_));
 sky130_fd_sc_hd__nand2_4 _41241_ (.A(_09849_),
    .B(_06327_),
    .Y(_10705_));
 sky130_vsdinv _41242_ (.A(_10705_),
    .Y(_10706_));
 sky130_fd_sc_hd__a21o_4 _41243_ (.A1(_10702_),
    .A2(_10704_),
    .B1(_10706_),
    .X(_10707_));
 sky130_fd_sc_hd__nand3_4 _41244_ (.A(_10702_),
    .B(_10704_),
    .C(_10706_),
    .Y(_10708_));
 sky130_fd_sc_hd__a21boi_4 _41245_ (.A1(_10391_),
    .A2(_10395_),
    .B1_N(_10392_),
    .Y(_10709_));
 sky130_fd_sc_hd__a21boi_4 _41246_ (.A1(_10707_),
    .A2(_10708_),
    .B1_N(_10709_),
    .Y(_10710_));
 sky130_fd_sc_hd__nand2_4 _41247_ (.A(_10707_),
    .B(_10708_),
    .Y(_10711_));
 sky130_fd_sc_hd__nor2_4 _41248_ (.A(_10709_),
    .B(_10711_),
    .Y(_10712_));
 sky130_fd_sc_hd__nand2_4 _41249_ (.A(_10406_),
    .B(_08043_),
    .Y(_10713_));
 sky130_fd_sc_hd__o21ai_4 _41250_ (.A1(_03394_),
    .A2(_05892_),
    .B1(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__buf_1 _41251_ (.A(_10408_),
    .X(_10715_));
 sky130_fd_sc_hd__nand4_4 _41252_ (.A(_10087_),
    .B(_10715_),
    .C(_07440_),
    .D(_03443_),
    .Y(_10716_));
 sky130_fd_sc_hd__nand2_4 _41253_ (.A(_03396_),
    .B(_03419_),
    .Y(_10717_));
 sky130_vsdinv _41254_ (.A(_10717_),
    .Y(_10718_));
 sky130_fd_sc_hd__a21o_4 _41255_ (.A1(_10714_),
    .A2(_10716_),
    .B1(_10718_),
    .X(_10719_));
 sky130_fd_sc_hd__nand3_4 _41256_ (.A(_10714_),
    .B(_10716_),
    .C(_10718_),
    .Y(_10720_));
 sky130_fd_sc_hd__and2_4 _41257_ (.A(_10719_),
    .B(_10720_),
    .X(_10721_));
 sky130_vsdinv _41258_ (.A(_10721_),
    .Y(_10722_));
 sky130_fd_sc_hd__o21ai_4 _41259_ (.A1(_10710_),
    .A2(_10712_),
    .B1(_10722_),
    .Y(_10723_));
 sky130_vsdinv _41260_ (.A(_10712_),
    .Y(_10724_));
 sky130_vsdinv _41261_ (.A(_10710_),
    .Y(_10725_));
 sky130_fd_sc_hd__nand3_4 _41262_ (.A(_10724_),
    .B(_10725_),
    .C(_10721_),
    .Y(_10726_));
 sky130_fd_sc_hd__nand3_4 _41263_ (.A(_10699_),
    .B(_10723_),
    .C(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__nand2_4 _41264_ (.A(_10723_),
    .B(_10726_),
    .Y(_10728_));
 sky130_fd_sc_hd__nand2_4 _41265_ (.A(_10728_),
    .B(_10698_),
    .Y(_10729_));
 sky130_fd_sc_hd__a21boi_4 _41266_ (.A1(_10404_),
    .A2(_10411_),
    .B1_N(_10407_),
    .Y(_10730_));
 sky130_vsdinv _41267_ (.A(_10730_),
    .Y(_10731_));
 sky130_fd_sc_hd__a21oi_4 _41268_ (.A1(_10727_),
    .A2(_10729_),
    .B1(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__nand3_4 _41269_ (.A(_10727_),
    .B(_10729_),
    .C(_10731_),
    .Y(_10733_));
 sky130_vsdinv _41270_ (.A(_10733_),
    .Y(_10734_));
 sky130_fd_sc_hd__nor2_4 _41271_ (.A(_10732_),
    .B(_10734_),
    .Y(_10735_));
 sky130_vsdinv _41272_ (.A(_10735_),
    .Y(_10736_));
 sky130_fd_sc_hd__nand2_4 _41273_ (.A(_10696_),
    .B(_10736_),
    .Y(_10737_));
 sky130_fd_sc_hd__nand3_4 _41274_ (.A(_10735_),
    .B(_10693_),
    .C(_10695_),
    .Y(_10738_));
 sky130_fd_sc_hd__nand2_4 _41275_ (.A(_10737_),
    .B(_10738_),
    .Y(_10739_));
 sky130_fd_sc_hd__a21boi_4 _41276_ (.A1(_10251_),
    .A2(_10257_),
    .B1_N(_10253_),
    .Y(_10740_));
 sky130_fd_sc_hd__nand2_4 _41277_ (.A(_10739_),
    .B(_10740_),
    .Y(_10741_));
 sky130_vsdinv _41278_ (.A(_10740_),
    .Y(_10742_));
 sky130_fd_sc_hd__nand3_4 _41279_ (.A(_10742_),
    .B(_10738_),
    .C(_10737_),
    .Y(_10743_));
 sky130_fd_sc_hd__nand2_4 _41280_ (.A(_10741_),
    .B(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__o21a_4 _41281_ (.A1(_10428_),
    .A2(_10388_),
    .B1(_10387_),
    .X(_10745_));
 sky130_fd_sc_hd__nand2_4 _41282_ (.A(_10744_),
    .B(_10745_),
    .Y(_10746_));
 sky130_vsdinv _41283_ (.A(_10745_),
    .Y(_10747_));
 sky130_fd_sc_hd__nand3_4 _41284_ (.A(_10741_),
    .B(_10747_),
    .C(_10743_),
    .Y(_10748_));
 sky130_fd_sc_hd__nand2_4 _41285_ (.A(_10746_),
    .B(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__nand2_4 _41286_ (.A(_10659_),
    .B(_10749_),
    .Y(_10750_));
 sky130_fd_sc_hd__nand4_4 _41287_ (.A(_10748_),
    .B(_10656_),
    .C(_10746_),
    .D(_10658_),
    .Y(_10751_));
 sky130_fd_sc_hd__nand2_4 _41288_ (.A(_10750_),
    .B(_10751_),
    .Y(_10752_));
 sky130_fd_sc_hd__nand2_4 _41289_ (.A(_10475_),
    .B(_10752_),
    .Y(_10753_));
 sky130_fd_sc_hd__nand2_4 _41290_ (.A(_10443_),
    .B(_10351_),
    .Y(_10754_));
 sky130_fd_sc_hd__nand3_4 _41291_ (.A(_10754_),
    .B(_10751_),
    .C(_10750_),
    .Y(_10755_));
 sky130_fd_sc_hd__nand2_4 _41292_ (.A(_10753_),
    .B(_10755_),
    .Y(_10756_));
 sky130_fd_sc_hd__o21a_4 _41293_ (.A1(_10423_),
    .A2(_10420_),
    .B1(_10421_),
    .X(_10757_));
 sky130_fd_sc_hd__a21boi_4 _41294_ (.A1(_10433_),
    .A2(_10439_),
    .B1_N(_10435_),
    .Y(_10758_));
 sky130_fd_sc_hd__xnor2_4 _41295_ (.A(_10757_),
    .B(_10758_),
    .Y(_10759_));
 sky130_fd_sc_hd__nand2_4 _41296_ (.A(_10756_),
    .B(_10759_),
    .Y(_10760_));
 sky130_vsdinv _41297_ (.A(_10759_),
    .Y(_10761_));
 sky130_fd_sc_hd__nand3_4 _41298_ (.A(_10753_),
    .B(_10755_),
    .C(_10761_),
    .Y(_10762_));
 sky130_fd_sc_hd__nand2_4 _41299_ (.A(_10760_),
    .B(_10762_),
    .Y(_10763_));
 sky130_fd_sc_hd__nand2_4 _41300_ (.A(_10456_),
    .B(_10449_),
    .Y(_10764_));
 sky130_vsdinv _41301_ (.A(_10764_),
    .Y(_10765_));
 sky130_fd_sc_hd__nand2_4 _41302_ (.A(_10763_),
    .B(_10765_),
    .Y(_10766_));
 sky130_fd_sc_hd__nand3_4 _41303_ (.A(_10764_),
    .B(_10760_),
    .C(_10762_),
    .Y(_10767_));
 sky130_fd_sc_hd__nand2_4 _41304_ (.A(_10766_),
    .B(_10767_),
    .Y(_10768_));
 sky130_fd_sc_hd__a21oi_4 _41305_ (.A1(_10156_),
    .A2(_10151_),
    .B1(_10451_),
    .Y(_10769_));
 sky130_vsdinv _41306_ (.A(_10769_),
    .Y(_10770_));
 sky130_fd_sc_hd__nand2_4 _41307_ (.A(_10768_),
    .B(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__nand3_4 _41308_ (.A(_10766_),
    .B(_10769_),
    .C(_10767_),
    .Y(_10772_));
 sky130_fd_sc_hd__nand2_4 _41309_ (.A(_10771_),
    .B(_10772_),
    .Y(_10773_));
 sky130_fd_sc_hd__nand2_4 _41310_ (.A(_10466_),
    .B(_10461_),
    .Y(_10774_));
 sky130_vsdinv _41311_ (.A(_10774_),
    .Y(_10775_));
 sky130_fd_sc_hd__nand2_4 _41312_ (.A(_10773_),
    .B(_10775_),
    .Y(_10776_));
 sky130_fd_sc_hd__nand3_4 _41313_ (.A(_10774_),
    .B(_10771_),
    .C(_10772_),
    .Y(_10777_));
 sky130_fd_sc_hd__and2_4 _41314_ (.A(_10776_),
    .B(_10777_),
    .X(_10778_));
 sky130_fd_sc_hd__buf_1 _41315_ (.A(_10778_),
    .X(_10779_));
 sky130_vsdinv _41316_ (.A(_10779_),
    .Y(_10780_));
 sky130_fd_sc_hd__o21ai_4 _41317_ (.A1(_10182_),
    .A2(_10181_),
    .B1(_10471_),
    .Y(_10781_));
 sky130_fd_sc_hd__a32oi_4 _41318_ (.A1(_10192_),
    .A2(_10187_),
    .A3(_10473_),
    .B1(_10470_),
    .B2(_10781_),
    .Y(_10782_));
 sky130_fd_sc_hd__xor2_4 _41319_ (.A(_10780_),
    .B(_10782_),
    .X(_01435_));
 sky130_fd_sc_hd__buf_1 _41320_ (.A(_09565_),
    .X(_10783_));
 sky130_fd_sc_hd__nand2_4 _41321_ (.A(_10783_),
    .B(_06789_),
    .Y(_10784_));
 sky130_fd_sc_hd__buf_1 _41322_ (.A(_09090_),
    .X(_10785_));
 sky130_fd_sc_hd__nand2_4 _41323_ (.A(_10785_),
    .B(_06947_),
    .Y(_10786_));
 sky130_fd_sc_hd__nand2_4 _41324_ (.A(_10784_),
    .B(_10786_),
    .Y(_10787_));
 sky130_fd_sc_hd__buf_1 _41325_ (.A(_08759_),
    .X(_10788_));
 sky130_fd_sc_hd__buf_1 _41326_ (.A(_09833_),
    .X(_10789_));
 sky130_fd_sc_hd__nand4_4 _41327_ (.A(_10788_),
    .B(_10789_),
    .C(_07097_),
    .D(_06794_),
    .Y(_10790_));
 sky130_fd_sc_hd__buf_1 _41328_ (.A(_03375_),
    .X(_10791_));
 sky130_fd_sc_hd__nand2_4 _41329_ (.A(_10791_),
    .B(_06797_),
    .Y(_10792_));
 sky130_vsdinv _41330_ (.A(_10792_),
    .Y(_10793_));
 sky130_fd_sc_hd__a21o_4 _41331_ (.A1(_10787_),
    .A2(_10790_),
    .B1(_10793_),
    .X(_10794_));
 sky130_fd_sc_hd__nand3_4 _41332_ (.A(_10787_),
    .B(_10790_),
    .C(_10793_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand2_4 _41333_ (.A(_10794_),
    .B(_10795_),
    .Y(_10796_));
 sky130_fd_sc_hd__a21boi_4 _41334_ (.A1(_10623_),
    .A2(_10628_),
    .B1_N(_10626_),
    .Y(_10797_));
 sky130_fd_sc_hd__nand2_4 _41335_ (.A(_10796_),
    .B(_10797_),
    .Y(_10798_));
 sky130_vsdinv _41336_ (.A(_10797_),
    .Y(_10799_));
 sky130_fd_sc_hd__nand3_4 _41337_ (.A(_10799_),
    .B(_10794_),
    .C(_10795_),
    .Y(_10800_));
 sky130_fd_sc_hd__a21boi_4 _41338_ (.A1(_10663_),
    .A2(_10668_),
    .B1_N(_10665_),
    .Y(_10801_));
 sky130_vsdinv _41339_ (.A(_10801_),
    .Y(_10802_));
 sky130_fd_sc_hd__a21o_4 _41340_ (.A1(_10798_),
    .A2(_10800_),
    .B1(_10802_),
    .X(_10803_));
 sky130_fd_sc_hd__nand3_4 _41341_ (.A(_10798_),
    .B(_10800_),
    .C(_10802_),
    .Y(_10804_));
 sky130_fd_sc_hd__nand2_4 _41342_ (.A(_10803_),
    .B(_10804_),
    .Y(_10805_));
 sky130_fd_sc_hd__a21boi_4 _41343_ (.A1(_10616_),
    .A2(_10632_),
    .B1_N(_10618_),
    .Y(_10806_));
 sky130_fd_sc_hd__nand2_4 _41344_ (.A(_10805_),
    .B(_10806_),
    .Y(_10807_));
 sky130_vsdinv _41345_ (.A(_10806_),
    .Y(_10808_));
 sky130_fd_sc_hd__nand3_4 _41346_ (.A(_10808_),
    .B(_10803_),
    .C(_10804_),
    .Y(_10809_));
 sky130_fd_sc_hd__a21boi_4 _41347_ (.A1(_10674_),
    .A2(_10678_),
    .B1_N(_10676_),
    .Y(_10810_));
 sky130_vsdinv _41348_ (.A(_10810_),
    .Y(_10811_));
 sky130_fd_sc_hd__a21o_4 _41349_ (.A1(_10807_),
    .A2(_10809_),
    .B1(_10811_),
    .X(_10812_));
 sky130_fd_sc_hd__nand3_4 _41350_ (.A(_10807_),
    .B(_10809_),
    .C(_10811_),
    .Y(_10813_));
 sky130_fd_sc_hd__nand2_4 _41351_ (.A(_10812_),
    .B(_10813_),
    .Y(_10814_));
 sky130_fd_sc_hd__a21boi_4 _41352_ (.A1(_10689_),
    .A2(_10685_),
    .B1_N(_10682_),
    .Y(_10815_));
 sky130_fd_sc_hd__nand2_4 _41353_ (.A(_10814_),
    .B(_10815_),
    .Y(_10816_));
 sky130_vsdinv _41354_ (.A(_10815_),
    .Y(_10817_));
 sky130_fd_sc_hd__nand3_4 _41355_ (.A(_10817_),
    .B(_10813_),
    .C(_10812_),
    .Y(_10818_));
 sky130_fd_sc_hd__nand2_4 _41356_ (.A(_10816_),
    .B(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__a21boi_4 _41357_ (.A1(_10702_),
    .A2(_10706_),
    .B1_N(_10704_),
    .Y(_10820_));
 sky130_fd_sc_hd__nand2_4 _41358_ (.A(_10080_),
    .B(_06315_),
    .Y(_10821_));
 sky130_fd_sc_hd__buf_1 _41359_ (.A(_03382_),
    .X(_10822_));
 sky130_fd_sc_hd__nand2_4 _41360_ (.A(_10822_),
    .B(_06136_),
    .Y(_10823_));
 sky130_fd_sc_hd__nand2_4 _41361_ (.A(_10821_),
    .B(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__nand4_4 _41362_ (.A(_10084_),
    .B(_10085_),
    .C(_06430_),
    .D(_06432_),
    .Y(_10825_));
 sky130_fd_sc_hd__buf_1 _41363_ (.A(\pcpi_mul.rs1[28] ),
    .X(_10826_));
 sky130_fd_sc_hd__buf_1 _41364_ (.A(_10826_),
    .X(_10827_));
 sky130_fd_sc_hd__nand2_4 _41365_ (.A(_10827_),
    .B(_06328_),
    .Y(_10828_));
 sky130_vsdinv _41366_ (.A(_10828_),
    .Y(_10829_));
 sky130_fd_sc_hd__a21o_4 _41367_ (.A1(_10824_),
    .A2(_10825_),
    .B1(_10829_),
    .X(_10830_));
 sky130_fd_sc_hd__nand3_4 _41368_ (.A(_10824_),
    .B(_10825_),
    .C(_10829_),
    .Y(_10831_));
 sky130_fd_sc_hd__nand2_4 _41369_ (.A(_10830_),
    .B(_10831_),
    .Y(_10832_));
 sky130_fd_sc_hd__nor2_4 _41370_ (.A(_10820_),
    .B(_10832_),
    .Y(_10833_));
 sky130_vsdinv _41371_ (.A(_10833_),
    .Y(_10834_));
 sky130_fd_sc_hd__nand2_4 _41372_ (.A(_10832_),
    .B(_10820_),
    .Y(_10835_));
 sky130_fd_sc_hd__buf_1 _41373_ (.A(\pcpi_mul.rs1[31] ),
    .X(_10836_));
 sky130_fd_sc_hd__buf_1 _41374_ (.A(_10836_),
    .X(_10837_));
 sky130_fd_sc_hd__buf_1 _41375_ (.A(_10837_),
    .X(_10838_));
 sky130_fd_sc_hd__nand2_4 _41376_ (.A(_10838_),
    .B(_03421_),
    .Y(_10839_));
 sky130_fd_sc_hd__buf_1 _41377_ (.A(_10715_),
    .X(_10840_));
 sky130_fd_sc_hd__nand2_4 _41378_ (.A(_10840_),
    .B(_03444_),
    .Y(_10841_));
 sky130_fd_sc_hd__o21ai_4 _41379_ (.A1(_03398_),
    .A2(_05893_),
    .B1(_10841_),
    .Y(_10842_));
 sky130_fd_sc_hd__buf_1 _41380_ (.A(_03393_),
    .X(_10843_));
 sky130_fd_sc_hd__buf_1 _41381_ (.A(_10843_),
    .X(_10844_));
 sky130_fd_sc_hd__buf_1 _41382_ (.A(\pcpi_mul.rs1[30] ),
    .X(_10845_));
 sky130_fd_sc_hd__buf_4 _41383_ (.A(_10845_),
    .X(_10846_));
 sky130_fd_sc_hd__buf_4 _41384_ (.A(_10846_),
    .X(_10847_));
 sky130_fd_sc_hd__nand4_4 _41385_ (.A(_10844_),
    .B(_10847_),
    .C(_05948_),
    .D(_05911_),
    .Y(_10848_));
 sky130_fd_sc_hd__nand2_4 _41386_ (.A(_10842_),
    .B(_10848_),
    .Y(_10849_));
 sky130_fd_sc_hd__xor2_4 _41387_ (.A(_10839_),
    .B(_10849_),
    .X(_10850_));
 sky130_fd_sc_hd__a21o_4 _41388_ (.A1(_10834_),
    .A2(_10835_),
    .B1(_10850_),
    .X(_10851_));
 sky130_fd_sc_hd__nand3_4 _41389_ (.A(_10834_),
    .B(_10850_),
    .C(_10835_),
    .Y(_10852_));
 sky130_fd_sc_hd__a21oi_4 _41390_ (.A1(_10725_),
    .A2(_10721_),
    .B1(_10712_),
    .Y(_10853_));
 sky130_vsdinv _41391_ (.A(_10853_),
    .Y(_10854_));
 sky130_fd_sc_hd__a21o_4 _41392_ (.A1(_10851_),
    .A2(_10852_),
    .B1(_10854_),
    .X(_10855_));
 sky130_fd_sc_hd__nand3_4 _41393_ (.A(_10854_),
    .B(_10851_),
    .C(_10852_),
    .Y(_10856_));
 sky130_fd_sc_hd__a21boi_4 _41394_ (.A1(_10714_),
    .A2(_10718_),
    .B1_N(_10716_),
    .Y(_10857_));
 sky130_vsdinv _41395_ (.A(_10857_),
    .Y(_10858_));
 sky130_fd_sc_hd__a21oi_4 _41396_ (.A1(_10855_),
    .A2(_10856_),
    .B1(_10858_),
    .Y(_10859_));
 sky130_vsdinv _41397_ (.A(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__nand3_4 _41398_ (.A(_10855_),
    .B(_10858_),
    .C(_10856_),
    .Y(_10861_));
 sky130_fd_sc_hd__nand2_4 _41399_ (.A(_10860_),
    .B(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__nand2_4 _41400_ (.A(_10819_),
    .B(_10862_),
    .Y(_10863_));
 sky130_vsdinv _41401_ (.A(_10861_),
    .Y(_10864_));
 sky130_fd_sc_hd__nor2_4 _41402_ (.A(_10859_),
    .B(_10864_),
    .Y(_10865_));
 sky130_fd_sc_hd__nand3_4 _41403_ (.A(_10865_),
    .B(_10816_),
    .C(_10818_),
    .Y(_10866_));
 sky130_fd_sc_hd__nand2_4 _41404_ (.A(_10863_),
    .B(_10866_),
    .Y(_10867_));
 sky130_fd_sc_hd__a21boi_4 _41405_ (.A1(_10642_),
    .A2(_10648_),
    .B1_N(_10644_),
    .Y(_10868_));
 sky130_fd_sc_hd__nand2_4 _41406_ (.A(_10867_),
    .B(_10868_),
    .Y(_10869_));
 sky130_vsdinv _41407_ (.A(_10868_),
    .Y(_10870_));
 sky130_fd_sc_hd__nand3_4 _41408_ (.A(_10870_),
    .B(_10863_),
    .C(_10866_),
    .Y(_10871_));
 sky130_fd_sc_hd__nand2_4 _41409_ (.A(_10869_),
    .B(_10871_),
    .Y(_10872_));
 sky130_fd_sc_hd__a21boi_4 _41410_ (.A1(_10735_),
    .A2(_10693_),
    .B1_N(_10695_),
    .Y(_10873_));
 sky130_fd_sc_hd__nand2_4 _41411_ (.A(_10872_),
    .B(_10873_),
    .Y(_10874_));
 sky130_vsdinv _41412_ (.A(_10873_),
    .Y(_10875_));
 sky130_fd_sc_hd__nand3_4 _41413_ (.A(_10869_),
    .B(_10875_),
    .C(_10871_),
    .Y(_10876_));
 sky130_fd_sc_hd__nand2_4 _41414_ (.A(_10874_),
    .B(_10876_),
    .Y(_10877_));
 sky130_fd_sc_hd__o21a_4 _41415_ (.A1(_10570_),
    .A2(_10530_),
    .B1(_10529_),
    .X(_10878_));
 sky130_fd_sc_hd__nand2_4 _41416_ (.A(_10496_),
    .B(_10491_),
    .Y(_10879_));
 sky130_vsdinv _41417_ (.A(_10879_),
    .Y(_10880_));
 sky130_fd_sc_hd__nand2_4 _41418_ (.A(_07758_),
    .B(_03576_),
    .Y(_10881_));
 sky130_fd_sc_hd__nand2_4 _41419_ (.A(_06451_),
    .B(_10536_),
    .Y(_10882_));
 sky130_fd_sc_hd__nand2_4 _41420_ (.A(_10881_),
    .B(_10882_),
    .Y(_10883_));
 sky130_fd_sc_hd__buf_1 _41421_ (.A(_08630_),
    .X(_10884_));
 sky130_fd_sc_hd__buf_1 _41422_ (.A(_10270_),
    .X(_10885_));
 sky130_fd_sc_hd__nand4_4 _41423_ (.A(_07959_),
    .B(_10265_),
    .C(_10884_),
    .D(_10885_),
    .Y(_10886_));
 sky130_fd_sc_hd__buf_1 _41424_ (.A(_08634_),
    .X(_10887_));
 sky130_fd_sc_hd__nand2_4 _41425_ (.A(_06567_),
    .B(_10887_),
    .Y(_10888_));
 sky130_vsdinv _41426_ (.A(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__a21o_4 _41427_ (.A1(_10883_),
    .A2(_10886_),
    .B1(_10889_),
    .X(_10890_));
 sky130_fd_sc_hd__nand3_4 _41428_ (.A(_10883_),
    .B(_10886_),
    .C(_10889_),
    .Y(_10891_));
 sky130_fd_sc_hd__nand2_4 _41429_ (.A(_10890_),
    .B(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__maj3_4 _41430_ (.A(_10541_),
    .B(_10533_),
    .C(_10534_),
    .X(_10893_));
 sky130_fd_sc_hd__nand2_4 _41431_ (.A(_10892_),
    .B(_10893_),
    .Y(_10894_));
 sky130_fd_sc_hd__nand2_4 _41432_ (.A(_10543_),
    .B(_10538_),
    .Y(_10895_));
 sky130_fd_sc_hd__nand3_4 _41433_ (.A(_10895_),
    .B(_10891_),
    .C(_10890_),
    .Y(_10896_));
 sky130_fd_sc_hd__nand2_4 _41434_ (.A(_10894_),
    .B(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__nand2_4 _41435_ (.A(_08392_),
    .B(_10262_),
    .Y(_10898_));
 sky130_fd_sc_hd__o21ai_4 _41436_ (.A1(_03299_),
    .A2(_03558_),
    .B1(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__buf_1 _41437_ (.A(_06846_),
    .X(_10900_));
 sky130_fd_sc_hd__nand4_4 _41438_ (.A(_10900_),
    .B(_07660_),
    .C(_08191_),
    .D(_08194_),
    .Y(_10901_));
 sky130_fd_sc_hd__nand2_4 _41439_ (.A(_10899_),
    .B(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__nand2_4 _41440_ (.A(_06999_),
    .B(_03544_),
    .Y(_10903_));
 sky130_fd_sc_hd__nand2_4 _41441_ (.A(_10902_),
    .B(_10903_),
    .Y(_10904_));
 sky130_vsdinv _41442_ (.A(_10903_),
    .Y(_10905_));
 sky130_fd_sc_hd__nand3_4 _41443_ (.A(_10899_),
    .B(_10901_),
    .C(_10905_),
    .Y(_10906_));
 sky130_fd_sc_hd__and2_4 _41444_ (.A(_10904_),
    .B(_10906_),
    .X(_10907_));
 sky130_vsdinv _41445_ (.A(_10907_),
    .Y(_10908_));
 sky130_fd_sc_hd__nand2_4 _41446_ (.A(_10897_),
    .B(_10908_),
    .Y(_10909_));
 sky130_fd_sc_hd__nand3_4 _41447_ (.A(_10907_),
    .B(_10894_),
    .C(_10896_),
    .Y(_10910_));
 sky130_fd_sc_hd__nand2_4 _41448_ (.A(_10909_),
    .B(_10910_),
    .Y(_10911_));
 sky130_fd_sc_hd__nand2_4 _41449_ (.A(_10880_),
    .B(_10911_),
    .Y(_10912_));
 sky130_fd_sc_hd__nand3_4 _41450_ (.A(_10879_),
    .B(_10909_),
    .C(_10910_),
    .Y(_10913_));
 sky130_fd_sc_hd__nand2_4 _41451_ (.A(_10912_),
    .B(_10913_),
    .Y(_10914_));
 sky130_fd_sc_hd__a21boi_4 _41452_ (.A1(_10558_),
    .A2(_10546_),
    .B1_N(_10548_),
    .Y(_10915_));
 sky130_fd_sc_hd__nand2_4 _41453_ (.A(_10914_),
    .B(_10915_),
    .Y(_10916_));
 sky130_vsdinv _41454_ (.A(_10915_),
    .Y(_10917_));
 sky130_fd_sc_hd__nand3_4 _41455_ (.A(_10912_),
    .B(_10917_),
    .C(_10913_),
    .Y(_10918_));
 sky130_fd_sc_hd__nand2_4 _41456_ (.A(_10916_),
    .B(_10918_),
    .Y(_10919_));
 sky130_fd_sc_hd__buf_1 _41457_ (.A(_09756_),
    .X(_10920_));
 sky130_fd_sc_hd__nand2_4 _41458_ (.A(_06160_),
    .B(_10920_),
    .Y(_10921_));
 sky130_fd_sc_hd__buf_1 _41459_ (.A(_09760_),
    .X(_10922_));
 sky130_fd_sc_hd__nand2_4 _41460_ (.A(_06163_),
    .B(_10922_),
    .Y(_10923_));
 sky130_fd_sc_hd__nand2_4 _41461_ (.A(_10921_),
    .B(_10923_),
    .Y(_10924_));
 sky130_fd_sc_hd__buf_1 _41462_ (.A(_10476_),
    .X(_10925_));
 sky130_fd_sc_hd__nand4_4 _41463_ (.A(_06076_),
    .B(_06938_),
    .C(_09344_),
    .D(_10925_),
    .Y(_10926_));
 sky130_fd_sc_hd__buf_1 _41464_ (.A(_09346_),
    .X(_10927_));
 sky130_fd_sc_hd__nand2_4 _41465_ (.A(_06942_),
    .B(_10927_),
    .Y(_10928_));
 sky130_vsdinv _41466_ (.A(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__a21o_4 _41467_ (.A1(_10924_),
    .A2(_10926_),
    .B1(_10929_),
    .X(_10930_));
 sky130_fd_sc_hd__nand3_4 _41468_ (.A(_10924_),
    .B(_10926_),
    .C(_10929_),
    .Y(_10931_));
 sky130_fd_sc_hd__nand2_4 _41469_ (.A(_10930_),
    .B(_10931_),
    .Y(_10932_));
 sky130_fd_sc_hd__maj3_4 _41470_ (.A(_10510_),
    .B(_10500_),
    .C(_10503_),
    .X(_10933_));
 sky130_fd_sc_hd__nand2_4 _41471_ (.A(_10932_),
    .B(_10933_),
    .Y(_10934_));
 sky130_fd_sc_hd__nand2_4 _41472_ (.A(_10514_),
    .B(_10507_),
    .Y(_10935_));
 sky130_fd_sc_hd__nand3_4 _41473_ (.A(_10935_),
    .B(_10931_),
    .C(_10930_),
    .Y(_10936_));
 sky130_fd_sc_hd__nand2_4 _41474_ (.A(_10934_),
    .B(_10936_),
    .Y(_10937_));
 sky130_fd_sc_hd__a21boi_4 _41475_ (.A1(_10479_),
    .A2(_10484_),
    .B1_N(_10482_),
    .Y(_10938_));
 sky130_fd_sc_hd__nand2_4 _41476_ (.A(_10937_),
    .B(_10938_),
    .Y(_10939_));
 sky130_vsdinv _41477_ (.A(_10938_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand3_4 _41478_ (.A(_10934_),
    .B(_10936_),
    .C(_10940_),
    .Y(_10941_));
 sky130_fd_sc_hd__nand2_4 _41479_ (.A(_10939_),
    .B(_10941_),
    .Y(_10942_));
 sky130_fd_sc_hd__nand2_4 _41480_ (.A(_06055_),
    .B(_10324_),
    .Y(_10943_));
 sky130_fd_sc_hd__nand2_4 _41481_ (.A(_05915_),
    .B(_10322_),
    .Y(_10944_));
 sky130_fd_sc_hd__nand2_4 _41482_ (.A(_10943_),
    .B(_10944_),
    .Y(_10945_));
 sky130_fd_sc_hd__buf_1 _41483_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10946_));
 sky130_fd_sc_hd__buf_1 _41484_ (.A(_10498_),
    .X(_10947_));
 sky130_fd_sc_hd__nand4_4 _41485_ (.A(_06055_),
    .B(_07360_),
    .C(_10946_),
    .D(_10947_),
    .Y(_10948_));
 sky130_fd_sc_hd__nand2_4 _41486_ (.A(_10945_),
    .B(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__nand2_4 _41487_ (.A(_06222_),
    .B(_10035_),
    .Y(_10950_));
 sky130_fd_sc_hd__nand2_4 _41488_ (.A(_10949_),
    .B(_10950_),
    .Y(_10951_));
 sky130_vsdinv _41489_ (.A(_10950_),
    .Y(_10952_));
 sky130_fd_sc_hd__nand3_4 _41490_ (.A(_10945_),
    .B(_10948_),
    .C(_10952_),
    .Y(_10953_));
 sky130_fd_sc_hd__nand2_4 _41491_ (.A(_10951_),
    .B(_10953_),
    .Y(_10954_));
 sky130_fd_sc_hd__buf_1 _41492_ (.A(_10515_),
    .X(_10955_));
 sky130_fd_sc_hd__nand2_4 _41493_ (.A(_05885_),
    .B(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__o21ai_4 _41494_ (.A1(_03229_),
    .A2(_03629_),
    .B1(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__buf_1 _41495_ (.A(\pcpi_mul.rs2[31] ),
    .X(_10958_));
 sky130_fd_sc_hd__buf_4 _41496_ (.A(_10958_),
    .X(_10959_));
 sky130_fd_sc_hd__nand4_4 _41497_ (.A(_06634_),
    .B(_07048_),
    .C(_03620_),
    .D(_10959_),
    .Y(_10960_));
 sky130_fd_sc_hd__nand2_4 _41498_ (.A(_10957_),
    .B(_10960_),
    .Y(_10961_));
 sky130_fd_sc_hd__nand2_4 _41499_ (.A(_10954_),
    .B(_10961_),
    .Y(_10962_));
 sky130_vsdinv _41500_ (.A(_10961_),
    .Y(_10963_));
 sky130_fd_sc_hd__nand3_4 _41501_ (.A(_10963_),
    .B(_10953_),
    .C(_10951_),
    .Y(_10964_));
 sky130_fd_sc_hd__nand2_4 _41502_ (.A(_10962_),
    .B(_10964_),
    .Y(_10965_));
 sky130_fd_sc_hd__nand2_4 _41503_ (.A(_10965_),
    .B(_10521_),
    .Y(_10966_));
 sky130_vsdinv _41504_ (.A(_10521_),
    .Y(_10967_));
 sky130_fd_sc_hd__nand3_4 _41505_ (.A(_10967_),
    .B(_10964_),
    .C(_10962_),
    .Y(_10968_));
 sky130_fd_sc_hd__nand2_4 _41506_ (.A(_10966_),
    .B(_10968_),
    .Y(_10969_));
 sky130_fd_sc_hd__nand2_4 _41507_ (.A(_10942_),
    .B(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__nand4_4 _41508_ (.A(_10941_),
    .B(_10939_),
    .C(_10968_),
    .D(_10966_),
    .Y(_10971_));
 sky130_fd_sc_hd__nand2_4 _41509_ (.A(_10970_),
    .B(_10971_),
    .Y(_10972_));
 sky130_fd_sc_hd__nand2_4 _41510_ (.A(_10972_),
    .B(_10525_),
    .Y(_10973_));
 sky130_vsdinv _41511_ (.A(_10525_),
    .Y(_10974_));
 sky130_fd_sc_hd__nand3_4 _41512_ (.A(_10974_),
    .B(_10970_),
    .C(_10971_),
    .Y(_10975_));
 sky130_fd_sc_hd__nand2_4 _41513_ (.A(_10973_),
    .B(_10975_),
    .Y(_10976_));
 sky130_fd_sc_hd__nand2_4 _41514_ (.A(_10919_),
    .B(_10976_),
    .Y(_10977_));
 sky130_fd_sc_hd__nand4_4 _41515_ (.A(_10918_),
    .B(_10916_),
    .C(_10973_),
    .D(_10975_),
    .Y(_10978_));
 sky130_fd_sc_hd__nand2_4 _41516_ (.A(_10977_),
    .B(_10978_),
    .Y(_10979_));
 sky130_fd_sc_hd__nand2_4 _41517_ (.A(_10878_),
    .B(_10979_),
    .Y(_10980_));
 sky130_fd_sc_hd__nand2_4 _41518_ (.A(_10572_),
    .B(_10529_),
    .Y(_10981_));
 sky130_fd_sc_hd__nand3_4 _41519_ (.A(_10981_),
    .B(_10978_),
    .C(_10977_),
    .Y(_10982_));
 sky130_fd_sc_hd__nand2_4 _41520_ (.A(_10980_),
    .B(_10982_),
    .Y(_10983_));
 sky130_fd_sc_hd__a21boi_4 _41521_ (.A1(_10552_),
    .A2(_10555_),
    .B1_N(_10553_),
    .Y(_10984_));
 sky130_vsdinv _41522_ (.A(_10984_),
    .Y(_10985_));
 sky130_fd_sc_hd__nand2_4 _41523_ (.A(_03314_),
    .B(_07922_),
    .Y(_10986_));
 sky130_fd_sc_hd__nand2_4 _41524_ (.A(_07157_),
    .B(_07713_),
    .Y(_10987_));
 sky130_fd_sc_hd__nand2_4 _41525_ (.A(_10986_),
    .B(_10987_),
    .Y(_10988_));
 sky130_fd_sc_hd__buf_1 _41526_ (.A(_07421_),
    .X(_10989_));
 sky130_fd_sc_hd__buf_1 _41527_ (.A(_08795_),
    .X(_10990_));
 sky130_fd_sc_hd__nand4_4 _41528_ (.A(_10989_),
    .B(_03318_),
    .C(_10990_),
    .D(_08125_),
    .Y(_10991_));
 sky130_fd_sc_hd__nand2_4 _41529_ (.A(_07620_),
    .B(_07562_),
    .Y(_10992_));
 sky130_vsdinv _41530_ (.A(_10992_),
    .Y(_10993_));
 sky130_fd_sc_hd__nand3_4 _41531_ (.A(_10988_),
    .B(_10991_),
    .C(_10993_),
    .Y(_10994_));
 sky130_fd_sc_hd__nand2_4 _41532_ (.A(_10988_),
    .B(_10991_),
    .Y(_10995_));
 sky130_fd_sc_hd__nand2_4 _41533_ (.A(_10995_),
    .B(_10992_),
    .Y(_10996_));
 sky130_fd_sc_hd__nand3_4 _41534_ (.A(_10985_),
    .B(_10994_),
    .C(_10996_),
    .Y(_10997_));
 sky130_fd_sc_hd__nand2_4 _41535_ (.A(_10996_),
    .B(_10994_),
    .Y(_10998_));
 sky130_fd_sc_hd__nand2_4 _41536_ (.A(_10998_),
    .B(_10984_),
    .Y(_10999_));
 sky130_fd_sc_hd__a21boi_4 _41537_ (.A1(_10583_),
    .A2(_10587_),
    .B1_N(_10585_),
    .Y(_11000_));
 sky130_vsdinv _41538_ (.A(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__a21o_4 _41539_ (.A1(_10997_),
    .A2(_10999_),
    .B1(_11001_),
    .X(_11002_));
 sky130_fd_sc_hd__nand3_4 _41540_ (.A(_10997_),
    .B(_10999_),
    .C(_11001_),
    .Y(_11003_));
 sky130_fd_sc_hd__nand2_4 _41541_ (.A(_11002_),
    .B(_11003_),
    .Y(_11004_));
 sky130_fd_sc_hd__a21boi_4 _41542_ (.A1(_10593_),
    .A2(_10597_),
    .B1_N(_10591_),
    .Y(_11005_));
 sky130_fd_sc_hd__nand2_4 _41543_ (.A(_11004_),
    .B(_11005_),
    .Y(_11006_));
 sky130_vsdinv _41544_ (.A(_11005_),
    .Y(_11007_));
 sky130_fd_sc_hd__nand3_4 _41545_ (.A(_11007_),
    .B(_11003_),
    .C(_11002_),
    .Y(_11008_));
 sky130_fd_sc_hd__nand2_4 _41546_ (.A(_11006_),
    .B(_11008_),
    .Y(_11009_));
 sky130_fd_sc_hd__buf_1 _41547_ (.A(_07443_),
    .X(_11010_));
 sky130_fd_sc_hd__nand2_4 _41548_ (.A(_11010_),
    .B(_07741_),
    .Y(_11011_));
 sky130_fd_sc_hd__nand2_4 _41549_ (.A(_10212_),
    .B(_07189_),
    .Y(_11012_));
 sky130_fd_sc_hd__nand2_4 _41550_ (.A(_11011_),
    .B(_11012_),
    .Y(_11013_));
 sky130_fd_sc_hd__buf_1 _41551_ (.A(_09038_),
    .X(_11014_));
 sky130_fd_sc_hd__buf_1 _41552_ (.A(_08510_),
    .X(_11015_));
 sky130_fd_sc_hd__buf_1 _41553_ (.A(_07356_),
    .X(_11016_));
 sky130_fd_sc_hd__buf_1 _41554_ (.A(_07734_),
    .X(_11017_));
 sky130_fd_sc_hd__nand4_4 _41555_ (.A(_11014_),
    .B(_11015_),
    .C(_11016_),
    .D(_11017_),
    .Y(_11018_));
 sky130_fd_sc_hd__buf_1 _41556_ (.A(_03341_),
    .X(_11019_));
 sky130_fd_sc_hd__nand2_4 _41557_ (.A(_11019_),
    .B(_07197_),
    .Y(_11020_));
 sky130_fd_sc_hd__a21bo_4 _41558_ (.A1(_11013_),
    .A2(_11018_),
    .B1_N(_11020_),
    .X(_11021_));
 sky130_fd_sc_hd__buf_1 _41559_ (.A(_03342_),
    .X(_11022_));
 sky130_fd_sc_hd__buf_1 _41560_ (.A(_06881_),
    .X(_11023_));
 sky130_fd_sc_hd__nand4_4 _41561_ (.A(_11022_),
    .B(_11013_),
    .C(_11018_),
    .D(_11023_),
    .Y(_11024_));
 sky130_fd_sc_hd__a21boi_4 _41562_ (.A1(_10608_),
    .A2(_10611_),
    .B1_N(_10609_),
    .Y(_11025_));
 sky130_vsdinv _41563_ (.A(_11025_),
    .Y(_11026_));
 sky130_fd_sc_hd__a21o_4 _41564_ (.A1(_11021_),
    .A2(_11024_),
    .B1(_11026_),
    .X(_11027_));
 sky130_fd_sc_hd__nand3_4 _41565_ (.A(_11026_),
    .B(_11021_),
    .C(_11024_),
    .Y(_11028_));
 sky130_fd_sc_hd__nand2_4 _41566_ (.A(_11027_),
    .B(_11028_),
    .Y(_11029_));
 sky130_fd_sc_hd__buf_1 _41567_ (.A(_03353_),
    .X(_11030_));
 sky130_fd_sc_hd__nand2_4 _41568_ (.A(_11030_),
    .B(_06887_),
    .Y(_11031_));
 sky130_fd_sc_hd__o21ai_4 _41569_ (.A1(_03347_),
    .A2(_03506_),
    .B1(_11031_),
    .Y(_11032_));
 sky130_fd_sc_hd__buf_1 _41570_ (.A(_09074_),
    .X(_11033_));
 sky130_fd_sc_hd__buf_1 _41571_ (.A(_08314_),
    .X(_11034_));
 sky130_fd_sc_hd__nand4_4 _41572_ (.A(_11033_),
    .B(_11034_),
    .C(_06506_),
    .D(_06637_),
    .Y(_11035_));
 sky130_fd_sc_hd__nand2_4 _41573_ (.A(_09830_),
    .B(_06751_),
    .Y(_11036_));
 sky130_vsdinv _41574_ (.A(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__a21oi_4 _41575_ (.A1(_11032_),
    .A2(_11035_),
    .B1(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__nand3_4 _41576_ (.A(_11032_),
    .B(_11035_),
    .C(_11037_),
    .Y(_11039_));
 sky130_vsdinv _41577_ (.A(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__nor2_4 _41578_ (.A(_11038_),
    .B(_11040_),
    .Y(_11041_));
 sky130_vsdinv _41579_ (.A(_11041_),
    .Y(_11042_));
 sky130_fd_sc_hd__nand2_4 _41580_ (.A(_11029_),
    .B(_11042_),
    .Y(_11043_));
 sky130_fd_sc_hd__nand3_4 _41581_ (.A(_11027_),
    .B(_11041_),
    .C(_11028_),
    .Y(_11044_));
 sky130_fd_sc_hd__and2_4 _41582_ (.A(_11043_),
    .B(_11044_),
    .X(_11045_));
 sky130_vsdinv _41583_ (.A(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__nand2_4 _41584_ (.A(_11009_),
    .B(_11046_),
    .Y(_11047_));
 sky130_fd_sc_hd__nand3_4 _41585_ (.A(_11045_),
    .B(_11006_),
    .C(_11008_),
    .Y(_11048_));
 sky130_fd_sc_hd__nand2_4 _41586_ (.A(_11047_),
    .B(_11048_),
    .Y(_11049_));
 sky130_fd_sc_hd__a21boi_4 _41587_ (.A1(_10568_),
    .A2(_10564_),
    .B1_N(_10562_),
    .Y(_11050_));
 sky130_fd_sc_hd__nand2_4 _41588_ (.A(_11049_),
    .B(_11050_),
    .Y(_11051_));
 sky130_vsdinv _41589_ (.A(_11050_),
    .Y(_11052_));
 sky130_fd_sc_hd__nand3_4 _41590_ (.A(_11052_),
    .B(_11048_),
    .C(_11047_),
    .Y(_11053_));
 sky130_fd_sc_hd__nand2_4 _41591_ (.A(_11051_),
    .B(_11053_),
    .Y(_11054_));
 sky130_fd_sc_hd__a21boi_4 _41592_ (.A1(_10635_),
    .A2(_10601_),
    .B1_N(_10603_),
    .Y(_11055_));
 sky130_fd_sc_hd__nand2_4 _41593_ (.A(_11054_),
    .B(_11055_),
    .Y(_11056_));
 sky130_vsdinv _41594_ (.A(_11055_),
    .Y(_11057_));
 sky130_fd_sc_hd__nand3_4 _41595_ (.A(_11051_),
    .B(_11053_),
    .C(_11057_),
    .Y(_11058_));
 sky130_fd_sc_hd__nand2_4 _41596_ (.A(_11056_),
    .B(_11058_),
    .Y(_11059_));
 sky130_fd_sc_hd__nand2_4 _41597_ (.A(_10983_),
    .B(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__nand4_4 _41598_ (.A(_11058_),
    .B(_10980_),
    .C(_10982_),
    .D(_11056_),
    .Y(_11061_));
 sky130_fd_sc_hd__nand2_4 _41599_ (.A(_11060_),
    .B(_11061_),
    .Y(_11062_));
 sky130_fd_sc_hd__a21oi_4 _41600_ (.A1(_10572_),
    .A2(_10571_),
    .B1(_10575_),
    .Y(_11063_));
 sky130_fd_sc_hd__o21a_4 _41601_ (.A1(_11063_),
    .A2(_10650_),
    .B1(_10576_),
    .X(_11064_));
 sky130_fd_sc_hd__nand2_4 _41602_ (.A(_11062_),
    .B(_11064_),
    .Y(_11065_));
 sky130_fd_sc_hd__o21ai_4 _41603_ (.A1(_11063_),
    .A2(_10650_),
    .B1(_10576_),
    .Y(_11066_));
 sky130_fd_sc_hd__nand3_4 _41604_ (.A(_11066_),
    .B(_11061_),
    .C(_11060_),
    .Y(_11067_));
 sky130_fd_sc_hd__nand2_4 _41605_ (.A(_11065_),
    .B(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__nand2_4 _41606_ (.A(_10877_),
    .B(_11068_),
    .Y(_11069_));
 sky130_fd_sc_hd__nand4_4 _41607_ (.A(_10876_),
    .B(_10874_),
    .C(_11065_),
    .D(_11067_),
    .Y(_11070_));
 sky130_fd_sc_hd__nand2_4 _41608_ (.A(_11069_),
    .B(_11070_),
    .Y(_11071_));
 sky130_fd_sc_hd__a21oi_4 _41609_ (.A1(_10651_),
    .A2(_10652_),
    .B1(_10657_),
    .Y(_11072_));
 sky130_fd_sc_hd__o21a_4 _41610_ (.A1(_11072_),
    .A2(_10749_),
    .B1(_10658_),
    .X(_11073_));
 sky130_fd_sc_hd__nand2_4 _41611_ (.A(_11071_),
    .B(_11073_),
    .Y(_11074_));
 sky130_fd_sc_hd__o21ai_4 _41612_ (.A1(_11072_),
    .A2(_10749_),
    .B1(_10658_),
    .Y(_11075_));
 sky130_fd_sc_hd__nand3_4 _41613_ (.A(_11075_),
    .B(_11070_),
    .C(_11069_),
    .Y(_11076_));
 sky130_fd_sc_hd__nand2_4 _41614_ (.A(_11074_),
    .B(_11076_),
    .Y(_11077_));
 sky130_fd_sc_hd__a21boi_4 _41615_ (.A1(_10731_),
    .A2(_10729_),
    .B1_N(_10727_),
    .Y(_11078_));
 sky130_fd_sc_hd__a21boi_4 _41616_ (.A1(_10741_),
    .A2(_10747_),
    .B1_N(_10743_),
    .Y(_11079_));
 sky130_fd_sc_hd__xnor2_4 _41617_ (.A(_11078_),
    .B(_11079_),
    .Y(_11080_));
 sky130_fd_sc_hd__nand2_4 _41618_ (.A(_11077_),
    .B(_11080_),
    .Y(_11081_));
 sky130_vsdinv _41619_ (.A(_11080_),
    .Y(_11082_));
 sky130_fd_sc_hd__nand3_4 _41620_ (.A(_11074_),
    .B(_11076_),
    .C(_11082_),
    .Y(_11083_));
 sky130_fd_sc_hd__nand2_4 _41621_ (.A(_11081_),
    .B(_11083_),
    .Y(_11084_));
 sky130_fd_sc_hd__a21boi_4 _41622_ (.A1(_10753_),
    .A2(_10761_),
    .B1_N(_10755_),
    .Y(_11085_));
 sky130_fd_sc_hd__nand2_4 _41623_ (.A(_11084_),
    .B(_11085_),
    .Y(_11086_));
 sky130_fd_sc_hd__nand2_4 _41624_ (.A(_10762_),
    .B(_10755_),
    .Y(_11087_));
 sky130_fd_sc_hd__nand3_4 _41625_ (.A(_11087_),
    .B(_11083_),
    .C(_11081_),
    .Y(_11088_));
 sky130_fd_sc_hd__nand2_4 _41626_ (.A(_11086_),
    .B(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__a21oi_4 _41627_ (.A1(_10440_),
    .A2(_10435_),
    .B1(_10757_),
    .Y(_11090_));
 sky130_vsdinv _41628_ (.A(_11090_),
    .Y(_11091_));
 sky130_fd_sc_hd__nand2_4 _41629_ (.A(_11089_),
    .B(_11091_),
    .Y(_11092_));
 sky130_fd_sc_hd__nand3_4 _41630_ (.A(_11086_),
    .B(_11088_),
    .C(_11090_),
    .Y(_11093_));
 sky130_fd_sc_hd__a21oi_4 _41631_ (.A1(_10760_),
    .A2(_10762_),
    .B1(_10764_),
    .Y(_11094_));
 sky130_fd_sc_hd__o21ai_4 _41632_ (.A1(_10770_),
    .A2(_11094_),
    .B1(_10767_),
    .Y(_11095_));
 sky130_fd_sc_hd__a21oi_4 _41633_ (.A1(_11092_),
    .A2(_11093_),
    .B1(_11095_),
    .Y(_11096_));
 sky130_fd_sc_hd__nand3_4 _41634_ (.A(_11092_),
    .B(_11095_),
    .C(_11093_),
    .Y(_11097_));
 sky130_vsdinv _41635_ (.A(_11097_),
    .Y(_11098_));
 sky130_fd_sc_hd__nor2_4 _41636_ (.A(_11096_),
    .B(_11098_),
    .Y(_11099_));
 sky130_fd_sc_hd__o21ai_4 _41637_ (.A1(_10780_),
    .A2(_10782_),
    .B1(_10777_),
    .Y(_11100_));
 sky130_fd_sc_hd__xor2_4 _41638_ (.A(_11099_),
    .B(_11100_),
    .X(_01436_));
 sky130_fd_sc_hd__buf_1 _41639_ (.A(_03632_),
    .X(_11101_));
 sky130_fd_sc_hd__buf_1 _41640_ (.A(_03627_),
    .X(_11102_));
 sky130_fd_sc_hd__nand2_4 _41641_ (.A(_06050_),
    .B(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__o21ai_4 _41642_ (.A1(_05961_),
    .A2(_11101_),
    .B1(_11103_),
    .Y(_11104_));
 sky130_fd_sc_hd__buf_1 _41643_ (.A(_10958_),
    .X(_11105_));
 sky130_fd_sc_hd__buf_1 _41644_ (.A(\pcpi_mul.rs2[32] ),
    .X(_11106_));
 sky130_fd_sc_hd__buf_1 _41645_ (.A(_11106_),
    .X(_11107_));
 sky130_fd_sc_hd__nand4_4 _41646_ (.A(_03229_),
    .B(_05987_),
    .C(_11105_),
    .D(_11107_),
    .Y(_11108_));
 sky130_fd_sc_hd__nand2_4 _41647_ (.A(_11104_),
    .B(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__nand2_4 _41648_ (.A(_06055_),
    .B(_10516_),
    .Y(_11110_));
 sky130_fd_sc_hd__nand2_4 _41649_ (.A(_11109_),
    .B(_11110_),
    .Y(_11111_));
 sky130_vsdinv _41650_ (.A(_11110_),
    .Y(_11112_));
 sky130_fd_sc_hd__nand3_4 _41651_ (.A(_11104_),
    .B(_11112_),
    .C(_11108_),
    .Y(_11113_));
 sky130_fd_sc_hd__nand2_4 _41652_ (.A(_11111_),
    .B(_11113_),
    .Y(_11114_));
 sky130_fd_sc_hd__nand2_4 _41653_ (.A(_11114_),
    .B(_10960_),
    .Y(_11115_));
 sky130_vsdinv _41654_ (.A(_10960_),
    .Y(_11116_));
 sky130_fd_sc_hd__nand3_4 _41655_ (.A(_11111_),
    .B(_11116_),
    .C(_11113_),
    .Y(_11117_));
 sky130_fd_sc_hd__nand2_4 _41656_ (.A(_11115_),
    .B(_11117_),
    .Y(_11118_));
 sky130_fd_sc_hd__buf_1 _41657_ (.A(_10498_),
    .X(_11119_));
 sky130_fd_sc_hd__nand2_4 _41658_ (.A(_06384_),
    .B(_11119_),
    .Y(_11120_));
 sky130_fd_sc_hd__buf_1 _41659_ (.A(_10501_),
    .X(_11121_));
 sky130_fd_sc_hd__nand2_4 _41660_ (.A(_10480_),
    .B(_11121_),
    .Y(_11122_));
 sky130_fd_sc_hd__nand2_4 _41661_ (.A(_11120_),
    .B(_11122_),
    .Y(_11123_));
 sky130_fd_sc_hd__nand4_4 _41662_ (.A(_07196_),
    .B(_07740_),
    .C(_10505_),
    .D(_10506_),
    .Y(_11124_));
 sky130_fd_sc_hd__buf_1 _41663_ (.A(_10035_),
    .X(_11125_));
 sky130_fd_sc_hd__nand2_4 _41664_ (.A(_06160_),
    .B(_11125_),
    .Y(_11126_));
 sky130_vsdinv _41665_ (.A(_11126_),
    .Y(_11127_));
 sky130_fd_sc_hd__a21o_4 _41666_ (.A1(_11123_),
    .A2(_11124_),
    .B1(_11127_),
    .X(_11128_));
 sky130_fd_sc_hd__nand3_4 _41667_ (.A(_11123_),
    .B(_11124_),
    .C(_11127_),
    .Y(_11129_));
 sky130_fd_sc_hd__and2_4 _41668_ (.A(_11128_),
    .B(_11129_),
    .X(_11130_));
 sky130_vsdinv _41669_ (.A(_11130_),
    .Y(_11131_));
 sky130_fd_sc_hd__nand2_4 _41670_ (.A(_11118_),
    .B(_11131_),
    .Y(_11132_));
 sky130_fd_sc_hd__nand3_4 _41671_ (.A(_11115_),
    .B(_11130_),
    .C(_11117_),
    .Y(_11133_));
 sky130_fd_sc_hd__nand2_4 _41672_ (.A(_11132_),
    .B(_11133_),
    .Y(_11134_));
 sky130_fd_sc_hd__nand2_4 _41673_ (.A(_11134_),
    .B(_10964_),
    .Y(_11135_));
 sky130_vsdinv _41674_ (.A(_10964_),
    .Y(_11136_));
 sky130_fd_sc_hd__nand3_4 _41675_ (.A(_11132_),
    .B(_11133_),
    .C(_11136_),
    .Y(_11137_));
 sky130_fd_sc_hd__nand2_4 _41676_ (.A(_11135_),
    .B(_11137_),
    .Y(_11138_));
 sky130_fd_sc_hd__nand2_4 _41677_ (.A(_07346_),
    .B(_10920_),
    .Y(_11139_));
 sky130_fd_sc_hd__nand2_4 _41678_ (.A(_08381_),
    .B(_10922_),
    .Y(_11140_));
 sky130_fd_sc_hd__nand2_4 _41679_ (.A(_11139_),
    .B(_11140_),
    .Y(_11141_));
 sky130_fd_sc_hd__buf_1 _41680_ (.A(_10476_),
    .X(_11142_));
 sky130_fd_sc_hd__nand4_4 _41681_ (.A(_06170_),
    .B(_06545_),
    .C(_09344_),
    .D(_11142_),
    .Y(_11143_));
 sky130_fd_sc_hd__nand2_4 _41682_ (.A(_07959_),
    .B(_10927_),
    .Y(_11144_));
 sky130_vsdinv _41683_ (.A(_11144_),
    .Y(_11145_));
 sky130_fd_sc_hd__a21o_4 _41684_ (.A1(_11141_),
    .A2(_11143_),
    .B1(_11145_),
    .X(_11146_));
 sky130_fd_sc_hd__nand3_4 _41685_ (.A(_11141_),
    .B(_11143_),
    .C(_11145_),
    .Y(_11147_));
 sky130_fd_sc_hd__nand2_4 _41686_ (.A(_11146_),
    .B(_11147_),
    .Y(_11148_));
 sky130_fd_sc_hd__a21boi_4 _41687_ (.A1(_10945_),
    .A2(_10952_),
    .B1_N(_10948_),
    .Y(_11149_));
 sky130_fd_sc_hd__nand2_4 _41688_ (.A(_11148_),
    .B(_11149_),
    .Y(_11150_));
 sky130_vsdinv _41689_ (.A(_11149_),
    .Y(_11151_));
 sky130_fd_sc_hd__nand3_4 _41690_ (.A(_11151_),
    .B(_11146_),
    .C(_11147_),
    .Y(_11152_));
 sky130_fd_sc_hd__a21boi_4 _41691_ (.A1(_10924_),
    .A2(_10929_),
    .B1_N(_10926_),
    .Y(_11153_));
 sky130_vsdinv _41692_ (.A(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__a21o_4 _41693_ (.A1(_11150_),
    .A2(_11152_),
    .B1(_11154_),
    .X(_11155_));
 sky130_fd_sc_hd__nand3_4 _41694_ (.A(_11150_),
    .B(_11152_),
    .C(_11154_),
    .Y(_11156_));
 sky130_fd_sc_hd__nand2_4 _41695_ (.A(_11155_),
    .B(_11156_),
    .Y(_11157_));
 sky130_fd_sc_hd__nand2_4 _41696_ (.A(_11138_),
    .B(_11157_),
    .Y(_11158_));
 sky130_vsdinv _41697_ (.A(_11157_),
    .Y(_11159_));
 sky130_fd_sc_hd__nand3_4 _41698_ (.A(_11135_),
    .B(_11159_),
    .C(_11137_),
    .Y(_11160_));
 sky130_fd_sc_hd__nand2_4 _41699_ (.A(_11158_),
    .B(_11160_),
    .Y(_11161_));
 sky130_fd_sc_hd__o21a_4 _41700_ (.A1(_10969_),
    .A2(_10942_),
    .B1(_10968_),
    .X(_11162_));
 sky130_fd_sc_hd__nand2_4 _41701_ (.A(_11161_),
    .B(_11162_),
    .Y(_11163_));
 sky130_vsdinv _41702_ (.A(_11162_),
    .Y(_11164_));
 sky130_fd_sc_hd__nand3_4 _41703_ (.A(_11158_),
    .B(_11164_),
    .C(_11160_),
    .Y(_11165_));
 sky130_fd_sc_hd__nand2_4 _41704_ (.A(_11163_),
    .B(_11165_),
    .Y(_11166_));
 sky130_fd_sc_hd__buf_1 _41705_ (.A(_10270_),
    .X(_11167_));
 sky130_fd_sc_hd__nand2_4 _41706_ (.A(_06447_),
    .B(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__buf_1 _41707_ (.A(_10272_),
    .X(_11169_));
 sky130_fd_sc_hd__nand2_4 _41708_ (.A(_06833_),
    .B(_11169_),
    .Y(_11170_));
 sky130_fd_sc_hd__nand2_4 _41709_ (.A(_11168_),
    .B(_11170_),
    .Y(_11171_));
 sky130_fd_sc_hd__buf_1 _41710_ (.A(_08631_),
    .X(_11172_));
 sky130_fd_sc_hd__buf_1 _41711_ (.A(_03576_),
    .X(_11173_));
 sky130_fd_sc_hd__nand4_4 _41712_ (.A(_06452_),
    .B(_06456_),
    .C(_11172_),
    .D(_11173_),
    .Y(_11174_));
 sky130_fd_sc_hd__buf_1 _41713_ (.A(_03563_),
    .X(_11175_));
 sky130_fd_sc_hd__nand2_4 _41714_ (.A(_06983_),
    .B(_11175_),
    .Y(_11176_));
 sky130_fd_sc_hd__a21bo_4 _41715_ (.A1(_11171_),
    .A2(_11174_),
    .B1_N(_11176_),
    .X(_11177_));
 sky130_fd_sc_hd__nand4_4 _41716_ (.A(_06572_),
    .B(_11171_),
    .C(_11174_),
    .D(_03565_),
    .Y(_11178_));
 sky130_fd_sc_hd__a21boi_4 _41717_ (.A1(_10883_),
    .A2(_10889_),
    .B1_N(_10886_),
    .Y(_11179_));
 sky130_vsdinv _41718_ (.A(_11179_),
    .Y(_11180_));
 sky130_fd_sc_hd__a21o_4 _41719_ (.A1(_11177_),
    .A2(_11178_),
    .B1(_11180_),
    .X(_11181_));
 sky130_fd_sc_hd__nand3_4 _41720_ (.A(_11180_),
    .B(_11177_),
    .C(_11178_),
    .Y(_11182_));
 sky130_fd_sc_hd__nand2_4 _41721_ (.A(_07605_),
    .B(_03545_),
    .Y(_11183_));
 sky130_fd_sc_hd__nand2_4 _41722_ (.A(_07000_),
    .B(_07977_),
    .Y(_11184_));
 sky130_fd_sc_hd__o21ai_4 _41723_ (.A1(_03304_),
    .A2(_03558_),
    .B1(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__buf_1 _41724_ (.A(_09416_),
    .X(_11186_));
 sky130_fd_sc_hd__buf_1 _41725_ (.A(_09415_),
    .X(_11187_));
 sky130_fd_sc_hd__nand4_4 _41726_ (.A(_06713_),
    .B(_07151_),
    .C(_11186_),
    .D(_11187_),
    .Y(_11188_));
 sky130_fd_sc_hd__nand2_4 _41727_ (.A(_11185_),
    .B(_11188_),
    .Y(_11189_));
 sky130_fd_sc_hd__xor2_4 _41728_ (.A(_11183_),
    .B(_11189_),
    .X(_11190_));
 sky130_fd_sc_hd__a21oi_4 _41729_ (.A1(_11181_),
    .A2(_11182_),
    .B1(_11190_),
    .Y(_11191_));
 sky130_fd_sc_hd__nand3_4 _41730_ (.A(_11190_),
    .B(_11181_),
    .C(_11182_),
    .Y(_11192_));
 sky130_vsdinv _41731_ (.A(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__a21boi_4 _41732_ (.A1(_10934_),
    .A2(_10940_),
    .B1_N(_10936_),
    .Y(_11194_));
 sky130_fd_sc_hd__o21ai_4 _41733_ (.A1(_11191_),
    .A2(_11193_),
    .B1(_11194_),
    .Y(_11195_));
 sky130_vsdinv _41734_ (.A(_11191_),
    .Y(_11196_));
 sky130_vsdinv _41735_ (.A(_11194_),
    .Y(_11197_));
 sky130_fd_sc_hd__nand3_4 _41736_ (.A(_11196_),
    .B(_11197_),
    .C(_11192_),
    .Y(_11198_));
 sky130_fd_sc_hd__a21boi_4 _41737_ (.A1(_10907_),
    .A2(_10894_),
    .B1_N(_10896_),
    .Y(_11199_));
 sky130_vsdinv _41738_ (.A(_11199_),
    .Y(_11200_));
 sky130_fd_sc_hd__a21o_4 _41739_ (.A1(_11195_),
    .A2(_11198_),
    .B1(_11200_),
    .X(_11201_));
 sky130_fd_sc_hd__nand3_4 _41740_ (.A(_11195_),
    .B(_11198_),
    .C(_11200_),
    .Y(_11202_));
 sky130_fd_sc_hd__nand2_4 _41741_ (.A(_11201_),
    .B(_11202_),
    .Y(_11203_));
 sky130_fd_sc_hd__nand2_4 _41742_ (.A(_11166_),
    .B(_11203_),
    .Y(_11204_));
 sky130_fd_sc_hd__nand4_4 _41743_ (.A(_11202_),
    .B(_11163_),
    .C(_11201_),
    .D(_11165_),
    .Y(_11205_));
 sky130_fd_sc_hd__nand2_4 _41744_ (.A(_11204_),
    .B(_11205_),
    .Y(_11206_));
 sky130_fd_sc_hd__o21a_4 _41745_ (.A1(_10976_),
    .A2(_10919_),
    .B1(_10975_),
    .X(_11207_));
 sky130_fd_sc_hd__nand2_4 _41746_ (.A(_11206_),
    .B(_11207_),
    .Y(_11208_));
 sky130_vsdinv _41747_ (.A(_11207_),
    .Y(_11209_));
 sky130_fd_sc_hd__nand3_4 _41748_ (.A(_11209_),
    .B(_11204_),
    .C(_11205_),
    .Y(_11210_));
 sky130_fd_sc_hd__nand2_4 _41749_ (.A(_11208_),
    .B(_11210_),
    .Y(_11211_));
 sky130_fd_sc_hd__nand2_4 _41750_ (.A(_08966_),
    .B(_08566_),
    .Y(_11212_));
 sky130_fd_sc_hd__nand2_4 _41751_ (.A(_09037_),
    .B(_07553_),
    .Y(_11213_));
 sky130_fd_sc_hd__nand2_4 _41752_ (.A(_11212_),
    .B(_11213_),
    .Y(_11214_));
 sky130_fd_sc_hd__nand4_4 _41753_ (.A(_10198_),
    .B(_07624_),
    .C(_08572_),
    .D(_07710_),
    .Y(_11215_));
 sky130_fd_sc_hd__nand2_4 _41754_ (.A(_03332_),
    .B(_07562_),
    .Y(_11216_));
 sky130_vsdinv _41755_ (.A(_11216_),
    .Y(_11217_));
 sky130_fd_sc_hd__a21o_4 _41756_ (.A1(_11214_),
    .A2(_11215_),
    .B1(_11217_),
    .X(_11218_));
 sky130_fd_sc_hd__nand3_4 _41757_ (.A(_11214_),
    .B(_11215_),
    .C(_11217_),
    .Y(_11219_));
 sky130_fd_sc_hd__nand2_4 _41758_ (.A(_11218_),
    .B(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__a21o_4 _41759_ (.A1(_10901_),
    .A2(_10906_),
    .B1(_11220_),
    .X(_11221_));
 sky130_fd_sc_hd__a21boi_4 _41760_ (.A1(_10899_),
    .A2(_10905_),
    .B1_N(_10901_),
    .Y(_11222_));
 sky130_fd_sc_hd__nand2_4 _41761_ (.A(_11220_),
    .B(_11222_),
    .Y(_11223_));
 sky130_fd_sc_hd__nand2_4 _41762_ (.A(_11221_),
    .B(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__a21boi_4 _41763_ (.A1(_10988_),
    .A2(_10993_),
    .B1_N(_10991_),
    .Y(_11225_));
 sky130_fd_sc_hd__nand2_4 _41764_ (.A(_11224_),
    .B(_11225_),
    .Y(_11226_));
 sky130_vsdinv _41765_ (.A(_11225_),
    .Y(_11227_));
 sky130_fd_sc_hd__nand3_4 _41766_ (.A(_11221_),
    .B(_11227_),
    .C(_11223_),
    .Y(_11228_));
 sky130_fd_sc_hd__nand2_4 _41767_ (.A(_11226_),
    .B(_11228_),
    .Y(_11229_));
 sky130_fd_sc_hd__a21boi_4 _41768_ (.A1(_11001_),
    .A2(_10999_),
    .B1_N(_10997_),
    .Y(_11230_));
 sky130_fd_sc_hd__nand2_4 _41769_ (.A(_11229_),
    .B(_11230_),
    .Y(_11231_));
 sky130_vsdinv _41770_ (.A(_11230_),
    .Y(_11232_));
 sky130_fd_sc_hd__nand3_4 _41771_ (.A(_11226_),
    .B(_11232_),
    .C(_11228_),
    .Y(_11233_));
 sky130_fd_sc_hd__nand2_4 _41772_ (.A(_11231_),
    .B(_11233_),
    .Y(_11234_));
 sky130_fd_sc_hd__maj3_4 _41773_ (.A(_11011_),
    .B(_11020_),
    .C(_11012_),
    .X(_11235_));
 sky130_fd_sc_hd__nand2_4 _41774_ (.A(_07871_),
    .B(_07362_),
    .Y(_11236_));
 sky130_fd_sc_hd__nand2_4 _41775_ (.A(_09070_),
    .B(_07737_),
    .Y(_11237_));
 sky130_fd_sc_hd__nand2_4 _41776_ (.A(_11236_),
    .B(_11237_),
    .Y(_11238_));
 sky130_fd_sc_hd__nand4_4 _41777_ (.A(_03337_),
    .B(_08052_),
    .C(_07518_),
    .D(_07187_),
    .Y(_11239_));
 sky130_fd_sc_hd__nand2_4 _41778_ (.A(_08523_),
    .B(_07744_),
    .Y(_11240_));
 sky130_fd_sc_hd__a21bo_4 _41779_ (.A1(_11238_),
    .A2(_11239_),
    .B1_N(_11240_),
    .X(_11241_));
 sky130_fd_sc_hd__buf_1 _41780_ (.A(_08055_),
    .X(_11242_));
 sky130_fd_sc_hd__buf_1 _41781_ (.A(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__nand4_4 _41782_ (.A(_11243_),
    .B(_11238_),
    .C(_11239_),
    .D(_07747_),
    .Y(_11244_));
 sky130_fd_sc_hd__nand2_4 _41783_ (.A(_11241_),
    .B(_11244_),
    .Y(_11245_));
 sky130_fd_sc_hd__nor2_4 _41784_ (.A(_11235_),
    .B(_11245_),
    .Y(_11246_));
 sky130_fd_sc_hd__a21boi_4 _41785_ (.A1(_11244_),
    .A2(_11241_),
    .B1_N(_11235_),
    .Y(_11247_));
 sky130_fd_sc_hd__nor2_4 _41786_ (.A(_11246_),
    .B(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__buf_1 _41787_ (.A(_08758_),
    .X(_11249_));
 sky130_fd_sc_hd__nand2_4 _41788_ (.A(_11249_),
    .B(_07205_),
    .Y(_11250_));
 sky130_fd_sc_hd__nand2_4 _41789_ (.A(_09087_),
    .B(_07541_),
    .Y(_11251_));
 sky130_fd_sc_hd__o21ai_4 _41790_ (.A1(_03354_),
    .A2(_03505_),
    .B1(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__nand4_4 _41791_ (.A(_08753_),
    .B(_10664_),
    .C(_03501_),
    .D(_06748_),
    .Y(_11253_));
 sky130_fd_sc_hd__nand2_4 _41792_ (.A(_11252_),
    .B(_11253_),
    .Y(_11254_));
 sky130_fd_sc_hd__xor2_4 _41793_ (.A(_11250_),
    .B(_11254_),
    .X(_11255_));
 sky130_fd_sc_hd__nand2_4 _41794_ (.A(_11248_),
    .B(_11255_),
    .Y(_11256_));
 sky130_vsdinv _41795_ (.A(_11255_),
    .Y(_11257_));
 sky130_fd_sc_hd__o21ai_4 _41796_ (.A1(_11246_),
    .A2(_11247_),
    .B1(_11257_),
    .Y(_11258_));
 sky130_fd_sc_hd__and2_4 _41797_ (.A(_11256_),
    .B(_11258_),
    .X(_11259_));
 sky130_vsdinv _41798_ (.A(_11259_),
    .Y(_11260_));
 sky130_fd_sc_hd__nand2_4 _41799_ (.A(_11234_),
    .B(_11260_),
    .Y(_11261_));
 sky130_fd_sc_hd__nand3_4 _41800_ (.A(_11231_),
    .B(_11259_),
    .C(_11233_),
    .Y(_11262_));
 sky130_fd_sc_hd__nand2_4 _41801_ (.A(_11261_),
    .B(_11262_),
    .Y(_11263_));
 sky130_fd_sc_hd__a21boi_4 _41802_ (.A1(_10912_),
    .A2(_10917_),
    .B1_N(_10913_),
    .Y(_11264_));
 sky130_fd_sc_hd__nand2_4 _41803_ (.A(_11263_),
    .B(_11264_),
    .Y(_11265_));
 sky130_vsdinv _41804_ (.A(_11264_),
    .Y(_11266_));
 sky130_fd_sc_hd__nand3_4 _41805_ (.A(_11261_),
    .B(_11266_),
    .C(_11262_),
    .Y(_11267_));
 sky130_fd_sc_hd__nand2_4 _41806_ (.A(_11265_),
    .B(_11267_),
    .Y(_11268_));
 sky130_fd_sc_hd__a21boi_4 _41807_ (.A1(_11045_),
    .A2(_11006_),
    .B1_N(_11008_),
    .Y(_11269_));
 sky130_fd_sc_hd__nand2_4 _41808_ (.A(_11268_),
    .B(_11269_),
    .Y(_11270_));
 sky130_vsdinv _41809_ (.A(_11269_),
    .Y(_11271_));
 sky130_fd_sc_hd__nand3_4 _41810_ (.A(_11265_),
    .B(_11271_),
    .C(_11267_),
    .Y(_11272_));
 sky130_fd_sc_hd__nand2_4 _41811_ (.A(_11270_),
    .B(_11272_),
    .Y(_11273_));
 sky130_fd_sc_hd__nand2_4 _41812_ (.A(_11211_),
    .B(_11273_),
    .Y(_11274_));
 sky130_vsdinv _41813_ (.A(_11273_),
    .Y(_11275_));
 sky130_fd_sc_hd__nand3_4 _41814_ (.A(_11275_),
    .B(_11210_),
    .C(_11208_),
    .Y(_11276_));
 sky130_fd_sc_hd__nand2_4 _41815_ (.A(_11274_),
    .B(_11276_),
    .Y(_11277_));
 sky130_fd_sc_hd__o21a_4 _41816_ (.A1(_11059_),
    .A2(_10983_),
    .B1(_10982_),
    .X(_11278_));
 sky130_fd_sc_hd__nand2_4 _41817_ (.A(_11277_),
    .B(_11278_),
    .Y(_11279_));
 sky130_vsdinv _41818_ (.A(_11278_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand3_4 _41819_ (.A(_11280_),
    .B(_11276_),
    .C(_11274_),
    .Y(_11281_));
 sky130_fd_sc_hd__nand2_4 _41820_ (.A(_11279_),
    .B(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__a21boi_4 _41821_ (.A1(_11032_),
    .A2(_11037_),
    .B1_N(_11035_),
    .Y(_11283_));
 sky130_fd_sc_hd__nand2_4 _41822_ (.A(_10666_),
    .B(_08082_),
    .Y(_11284_));
 sky130_fd_sc_hd__nand2_4 _41823_ (.A(_03375_),
    .B(_07096_),
    .Y(_11285_));
 sky130_fd_sc_hd__nand2_4 _41824_ (.A(_11284_),
    .B(_11285_),
    .Y(_11286_));
 sky130_fd_sc_hd__buf_1 _41825_ (.A(_09090_),
    .X(_11287_));
 sky130_fd_sc_hd__nand4_4 _41826_ (.A(_11287_),
    .B(_09846_),
    .C(_06600_),
    .D(_06594_),
    .Y(_11288_));
 sky130_fd_sc_hd__nand2_4 _41827_ (.A(_09847_),
    .B(_06949_),
    .Y(_11289_));
 sky130_vsdinv _41828_ (.A(_11289_),
    .Y(_11290_));
 sky130_fd_sc_hd__a21o_4 _41829_ (.A1(_11286_),
    .A2(_11288_),
    .B1(_11290_),
    .X(_11291_));
 sky130_fd_sc_hd__nand3_4 _41830_ (.A(_11286_),
    .B(_11288_),
    .C(_11290_),
    .Y(_11292_));
 sky130_fd_sc_hd__nand2_4 _41831_ (.A(_11291_),
    .B(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__nor2_4 _41832_ (.A(_11283_),
    .B(_11293_),
    .Y(_11294_));
 sky130_vsdinv _41833_ (.A(_11294_),
    .Y(_11295_));
 sky130_fd_sc_hd__nand2_4 _41834_ (.A(_11293_),
    .B(_11283_),
    .Y(_11296_));
 sky130_fd_sc_hd__a21boi_4 _41835_ (.A1(_10787_),
    .A2(_10793_),
    .B1_N(_10790_),
    .Y(_11297_));
 sky130_vsdinv _41836_ (.A(_11297_),
    .Y(_11298_));
 sky130_fd_sc_hd__a21o_4 _41837_ (.A1(_11295_),
    .A2(_11296_),
    .B1(_11298_),
    .X(_11299_));
 sky130_fd_sc_hd__nand3_4 _41838_ (.A(_11295_),
    .B(_11296_),
    .C(_11298_),
    .Y(_11300_));
 sky130_fd_sc_hd__nand2_4 _41839_ (.A(_11299_),
    .B(_11300_),
    .Y(_11301_));
 sky130_fd_sc_hd__a21boi_4 _41840_ (.A1(_11027_),
    .A2(_11041_),
    .B1_N(_11028_),
    .Y(_11302_));
 sky130_fd_sc_hd__nand2_4 _41841_ (.A(_11301_),
    .B(_11302_),
    .Y(_11303_));
 sky130_vsdinv _41842_ (.A(_11302_),
    .Y(_11304_));
 sky130_fd_sc_hd__nand3_4 _41843_ (.A(_11299_),
    .B(_11304_),
    .C(_11300_),
    .Y(_11305_));
 sky130_fd_sc_hd__nand2_4 _41844_ (.A(_11303_),
    .B(_11305_),
    .Y(_11306_));
 sky130_fd_sc_hd__a21boi_4 _41845_ (.A1(_10798_),
    .A2(_10802_),
    .B1_N(_10800_),
    .Y(_11307_));
 sky130_fd_sc_hd__nand2_4 _41846_ (.A(_11306_),
    .B(_11307_),
    .Y(_11308_));
 sky130_vsdinv _41847_ (.A(_11307_),
    .Y(_11309_));
 sky130_fd_sc_hd__nand3_4 _41848_ (.A(_11303_),
    .B(_11309_),
    .C(_11305_),
    .Y(_11310_));
 sky130_fd_sc_hd__nand2_4 _41849_ (.A(_11308_),
    .B(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__a21boi_4 _41850_ (.A1(_10807_),
    .A2(_10811_),
    .B1_N(_10809_),
    .Y(_11312_));
 sky130_fd_sc_hd__nand2_4 _41851_ (.A(_11311_),
    .B(_11312_),
    .Y(_11313_));
 sky130_vsdinv _41852_ (.A(_11312_),
    .Y(_11314_));
 sky130_fd_sc_hd__nand3_4 _41853_ (.A(_11308_),
    .B(_11314_),
    .C(_11310_),
    .Y(_11315_));
 sky130_fd_sc_hd__nand2_4 _41854_ (.A(_11313_),
    .B(_11315_),
    .Y(_11316_));
 sky130_fd_sc_hd__buf_1 _41855_ (.A(_03382_),
    .X(_11317_));
 sky130_fd_sc_hd__nand2_4 _41856_ (.A(_11317_),
    .B(_03472_),
    .Y(_11318_));
 sky130_fd_sc_hd__buf_1 _41857_ (.A(_03387_),
    .X(_11319_));
 sky130_fd_sc_hd__nand2_4 _41858_ (.A(_11319_),
    .B(_05992_),
    .Y(_11320_));
 sky130_fd_sc_hd__nand2_4 _41859_ (.A(_11318_),
    .B(_11320_),
    .Y(_11321_));
 sky130_fd_sc_hd__nand4_4 _41860_ (.A(_11317_),
    .B(_10087_),
    .C(_06228_),
    .D(_06220_),
    .Y(_11322_));
 sky130_fd_sc_hd__buf_1 _41861_ (.A(_10408_),
    .X(_11323_));
 sky130_fd_sc_hd__nand2_4 _41862_ (.A(_11323_),
    .B(_06232_),
    .Y(_11324_));
 sky130_vsdinv _41863_ (.A(_11324_),
    .Y(_11325_));
 sky130_fd_sc_hd__a21o_4 _41864_ (.A1(_11321_),
    .A2(_11322_),
    .B1(_11325_),
    .X(_11326_));
 sky130_fd_sc_hd__nand3_4 _41865_ (.A(_11321_),
    .B(_11322_),
    .C(_11325_),
    .Y(_11327_));
 sky130_fd_sc_hd__a21boi_4 _41866_ (.A1(_10824_),
    .A2(_10829_),
    .B1_N(_10825_),
    .Y(_11328_));
 sky130_fd_sc_hd__a21boi_4 _41867_ (.A1(_11326_),
    .A2(_11327_),
    .B1_N(_11328_),
    .Y(_11329_));
 sky130_vsdinv _41868_ (.A(_11329_),
    .Y(_11330_));
 sky130_vsdinv _41869_ (.A(_11328_),
    .Y(_11331_));
 sky130_fd_sc_hd__nand3_4 _41870_ (.A(_11331_),
    .B(_11326_),
    .C(_11327_),
    .Y(_11332_));
 sky130_fd_sc_hd__buf_1 _41871_ (.A(\pcpi_mul.rs1[30] ),
    .X(_11333_));
 sky130_fd_sc_hd__buf_1 _41872_ (.A(_11333_),
    .X(_11334_));
 sky130_fd_sc_hd__nand2_4 _41873_ (.A(_11334_),
    .B(_06003_),
    .Y(_11335_));
 sky130_fd_sc_hd__o21ai_4 _41874_ (.A1(_03401_),
    .A2(_07619_),
    .B1(_11335_),
    .Y(_11336_));
 sky130_fd_sc_hd__buf_1 _41875_ (.A(_10836_),
    .X(_11337_));
 sky130_fd_sc_hd__nand4_4 _41876_ (.A(_03397_),
    .B(_11337_),
    .C(_06165_),
    .D(_06706_),
    .Y(_11338_));
 sky130_fd_sc_hd__buf_1 _41877_ (.A(\pcpi_mul.rs1[32] ),
    .X(_11339_));
 sky130_fd_sc_hd__nand2_4 _41878_ (.A(_11339_),
    .B(\pcpi_mul.rs2[0] ),
    .Y(_11340_));
 sky130_vsdinv _41879_ (.A(_11340_),
    .Y(_11341_));
 sky130_fd_sc_hd__buf_4 _41880_ (.A(_11341_),
    .X(_11342_));
 sky130_fd_sc_hd__a21o_4 _41881_ (.A1(_11336_),
    .A2(_11338_),
    .B1(_11342_),
    .X(_11343_));
 sky130_fd_sc_hd__buf_1 _41882_ (.A(_11342_),
    .X(_11344_));
 sky130_fd_sc_hd__nand3_4 _41883_ (.A(_11336_),
    .B(_11338_),
    .C(_11344_),
    .Y(_11345_));
 sky130_fd_sc_hd__and2_4 _41884_ (.A(_11343_),
    .B(_11345_),
    .X(_11346_));
 sky130_fd_sc_hd__buf_1 _41885_ (.A(_11346_),
    .X(_11347_));
 sky130_fd_sc_hd__a21o_4 _41886_ (.A1(_11330_),
    .A2(_11332_),
    .B1(_11347_),
    .X(_11348_));
 sky130_fd_sc_hd__nand3_4 _41887_ (.A(_11330_),
    .B(_11347_),
    .C(_11332_),
    .Y(_11349_));
 sky130_fd_sc_hd__a21oi_4 _41888_ (.A1(_10850_),
    .A2(_10835_),
    .B1(_10833_),
    .Y(_11350_));
 sky130_vsdinv _41889_ (.A(_11350_),
    .Y(_11351_));
 sky130_fd_sc_hd__a21o_4 _41890_ (.A1(_11348_),
    .A2(_11349_),
    .B1(_11351_),
    .X(_11352_));
 sky130_fd_sc_hd__nand3_4 _41891_ (.A(_11351_),
    .B(_11349_),
    .C(_11348_),
    .Y(_11353_));
 sky130_vsdinv _41892_ (.A(_10839_),
    .Y(_11354_));
 sky130_fd_sc_hd__a21boi_4 _41893_ (.A1(_10842_),
    .A2(_11354_),
    .B1_N(_10848_),
    .Y(_11355_));
 sky130_vsdinv _41894_ (.A(_11355_),
    .Y(_11356_));
 sky130_fd_sc_hd__a21o_4 _41895_ (.A1(_11352_),
    .A2(_11353_),
    .B1(_11356_),
    .X(_11357_));
 sky130_fd_sc_hd__nand3_4 _41896_ (.A(_11352_),
    .B(_11356_),
    .C(_11353_),
    .Y(_11358_));
 sky130_fd_sc_hd__and2_4 _41897_ (.A(_11357_),
    .B(_11358_),
    .X(_11359_));
 sky130_vsdinv _41898_ (.A(_11359_),
    .Y(_11360_));
 sky130_fd_sc_hd__nand2_4 _41899_ (.A(_11316_),
    .B(_11360_),
    .Y(_11361_));
 sky130_fd_sc_hd__nand3_4 _41900_ (.A(_11359_),
    .B(_11313_),
    .C(_11315_),
    .Y(_11362_));
 sky130_fd_sc_hd__nand2_4 _41901_ (.A(_11361_),
    .B(_11362_),
    .Y(_11363_));
 sky130_fd_sc_hd__a21boi_4 _41902_ (.A1(_11051_),
    .A2(_11057_),
    .B1_N(_11053_),
    .Y(_11364_));
 sky130_fd_sc_hd__nand2_4 _41903_ (.A(_11363_),
    .B(_11364_),
    .Y(_11365_));
 sky130_vsdinv _41904_ (.A(_11364_),
    .Y(_11366_));
 sky130_fd_sc_hd__nand3_4 _41905_ (.A(_11361_),
    .B(_11366_),
    .C(_11362_),
    .Y(_11367_));
 sky130_fd_sc_hd__a21boi_4 _41906_ (.A1(_10865_),
    .A2(_10816_),
    .B1_N(_10818_),
    .Y(_11368_));
 sky130_vsdinv _41907_ (.A(_11368_),
    .Y(_11369_));
 sky130_fd_sc_hd__a21o_4 _41908_ (.A1(_11365_),
    .A2(_11367_),
    .B1(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__nand3_4 _41909_ (.A(_11365_),
    .B(_11369_),
    .C(_11367_),
    .Y(_11371_));
 sky130_fd_sc_hd__nand2_4 _41910_ (.A(_11370_),
    .B(_11371_),
    .Y(_11372_));
 sky130_fd_sc_hd__nand2_4 _41911_ (.A(_11282_),
    .B(_11372_),
    .Y(_11373_));
 sky130_fd_sc_hd__nand4_4 _41912_ (.A(_11371_),
    .B(_11279_),
    .C(_11370_),
    .D(_11281_),
    .Y(_11374_));
 sky130_fd_sc_hd__nand2_4 _41913_ (.A(_11373_),
    .B(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__nand2_4 _41914_ (.A(_11070_),
    .B(_11067_),
    .Y(_11376_));
 sky130_vsdinv _41915_ (.A(_11376_),
    .Y(_11377_));
 sky130_fd_sc_hd__nand2_4 _41916_ (.A(_11375_),
    .B(_11377_),
    .Y(_11378_));
 sky130_fd_sc_hd__nand3_4 _41917_ (.A(_11373_),
    .B(_11374_),
    .C(_11376_),
    .Y(_11379_));
 sky130_fd_sc_hd__nand2_4 _41918_ (.A(_11378_),
    .B(_11379_),
    .Y(_11380_));
 sky130_fd_sc_hd__a21boi_4 _41919_ (.A1(_10855_),
    .A2(_10858_),
    .B1_N(_10856_),
    .Y(_11381_));
 sky130_fd_sc_hd__a21o_4 _41920_ (.A1(_10876_),
    .A2(_10871_),
    .B1(_11381_),
    .X(_11382_));
 sky130_fd_sc_hd__nand3_4 _41921_ (.A(_10876_),
    .B(_10871_),
    .C(_11381_),
    .Y(_11383_));
 sky130_fd_sc_hd__buf_4 _41922_ (.A(_11106_),
    .X(_11384_));
 sky130_fd_sc_hd__buf_1 _41923_ (.A(_11384_),
    .X(_11385_));
 sky130_fd_sc_hd__buf_1 _41924_ (.A(_11385_),
    .X(_11386_));
 sky130_fd_sc_hd__buf_1 _41925_ (.A(_11386_),
    .X(_11387_));
 sky130_fd_sc_hd__buf_1 _41926_ (.A(_11387_),
    .X(_11388_));
 sky130_fd_sc_hd__a21o_4 _41927_ (.A1(_11382_),
    .A2(_11383_),
    .B1(_11388_),
    .X(_11389_));
 sky130_fd_sc_hd__nand3_4 _41928_ (.A(_11382_),
    .B(_11388_),
    .C(_11383_),
    .Y(_11390_));
 sky130_fd_sc_hd__nand2_4 _41929_ (.A(_11389_),
    .B(_11390_),
    .Y(_11391_));
 sky130_fd_sc_hd__nand2_4 _41930_ (.A(_11380_),
    .B(_11391_),
    .Y(_11392_));
 sky130_vsdinv _41931_ (.A(_11391_),
    .Y(_11393_));
 sky130_fd_sc_hd__nand3_4 _41932_ (.A(_11393_),
    .B(_11378_),
    .C(_11379_),
    .Y(_11394_));
 sky130_fd_sc_hd__nand2_4 _41933_ (.A(_11392_),
    .B(_11394_),
    .Y(_11395_));
 sky130_fd_sc_hd__a21boi_4 _41934_ (.A1(_11074_),
    .A2(_11082_),
    .B1_N(_11076_),
    .Y(_11396_));
 sky130_fd_sc_hd__nand2_4 _41935_ (.A(_11395_),
    .B(_11396_),
    .Y(_11397_));
 sky130_vsdinv _41936_ (.A(_11396_),
    .Y(_11398_));
 sky130_fd_sc_hd__nand3_4 _41937_ (.A(_11392_),
    .B(_11394_),
    .C(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__nand2_4 _41938_ (.A(_11397_),
    .B(_11399_),
    .Y(_11400_));
 sky130_fd_sc_hd__a21oi_4 _41939_ (.A1(_10748_),
    .A2(_10743_),
    .B1(_11078_),
    .Y(_11401_));
 sky130_vsdinv _41940_ (.A(_11401_),
    .Y(_11402_));
 sky130_fd_sc_hd__nand2_4 _41941_ (.A(_11400_),
    .B(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__nand3_4 _41942_ (.A(_11397_),
    .B(_11401_),
    .C(_11399_),
    .Y(_11404_));
 sky130_fd_sc_hd__a21boi_4 _41943_ (.A1(_11086_),
    .A2(_11090_),
    .B1_N(_11088_),
    .Y(_11405_));
 sky130_vsdinv _41944_ (.A(_11405_),
    .Y(_11406_));
 sky130_fd_sc_hd__a21o_4 _41945_ (.A1(_11403_),
    .A2(_11404_),
    .B1(_11406_),
    .X(_11407_));
 sky130_fd_sc_hd__nand3_4 _41946_ (.A(_11403_),
    .B(_11404_),
    .C(_11406_),
    .Y(_11408_));
 sky130_fd_sc_hd__nand2_4 _41947_ (.A(_11407_),
    .B(_11408_),
    .Y(_11409_));
 sky130_fd_sc_hd__nand4_4 _41948_ (.A(_09149_),
    .B(_09645_),
    .C(_09398_),
    .D(_09916_),
    .Y(_11410_));
 sky130_fd_sc_hd__nand4_4 _41949_ (.A(_10187_),
    .B(_10779_),
    .C(_10473_),
    .D(_11099_),
    .Y(_11411_));
 sky130_fd_sc_hd__nor2_4 _41950_ (.A(_11410_),
    .B(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__nand4_4 _41951_ (.A(_10185_),
    .B(_10470_),
    .C(_10183_),
    .D(_10471_),
    .Y(_11413_));
 sky130_fd_sc_hd__nand2_4 _41952_ (.A(_11092_),
    .B(_11093_),
    .Y(_11414_));
 sky130_vsdinv _41953_ (.A(_11095_),
    .Y(_11415_));
 sky130_fd_sc_hd__nand2_4 _41954_ (.A(_11414_),
    .B(_11415_),
    .Y(_11416_));
 sky130_fd_sc_hd__nand4_4 _41955_ (.A(_10777_),
    .B(_10776_),
    .C(_11416_),
    .D(_11097_),
    .Y(_11417_));
 sky130_fd_sc_hd__nor2_4 _41956_ (.A(_11413_),
    .B(_11417_),
    .Y(_11418_));
 sky130_fd_sc_hd__nand2_4 _41957_ (.A(_10191_),
    .B(_11418_),
    .Y(_11419_));
 sky130_fd_sc_hd__nand2_4 _41958_ (.A(_10781_),
    .B(_10470_),
    .Y(_11420_));
 sky130_fd_sc_hd__o21a_4 _41959_ (.A1(_10777_),
    .A2(_11096_),
    .B1(_11097_),
    .X(_11421_));
 sky130_fd_sc_hd__o21a_4 _41960_ (.A1(_11420_),
    .A2(_11417_),
    .B1(_11421_),
    .X(_11422_));
 sky130_fd_sc_hd__nand2_4 _41961_ (.A(_11419_),
    .B(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__a21oi_4 _41962_ (.A1(_09156_),
    .A2(_11412_),
    .B1(_11423_),
    .Y(_11424_));
 vsdcell_nand3_2x _41963_ (.A(_07414_),
    .B(_09152_),
    .C(_11412_),
    .Y(_11425_));
 sky130_fd_sc_hd__nand2_4 _41964_ (.A(_11424_),
    .B(_11425_),
    .Y(_11426_));
 sky130_fd_sc_hd__buf_8 _41965_ (.A(_11426_),
    .X(_11427_));
 sky130_fd_sc_hd__xnor2_4 _41966_ (.A(_11409_),
    .B(_11427_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_4 _41967_ (.A(_11394_),
    .B(_11379_),
    .Y(_11428_));
 sky130_vsdinv _41968_ (.A(_11428_),
    .Y(_11429_));
 sky130_fd_sc_hd__a21boi_4 _41969_ (.A1(_11104_),
    .A2(_11112_),
    .B1_N(_11108_),
    .Y(_11430_));
 sky130_vsdinv _41970_ (.A(_11430_),
    .Y(_11431_));
 sky130_fd_sc_hd__buf_1 _41971_ (.A(_03632_),
    .X(_11432_));
 sky130_fd_sc_hd__buf_1 _41972_ (.A(_03627_),
    .X(_11433_));
 sky130_fd_sc_hd__nand2_4 _41973_ (.A(_05900_),
    .B(_11433_),
    .Y(_11434_));
 sky130_fd_sc_hd__o21ai_4 _41974_ (.A1(_07048_),
    .A2(_11432_),
    .B1(_11434_),
    .Y(_11435_));
 sky130_fd_sc_hd__nand2_4 _41975_ (.A(_07360_),
    .B(_10516_),
    .Y(_11436_));
 sky130_vsdinv _41976_ (.A(_11436_),
    .Y(_11437_));
 sky130_fd_sc_hd__buf_1 _41977_ (.A(_10958_),
    .X(_11438_));
 sky130_fd_sc_hd__nand4_4 _41978_ (.A(_03249_),
    .B(_07359_),
    .C(_11438_),
    .D(_11107_),
    .Y(_11439_));
 sky130_fd_sc_hd__nand3_4 _41979_ (.A(_11435_),
    .B(_11437_),
    .C(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__nand2_4 _41980_ (.A(_11435_),
    .B(_11439_),
    .Y(_11441_));
 sky130_fd_sc_hd__nand2_4 _41981_ (.A(_11441_),
    .B(_11436_),
    .Y(_11442_));
 sky130_fd_sc_hd__nand3_4 _41982_ (.A(_11431_),
    .B(_11440_),
    .C(_11442_),
    .Y(_11443_));
 sky130_fd_sc_hd__nand2_4 _41983_ (.A(_11442_),
    .B(_11440_),
    .Y(_11444_));
 sky130_fd_sc_hd__nand2_4 _41984_ (.A(_11444_),
    .B(_11430_),
    .Y(_11445_));
 sky130_fd_sc_hd__nand2_4 _41985_ (.A(_11443_),
    .B(_11445_),
    .Y(_11446_));
 sky130_fd_sc_hd__buf_1 _41986_ (.A(_10498_),
    .X(_11447_));
 sky130_fd_sc_hd__nand2_4 _41987_ (.A(_10480_),
    .B(_11447_),
    .Y(_11448_));
 sky130_fd_sc_hd__buf_1 _41988_ (.A(_10501_),
    .X(_11449_));
 sky130_fd_sc_hd__nand2_4 _41989_ (.A(_08565_),
    .B(_11449_),
    .Y(_11450_));
 sky130_fd_sc_hd__nand2_4 _41990_ (.A(_11448_),
    .B(_11450_),
    .Y(_11451_));
 sky130_fd_sc_hd__nand4_4 _41991_ (.A(_07740_),
    .B(_07526_),
    .C(_03606_),
    .D(_03613_),
    .Y(_11452_));
 sky130_fd_sc_hd__nand2_4 _41992_ (.A(_07346_),
    .B(_11125_),
    .Y(_11453_));
 sky130_vsdinv _41993_ (.A(_11453_),
    .Y(_11454_));
 sky130_fd_sc_hd__a21o_4 _41994_ (.A1(_11451_),
    .A2(_11452_),
    .B1(_11454_),
    .X(_11455_));
 sky130_fd_sc_hd__nand3_4 _41995_ (.A(_11451_),
    .B(_11452_),
    .C(_11454_),
    .Y(_11456_));
 sky130_fd_sc_hd__nand2_4 _41996_ (.A(_11455_),
    .B(_11456_),
    .Y(_11457_));
 sky130_fd_sc_hd__nand2_4 _41997_ (.A(_11446_),
    .B(_11457_),
    .Y(_11458_));
 sky130_vsdinv _41998_ (.A(_11457_),
    .Y(_11459_));
 sky130_fd_sc_hd__nand3_4 _41999_ (.A(_11443_),
    .B(_11445_),
    .C(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__nand2_4 _42000_ (.A(_11458_),
    .B(_11460_),
    .Y(_11461_));
 sky130_vsdinv _42001_ (.A(_11117_),
    .Y(_11462_));
 sky130_fd_sc_hd__a21oi_4 _42002_ (.A1(_11115_),
    .A2(_11130_),
    .B1(_11462_),
    .Y(_11463_));
 sky130_fd_sc_hd__nand2_4 _42003_ (.A(_11461_),
    .B(_11463_),
    .Y(_11464_));
 sky130_vsdinv _42004_ (.A(_11463_),
    .Y(_11465_));
 sky130_fd_sc_hd__nand3_4 _42005_ (.A(_11465_),
    .B(_11460_),
    .C(_11458_),
    .Y(_11466_));
 sky130_fd_sc_hd__nand2_4 _42006_ (.A(_11464_),
    .B(_11466_),
    .Y(_11467_));
 sky130_fd_sc_hd__a21boi_4 _42007_ (.A1(_11123_),
    .A2(_11127_),
    .B1_N(_11124_),
    .Y(_11468_));
 sky130_fd_sc_hd__nand2_4 _42008_ (.A(_06155_),
    .B(_10920_),
    .Y(_11469_));
 sky130_fd_sc_hd__nand2_4 _42009_ (.A(_07758_),
    .B(_03587_),
    .Y(_11470_));
 sky130_fd_sc_hd__nand2_4 _42010_ (.A(_11469_),
    .B(_11470_),
    .Y(_11471_));
 sky130_fd_sc_hd__nand4_4 _42011_ (.A(_06340_),
    .B(_07959_),
    .C(_09344_),
    .D(_10925_),
    .Y(_11472_));
 sky130_fd_sc_hd__buf_1 _42012_ (.A(_03580_),
    .X(_11473_));
 sky130_fd_sc_hd__nand2_4 _42013_ (.A(_10265_),
    .B(_11473_),
    .Y(_11474_));
 sky130_vsdinv _42014_ (.A(_11474_),
    .Y(_11475_));
 sky130_fd_sc_hd__a21o_4 _42015_ (.A1(_11471_),
    .A2(_11472_),
    .B1(_11475_),
    .X(_11476_));
 sky130_fd_sc_hd__nand3_4 _42016_ (.A(_11471_),
    .B(_11472_),
    .C(_11475_),
    .Y(_11477_));
 sky130_fd_sc_hd__nand2_4 _42017_ (.A(_11476_),
    .B(_11477_),
    .Y(_11478_));
 sky130_fd_sc_hd__nor2_4 _42018_ (.A(_11468_),
    .B(_11478_),
    .Y(_11479_));
 sky130_vsdinv _42019_ (.A(_11479_),
    .Y(_11480_));
 sky130_fd_sc_hd__a21boi_4 _42020_ (.A1(_11141_),
    .A2(_11145_),
    .B1_N(_11143_),
    .Y(_11481_));
 sky130_vsdinv _42021_ (.A(_11481_),
    .Y(_11482_));
 sky130_fd_sc_hd__nand2_4 _42022_ (.A(_11478_),
    .B(_11468_),
    .Y(_11483_));
 sky130_fd_sc_hd__nand3_4 _42023_ (.A(_11480_),
    .B(_11482_),
    .C(_11483_),
    .Y(_11484_));
 sky130_fd_sc_hd__a21boi_4 _42024_ (.A1(_11476_),
    .A2(_11477_),
    .B1_N(_11468_),
    .Y(_11485_));
 sky130_fd_sc_hd__o21ai_4 _42025_ (.A1(_11485_),
    .A2(_11479_),
    .B1(_11481_),
    .Y(_11486_));
 sky130_fd_sc_hd__nand2_4 _42026_ (.A(_11484_),
    .B(_11486_),
    .Y(_11487_));
 sky130_fd_sc_hd__nand2_4 _42027_ (.A(_11467_),
    .B(_11487_),
    .Y(_11488_));
 sky130_vsdinv _42028_ (.A(_11487_),
    .Y(_11489_));
 sky130_fd_sc_hd__nand3_4 _42029_ (.A(_11464_),
    .B(_11489_),
    .C(_11466_),
    .Y(_11490_));
 sky130_fd_sc_hd__nand2_4 _42030_ (.A(_11488_),
    .B(_11490_),
    .Y(_11491_));
 sky130_vsdinv _42031_ (.A(_11137_),
    .Y(_11492_));
 sky130_fd_sc_hd__a21o_4 _42032_ (.A1(_11135_),
    .A2(_11159_),
    .B1(_11492_),
    .X(_11493_));
 sky130_vsdinv _42033_ (.A(_11493_),
    .Y(_11494_));
 sky130_fd_sc_hd__nand2_4 _42034_ (.A(_11491_),
    .B(_11494_),
    .Y(_11495_));
 sky130_fd_sc_hd__nand3_4 _42035_ (.A(_11493_),
    .B(_11488_),
    .C(_11490_),
    .Y(_11496_));
 sky130_fd_sc_hd__nand2_4 _42036_ (.A(_11495_),
    .B(_11496_),
    .Y(_11497_));
 sky130_fd_sc_hd__maj3_4 _42037_ (.A(_11168_),
    .B(_11176_),
    .C(_11170_),
    .X(_11498_));
 sky130_vsdinv _42038_ (.A(_11498_),
    .Y(_11499_));
 sky130_fd_sc_hd__nand2_4 _42039_ (.A(_07130_),
    .B(_11169_),
    .Y(_11500_));
 sky130_fd_sc_hd__o21ai_4 _42040_ (.A1(_03295_),
    .A2(_03577_),
    .B1(_11500_),
    .Y(_11501_));
 sky130_fd_sc_hd__buf_1 _42041_ (.A(_03569_),
    .X(_11502_));
 sky130_fd_sc_hd__buf_1 _42042_ (.A(_10275_),
    .X(_11503_));
 sky130_fd_sc_hd__nand4_4 _42043_ (.A(_06981_),
    .B(_07130_),
    .C(_11502_),
    .D(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__nand2_4 _42044_ (.A(_07416_),
    .B(_10540_),
    .Y(_11505_));
 sky130_vsdinv _42045_ (.A(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__nand3_4 _42046_ (.A(_11501_),
    .B(_11504_),
    .C(_11506_),
    .Y(_11507_));
 sky130_fd_sc_hd__nand2_4 _42047_ (.A(_11501_),
    .B(_11504_),
    .Y(_11508_));
 sky130_fd_sc_hd__nand2_4 _42048_ (.A(_11508_),
    .B(_11505_),
    .Y(_11509_));
 sky130_fd_sc_hd__nand3_4 _42049_ (.A(_11499_),
    .B(_11507_),
    .C(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__nand2_4 _42050_ (.A(_11509_),
    .B(_11507_),
    .Y(_11511_));
 sky130_fd_sc_hd__nand2_4 _42051_ (.A(_11511_),
    .B(_11498_),
    .Y(_11512_));
 sky130_fd_sc_hd__buf_1 _42052_ (.A(_08026_),
    .X(_11513_));
 sky130_fd_sc_hd__buf_1 _42053_ (.A(_07979_),
    .X(_11514_));
 sky130_fd_sc_hd__nand2_4 _42054_ (.A(_11513_),
    .B(_11514_),
    .Y(_11515_));
 sky130_fd_sc_hd__buf_1 _42055_ (.A(_08194_),
    .X(_11516_));
 sky130_fd_sc_hd__nand2_4 _42056_ (.A(_07006_),
    .B(_11516_),
    .Y(_11517_));
 sky130_fd_sc_hd__buf_1 _42057_ (.A(_10262_),
    .X(_11518_));
 sky130_fd_sc_hd__nand2_4 _42058_ (.A(_06993_),
    .B(_11518_),
    .Y(_11519_));
 sky130_fd_sc_hd__nand2_4 _42059_ (.A(_11517_),
    .B(_11519_),
    .Y(_11520_));
 sky130_fd_sc_hd__buf_1 _42060_ (.A(_08191_),
    .X(_11521_));
 sky130_fd_sc_hd__buf_1 _42061_ (.A(_08647_),
    .X(_11522_));
 sky130_fd_sc_hd__buf_1 _42062_ (.A(_11522_),
    .X(_11523_));
 sky130_fd_sc_hd__nand4_4 _42063_ (.A(_07006_),
    .B(_06993_),
    .C(_11521_),
    .D(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__nand2_4 _42064_ (.A(_11520_),
    .B(_11524_),
    .Y(_11525_));
 sky130_fd_sc_hd__xor2_4 _42065_ (.A(_11515_),
    .B(_11525_),
    .X(_11526_));
 sky130_fd_sc_hd__a21o_4 _42066_ (.A1(_11510_),
    .A2(_11512_),
    .B1(_11526_),
    .X(_11527_));
 sky130_fd_sc_hd__nand3_4 _42067_ (.A(_11510_),
    .B(_11512_),
    .C(_11526_),
    .Y(_11528_));
 sky130_fd_sc_hd__a21boi_4 _42068_ (.A1(_11150_),
    .A2(_11154_),
    .B1_N(_11152_),
    .Y(_11529_));
 sky130_vsdinv _42069_ (.A(_11529_),
    .Y(_11530_));
 sky130_fd_sc_hd__a21oi_4 _42070_ (.A1(_11527_),
    .A2(_11528_),
    .B1(_11530_),
    .Y(_11531_));
 sky130_fd_sc_hd__nand3_4 _42071_ (.A(_11527_),
    .B(_11530_),
    .C(_11528_),
    .Y(_11532_));
 sky130_vsdinv _42072_ (.A(_11532_),
    .Y(_11533_));
 sky130_vsdinv _42073_ (.A(_11182_),
    .Y(_11534_));
 sky130_fd_sc_hd__a21oi_4 _42074_ (.A1(_11190_),
    .A2(_11181_),
    .B1(_11534_),
    .Y(_11535_));
 sky130_fd_sc_hd__o21ai_4 _42075_ (.A1(_11531_),
    .A2(_11533_),
    .B1(_11535_),
    .Y(_11536_));
 sky130_vsdinv _42076_ (.A(_11531_),
    .Y(_11537_));
 sky130_vsdinv _42077_ (.A(_11535_),
    .Y(_11538_));
 sky130_fd_sc_hd__nand3_4 _42078_ (.A(_11537_),
    .B(_11538_),
    .C(_11532_),
    .Y(_11539_));
 sky130_fd_sc_hd__nand2_4 _42079_ (.A(_11536_),
    .B(_11539_),
    .Y(_11540_));
 sky130_fd_sc_hd__nand2_4 _42080_ (.A(_11497_),
    .B(_11540_),
    .Y(_11541_));
 sky130_vsdinv _42081_ (.A(_11540_),
    .Y(_11542_));
 sky130_fd_sc_hd__nand3_4 _42082_ (.A(_11542_),
    .B(_11496_),
    .C(_11495_),
    .Y(_11543_));
 sky130_fd_sc_hd__nand2_4 _42083_ (.A(_11541_),
    .B(_11543_),
    .Y(_11544_));
 sky130_vsdinv _42084_ (.A(_11163_),
    .Y(_11545_));
 sky130_fd_sc_hd__o21a_4 _42085_ (.A1(_11203_),
    .A2(_11545_),
    .B1(_11165_),
    .X(_11546_));
 sky130_fd_sc_hd__nand2_4 _42086_ (.A(_11544_),
    .B(_11546_),
    .Y(_11547_));
 sky130_fd_sc_hd__o21ai_4 _42087_ (.A1(_11203_),
    .A2(_11545_),
    .B1(_11165_),
    .Y(_11548_));
 sky130_fd_sc_hd__nand3_4 _42088_ (.A(_11548_),
    .B(_11543_),
    .C(_11541_),
    .Y(_11549_));
 sky130_fd_sc_hd__nand2_4 _42089_ (.A(_11547_),
    .B(_11549_),
    .Y(_11550_));
 sky130_vsdinv _42090_ (.A(_11183_),
    .Y(_11551_));
 sky130_fd_sc_hd__a21boi_4 _42091_ (.A1(_11185_),
    .A2(_11551_),
    .B1_N(_11188_),
    .Y(_11552_));
 sky130_fd_sc_hd__nand2_4 _42092_ (.A(_10605_),
    .B(_03541_),
    .Y(_11553_));
 sky130_fd_sc_hd__nand2_4 _42093_ (.A(_07444_),
    .B(_08128_),
    .Y(_11554_));
 sky130_fd_sc_hd__nand2_4 _42094_ (.A(_11553_),
    .B(_11554_),
    .Y(_11555_));
 sky130_fd_sc_hd__buf_1 _42095_ (.A(_09037_),
    .X(_11556_));
 sky130_fd_sc_hd__buf_1 _42096_ (.A(_07874_),
    .X(_11557_));
 sky130_fd_sc_hd__nand4_4 _42097_ (.A(_11556_),
    .B(_11557_),
    .C(_07917_),
    .D(_07915_),
    .Y(_11558_));
 sky130_fd_sc_hd__buf_1 _42098_ (.A(_03336_),
    .X(_11559_));
 sky130_fd_sc_hd__nand2_4 _42099_ (.A(_11559_),
    .B(_08132_),
    .Y(_11560_));
 sky130_vsdinv _42100_ (.A(_11560_),
    .Y(_11561_));
 sky130_fd_sc_hd__a21o_4 _42101_ (.A1(_11555_),
    .A2(_11558_),
    .B1(_11561_),
    .X(_11562_));
 sky130_fd_sc_hd__nand3_4 _42102_ (.A(_11555_),
    .B(_11558_),
    .C(_11561_),
    .Y(_11563_));
 sky130_fd_sc_hd__nand2_4 _42103_ (.A(_11562_),
    .B(_11563_),
    .Y(_11564_));
 sky130_fd_sc_hd__nor2_4 _42104_ (.A(_11552_),
    .B(_11564_),
    .Y(_11565_));
 sky130_vsdinv _42105_ (.A(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__nand2_4 _42106_ (.A(_11564_),
    .B(_11552_),
    .Y(_11567_));
 sky130_fd_sc_hd__a21boi_4 _42107_ (.A1(_11214_),
    .A2(_11217_),
    .B1_N(_11215_),
    .Y(_11568_));
 sky130_vsdinv _42108_ (.A(_11568_),
    .Y(_11569_));
 sky130_fd_sc_hd__a21o_4 _42109_ (.A1(_11566_),
    .A2(_11567_),
    .B1(_11569_),
    .X(_11570_));
 sky130_fd_sc_hd__nand3_4 _42110_ (.A(_11566_),
    .B(_11567_),
    .C(_11569_),
    .Y(_11571_));
 sky130_fd_sc_hd__nand2_4 _42111_ (.A(_11570_),
    .B(_11571_),
    .Y(_11572_));
 sky130_fd_sc_hd__maj3_4 _42112_ (.A(_11225_),
    .B(_11220_),
    .C(_11222_),
    .X(_11573_));
 sky130_fd_sc_hd__nand2_4 _42113_ (.A(_11572_),
    .B(_11573_),
    .Y(_11574_));
 sky130_vsdinv _42114_ (.A(_11573_),
    .Y(_11575_));
 sky130_fd_sc_hd__nand3_4 _42115_ (.A(_11570_),
    .B(_11575_),
    .C(_11571_),
    .Y(_11576_));
 sky130_fd_sc_hd__nand2_4 _42116_ (.A(_11574_),
    .B(_11576_),
    .Y(_11577_));
 sky130_fd_sc_hd__maj3_4 _42117_ (.A(_11240_),
    .B(_11236_),
    .C(_11237_),
    .X(_11578_));
 sky130_fd_sc_hd__nand2_4 _42118_ (.A(_11019_),
    .B(_07055_),
    .Y(_11579_));
 sky130_fd_sc_hd__nand2_4 _42119_ (.A(_11242_),
    .B(_07059_),
    .Y(_11580_));
 sky130_fd_sc_hd__nand2_4 _42120_ (.A(_11579_),
    .B(_11580_),
    .Y(_11581_));
 sky130_fd_sc_hd__nand4_4 _42121_ (.A(_10624_),
    .B(_11033_),
    .C(_07522_),
    .D(_07523_),
    .Y(_11582_));
 sky130_fd_sc_hd__nand2_4 _42122_ (.A(_11034_),
    .B(_07744_),
    .Y(_11583_));
 sky130_vsdinv _42123_ (.A(_11583_),
    .Y(_11584_));
 sky130_fd_sc_hd__a21o_4 _42124_ (.A1(_11581_),
    .A2(_11582_),
    .B1(_11584_),
    .X(_11585_));
 sky130_fd_sc_hd__nand3_4 _42125_ (.A(_11581_),
    .B(_11582_),
    .C(_11584_),
    .Y(_11586_));
 sky130_fd_sc_hd__nand2_4 _42126_ (.A(_11585_),
    .B(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__nor2_4 _42127_ (.A(_11578_),
    .B(_11587_),
    .Y(_11588_));
 sky130_fd_sc_hd__a21boi_4 _42128_ (.A1(_11586_),
    .A2(_11585_),
    .B1_N(_11578_),
    .Y(_11589_));
 sky130_fd_sc_hd__buf_1 _42129_ (.A(_07754_),
    .X(_11590_));
 sky130_fd_sc_hd__nand2_4 _42130_ (.A(_09577_),
    .B(_11590_),
    .Y(_11591_));
 sky130_vsdinv _42131_ (.A(_11591_),
    .Y(_11592_));
 sky130_fd_sc_hd__buf_1 _42132_ (.A(_09202_),
    .X(_11593_));
 sky130_fd_sc_hd__nand2_4 _42133_ (.A(_11593_),
    .B(_07544_),
    .Y(_11594_));
 sky130_fd_sc_hd__buf_1 _42134_ (.A(_09088_),
    .X(_11595_));
 sky130_fd_sc_hd__nand2_4 _42135_ (.A(_11595_),
    .B(_07542_),
    .Y(_11596_));
 sky130_fd_sc_hd__xnor2_4 _42136_ (.A(_11594_),
    .B(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__xor2_4 _42137_ (.A(_11592_),
    .B(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__o21a_4 _42138_ (.A1(_11588_),
    .A2(_11589_),
    .B1(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__xor2_4 _42139_ (.A(_11591_),
    .B(_11597_),
    .X(_11600_));
 sky130_vsdinv _42140_ (.A(_11589_),
    .Y(_11601_));
 sky130_vsdinv _42141_ (.A(_11588_),
    .Y(_11602_));
 sky130_fd_sc_hd__nand3_4 _42142_ (.A(_11600_),
    .B(_11601_),
    .C(_11602_),
    .Y(_11603_));
 sky130_vsdinv _42143_ (.A(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__nor2_4 _42144_ (.A(_11599_),
    .B(_11604_),
    .Y(_11605_));
 sky130_vsdinv _42145_ (.A(_11605_),
    .Y(_11606_));
 sky130_fd_sc_hd__nand2_4 _42146_ (.A(_11577_),
    .B(_11606_),
    .Y(_11607_));
 sky130_fd_sc_hd__nand3_4 _42147_ (.A(_11574_),
    .B(_11605_),
    .C(_11576_),
    .Y(_11608_));
 sky130_fd_sc_hd__nand2_4 _42148_ (.A(_11607_),
    .B(_11608_),
    .Y(_11609_));
 sky130_fd_sc_hd__a21boi_4 _42149_ (.A1(_11195_),
    .A2(_11200_),
    .B1_N(_11198_),
    .Y(_11610_));
 sky130_fd_sc_hd__nand2_4 _42150_ (.A(_11609_),
    .B(_11610_),
    .Y(_11611_));
 sky130_vsdinv _42151_ (.A(_11610_),
    .Y(_11612_));
 sky130_fd_sc_hd__nand3_4 _42152_ (.A(_11612_),
    .B(_11607_),
    .C(_11608_),
    .Y(_11613_));
 sky130_fd_sc_hd__nand2_4 _42153_ (.A(_11611_),
    .B(_11613_),
    .Y(_11614_));
 sky130_fd_sc_hd__a21boi_4 _42154_ (.A1(_11231_),
    .A2(_11259_),
    .B1_N(_11233_),
    .Y(_11615_));
 sky130_fd_sc_hd__nand2_4 _42155_ (.A(_11614_),
    .B(_11615_),
    .Y(_11616_));
 sky130_vsdinv _42156_ (.A(_11615_),
    .Y(_11617_));
 sky130_fd_sc_hd__nand3_4 _42157_ (.A(_11611_),
    .B(_11617_),
    .C(_11613_),
    .Y(_11618_));
 sky130_fd_sc_hd__nand2_4 _42158_ (.A(_11616_),
    .B(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__nand2_4 _42159_ (.A(_11550_),
    .B(_11619_),
    .Y(_11620_));
 sky130_fd_sc_hd__a21oi_4 _42160_ (.A1(_11611_),
    .A2(_11613_),
    .B1(_11617_),
    .Y(_11621_));
 sky130_vsdinv _42161_ (.A(_11618_),
    .Y(_11622_));
 sky130_fd_sc_hd__nor2_4 _42162_ (.A(_11621_),
    .B(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__nand3_4 _42163_ (.A(_11623_),
    .B(_11549_),
    .C(_11547_),
    .Y(_11624_));
 sky130_fd_sc_hd__nand2_4 _42164_ (.A(_11620_),
    .B(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__a21boi_4 _42165_ (.A1(_11275_),
    .A2(_11208_),
    .B1_N(_11210_),
    .Y(_11626_));
 sky130_fd_sc_hd__nand2_4 _42166_ (.A(_11625_),
    .B(_11626_),
    .Y(_11627_));
 sky130_vsdinv _42167_ (.A(_11208_),
    .Y(_11628_));
 sky130_fd_sc_hd__o21ai_4 _42168_ (.A1(_11273_),
    .A2(_11628_),
    .B1(_11210_),
    .Y(_11629_));
 sky130_fd_sc_hd__nand3_4 _42169_ (.A(_11629_),
    .B(_11624_),
    .C(_11620_),
    .Y(_11630_));
 sky130_fd_sc_hd__nand2_4 _42170_ (.A(_11627_),
    .B(_11630_),
    .Y(_11631_));
 sky130_vsdinv _42171_ (.A(_11250_),
    .Y(_11632_));
 sky130_fd_sc_hd__a21boi_4 _42172_ (.A1(_11252_),
    .A2(_11632_),
    .B1_N(_11253_),
    .Y(_11633_));
 sky130_vsdinv _42173_ (.A(_11633_),
    .Y(_11634_));
 sky130_fd_sc_hd__buf_1 _42174_ (.A(_09214_),
    .X(_11635_));
 sky130_fd_sc_hd__nand2_4 _42175_ (.A(_11635_),
    .B(_07470_),
    .Y(_11636_));
 sky130_fd_sc_hd__nand2_4 _42176_ (.A(_10080_),
    .B(_06791_),
    .Y(_11637_));
 sky130_fd_sc_hd__nand2_4 _42177_ (.A(_11636_),
    .B(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__buf_1 _42178_ (.A(_10393_),
    .X(_11639_));
 sky130_fd_sc_hd__nand4_4 _42179_ (.A(_10791_),
    .B(_11639_),
    .C(_06478_),
    .D(_06373_),
    .Y(_11640_));
 sky130_fd_sc_hd__nand2_4 _42180_ (.A(_11638_),
    .B(_11640_),
    .Y(_11641_));
 sky130_fd_sc_hd__nand2_4 _42181_ (.A(_10822_),
    .B(_06797_),
    .Y(_11642_));
 sky130_fd_sc_hd__nand2_4 _42182_ (.A(_11641_),
    .B(_11642_),
    .Y(_11643_));
 sky130_vsdinv _42183_ (.A(_11642_),
    .Y(_11644_));
 sky130_fd_sc_hd__nand3_4 _42184_ (.A(_11638_),
    .B(_11640_),
    .C(_11644_),
    .Y(_11645_));
 sky130_fd_sc_hd__nand3_4 _42185_ (.A(_11634_),
    .B(_11643_),
    .C(_11645_),
    .Y(_11646_));
 sky130_fd_sc_hd__nand2_4 _42186_ (.A(_11643_),
    .B(_11645_),
    .Y(_11647_));
 sky130_fd_sc_hd__nand2_4 _42187_ (.A(_11647_),
    .B(_11633_),
    .Y(_11648_));
 sky130_fd_sc_hd__a21boi_4 _42188_ (.A1(_11286_),
    .A2(_11290_),
    .B1_N(_11288_),
    .Y(_11649_));
 sky130_vsdinv _42189_ (.A(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__a21o_4 _42190_ (.A1(_11646_),
    .A2(_11648_),
    .B1(_11650_),
    .X(_11651_));
 sky130_fd_sc_hd__nand3_4 _42191_ (.A(_11646_),
    .B(_11648_),
    .C(_11650_),
    .Y(_11652_));
 sky130_fd_sc_hd__nand2_4 _42192_ (.A(_11651_),
    .B(_11652_),
    .Y(_11653_));
 sky130_vsdinv _42193_ (.A(_11246_),
    .Y(_11654_));
 sky130_fd_sc_hd__nand3_4 _42194_ (.A(_11653_),
    .B(_11654_),
    .C(_11256_),
    .Y(_11655_));
 sky130_fd_sc_hd__o21ai_4 _42195_ (.A1(_11247_),
    .A2(_11257_),
    .B1(_11654_),
    .Y(_11656_));
 sky130_fd_sc_hd__nand3_4 _42196_ (.A(_11656_),
    .B(_11652_),
    .C(_11651_),
    .Y(_11657_));
 sky130_fd_sc_hd__nand2_4 _42197_ (.A(_11655_),
    .B(_11657_),
    .Y(_11658_));
 sky130_fd_sc_hd__a21oi_4 _42198_ (.A1(_11296_),
    .A2(_11298_),
    .B1(_11294_),
    .Y(_11659_));
 sky130_fd_sc_hd__nand2_4 _42199_ (.A(_11658_),
    .B(_11659_),
    .Y(_11660_));
 sky130_vsdinv _42200_ (.A(_11659_),
    .Y(_11661_));
 sky130_fd_sc_hd__nand3_4 _42201_ (.A(_11655_),
    .B(_11661_),
    .C(_11657_),
    .Y(_11662_));
 sky130_fd_sc_hd__nand2_4 _42202_ (.A(_11660_),
    .B(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__a21boi_4 _42203_ (.A1(_11303_),
    .A2(_11309_),
    .B1_N(_11305_),
    .Y(_11664_));
 sky130_fd_sc_hd__nand2_4 _42204_ (.A(_11663_),
    .B(_11664_),
    .Y(_11665_));
 sky130_fd_sc_hd__nand2_4 _42205_ (.A(_11310_),
    .B(_11305_),
    .Y(_11666_));
 sky130_fd_sc_hd__nand3_4 _42206_ (.A(_11666_),
    .B(_11662_),
    .C(_11660_),
    .Y(_11667_));
 sky130_fd_sc_hd__nand2_4 _42207_ (.A(_11665_),
    .B(_11667_),
    .Y(_11668_));
 sky130_fd_sc_hd__a21boi_4 _42208_ (.A1(_11321_),
    .A2(_11325_),
    .B1_N(_11322_),
    .Y(_11669_));
 sky130_fd_sc_hd__nand2_4 _42209_ (.A(_11319_),
    .B(_06128_),
    .Y(_11670_));
 sky130_fd_sc_hd__nand2_4 _42210_ (.A(_10715_),
    .B(_06130_),
    .Y(_11671_));
 sky130_fd_sc_hd__nand2_4 _42211_ (.A(_11670_),
    .B(_11671_),
    .Y(_11672_));
 sky130_fd_sc_hd__buf_1 _42212_ (.A(_03393_),
    .X(_11673_));
 sky130_fd_sc_hd__nand4_4 _42213_ (.A(_10827_),
    .B(_11673_),
    .C(_07132_),
    .D(_07128_),
    .Y(_11674_));
 sky130_fd_sc_hd__buf_1 _42214_ (.A(_11333_),
    .X(_11675_));
 sky130_fd_sc_hd__nand2_4 _42215_ (.A(_11675_),
    .B(_06232_),
    .Y(_11676_));
 sky130_vsdinv _42216_ (.A(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__a21o_4 _42217_ (.A1(_11672_),
    .A2(_11674_),
    .B1(_11677_),
    .X(_11678_));
 sky130_fd_sc_hd__nand3_4 _42218_ (.A(_11672_),
    .B(_11674_),
    .C(_11677_),
    .Y(_11679_));
 sky130_fd_sc_hd__nand2_4 _42219_ (.A(_11678_),
    .B(_11679_),
    .Y(_11680_));
 sky130_fd_sc_hd__nor2_4 _42220_ (.A(_11669_),
    .B(_11680_),
    .Y(_11681_));
 sky130_vsdinv _42221_ (.A(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__buf_1 _42222_ (.A(\pcpi_mul.rs1[31] ),
    .X(_11683_));
 sky130_fd_sc_hd__buf_1 _42223_ (.A(_11683_),
    .X(_11684_));
 sky130_fd_sc_hd__nand2_4 _42224_ (.A(_11684_),
    .B(_06073_),
    .Y(_11685_));
 sky130_fd_sc_hd__buf_1 _42225_ (.A(_03405_),
    .X(_11686_));
 sky130_fd_sc_hd__buf_1 _42226_ (.A(_11686_),
    .X(_11687_));
 sky130_fd_sc_hd__nand2_4 _42227_ (.A(_11687_),
    .B(_05947_),
    .Y(_11688_));
 sky130_fd_sc_hd__nand2_4 _42228_ (.A(_11685_),
    .B(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__buf_1 _42229_ (.A(_10836_),
    .X(_11690_));
 sky130_fd_sc_hd__buf_4 _42230_ (.A(_03405_),
    .X(_11691_));
 sky130_fd_sc_hd__buf_4 _42231_ (.A(_11691_),
    .X(_11692_));
 sky130_fd_sc_hd__nand4_4 _42232_ (.A(_11690_),
    .B(_11692_),
    .C(_08310_),
    .D(_08311_),
    .Y(_11693_));
 sky130_fd_sc_hd__a21o_4 _42233_ (.A1(_11689_),
    .A2(_11693_),
    .B1(_11342_),
    .X(_11694_));
 sky130_fd_sc_hd__nand3_4 _42234_ (.A(_11689_),
    .B(_11693_),
    .C(_11342_),
    .Y(_11695_));
 sky130_fd_sc_hd__and2_4 _42235_ (.A(_11694_),
    .B(_11695_),
    .X(_11696_));
 sky130_fd_sc_hd__a21boi_4 _42236_ (.A1(_11678_),
    .A2(_11679_),
    .B1_N(_11669_),
    .Y(_11697_));
 sky130_vsdinv _42237_ (.A(_11697_),
    .Y(_11698_));
 sky130_fd_sc_hd__nand3_4 _42238_ (.A(_11682_),
    .B(_11696_),
    .C(_11698_),
    .Y(_11699_));
 sky130_vsdinv _42239_ (.A(_11696_),
    .Y(_11700_));
 sky130_fd_sc_hd__o21ai_4 _42240_ (.A1(_11697_),
    .A2(_11681_),
    .B1(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__nand2_4 _42241_ (.A(_11699_),
    .B(_11701_),
    .Y(_11702_));
 sky130_fd_sc_hd__a21o_4 _42242_ (.A1(_11332_),
    .A2(_11349_),
    .B1(_11702_),
    .X(_11703_));
 sky130_fd_sc_hd__a21boi_4 _42243_ (.A1(_11330_),
    .A2(_11347_),
    .B1_N(_11332_),
    .Y(_11704_));
 sky130_fd_sc_hd__nand2_4 _42244_ (.A(_11702_),
    .B(_11704_),
    .Y(_11705_));
 sky130_fd_sc_hd__a21boi_4 _42245_ (.A1(_11336_),
    .A2(_11344_),
    .B1_N(_11338_),
    .Y(_11706_));
 sky130_vsdinv _42246_ (.A(_11706_),
    .Y(_11707_));
 sky130_fd_sc_hd__a21oi_4 _42247_ (.A1(_11703_),
    .A2(_11705_),
    .B1(_11707_),
    .Y(_11708_));
 sky130_fd_sc_hd__nand3_4 _42248_ (.A(_11703_),
    .B(_11707_),
    .C(_11705_),
    .Y(_11709_));
 sky130_vsdinv _42249_ (.A(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__nor2_4 _42250_ (.A(_11708_),
    .B(_11710_),
    .Y(_11711_));
 sky130_vsdinv _42251_ (.A(_11711_),
    .Y(_11712_));
 sky130_fd_sc_hd__nand2_4 _42252_ (.A(_11668_),
    .B(_11712_),
    .Y(_11713_));
 sky130_fd_sc_hd__nand3_4 _42253_ (.A(_11665_),
    .B(_11667_),
    .C(_11711_),
    .Y(_11714_));
 sky130_fd_sc_hd__nand2_4 _42254_ (.A(_11713_),
    .B(_11714_),
    .Y(_11715_));
 sky130_fd_sc_hd__a21boi_4 _42255_ (.A1(_11265_),
    .A2(_11271_),
    .B1_N(_11267_),
    .Y(_11716_));
 sky130_fd_sc_hd__nand2_4 _42256_ (.A(_11715_),
    .B(_11716_),
    .Y(_11717_));
 sky130_vsdinv _42257_ (.A(_11716_),
    .Y(_11718_));
 sky130_fd_sc_hd__nand3_4 _42258_ (.A(_11718_),
    .B(_11714_),
    .C(_11713_),
    .Y(_11719_));
 sky130_fd_sc_hd__nand2_4 _42259_ (.A(_11717_),
    .B(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__a21boi_4 _42260_ (.A1(_11359_),
    .A2(_11313_),
    .B1_N(_11315_),
    .Y(_11721_));
 sky130_fd_sc_hd__nand2_4 _42261_ (.A(_11720_),
    .B(_11721_),
    .Y(_11722_));
 sky130_vsdinv _42262_ (.A(_11721_),
    .Y(_11723_));
 sky130_fd_sc_hd__nand3_4 _42263_ (.A(_11717_),
    .B(_11719_),
    .C(_11723_),
    .Y(_11724_));
 sky130_fd_sc_hd__nand2_4 _42264_ (.A(_11722_),
    .B(_11724_),
    .Y(_11725_));
 sky130_fd_sc_hd__nand2_4 _42265_ (.A(_11631_),
    .B(_11725_),
    .Y(_11726_));
 sky130_vsdinv _42266_ (.A(_11725_),
    .Y(_11727_));
 sky130_fd_sc_hd__nand3_4 _42267_ (.A(_11727_),
    .B(_11630_),
    .C(_11627_),
    .Y(_11728_));
 sky130_fd_sc_hd__nand2_4 _42268_ (.A(_11726_),
    .B(_11728_),
    .Y(_11729_));
 sky130_vsdinv _42269_ (.A(_11279_),
    .Y(_11730_));
 sky130_fd_sc_hd__o21a_4 _42270_ (.A1(_11372_),
    .A2(_11730_),
    .B1(_11281_),
    .X(_11731_));
 sky130_fd_sc_hd__nand2_4 _42271_ (.A(_11729_),
    .B(_11731_),
    .Y(_11732_));
 sky130_fd_sc_hd__o21ai_4 _42272_ (.A1(_11372_),
    .A2(_11730_),
    .B1(_11281_),
    .Y(_11733_));
 sky130_fd_sc_hd__nand3_4 _42273_ (.A(_11733_),
    .B(_11726_),
    .C(_11728_),
    .Y(_11734_));
 sky130_fd_sc_hd__nand2_4 _42274_ (.A(_11732_),
    .B(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__a21boi_4 _42275_ (.A1(_11352_),
    .A2(_11356_),
    .B1_N(_11353_),
    .Y(_11736_));
 sky130_fd_sc_hd__a21boi_4 _42276_ (.A1(_11365_),
    .A2(_11369_),
    .B1_N(_11367_),
    .Y(_11737_));
 sky130_fd_sc_hd__xnor2_4 _42277_ (.A(_11736_),
    .B(_11737_),
    .Y(_11738_));
 sky130_fd_sc_hd__nand2_4 _42278_ (.A(_11735_),
    .B(_11738_),
    .Y(_11739_));
 sky130_vsdinv _42279_ (.A(_11738_),
    .Y(_11740_));
 sky130_fd_sc_hd__nand3_4 _42280_ (.A(_11732_),
    .B(_11734_),
    .C(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__nand2_4 _42281_ (.A(_11739_),
    .B(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__nand2_4 _42282_ (.A(_11429_),
    .B(_11742_),
    .Y(_11743_));
 sky130_fd_sc_hd__nand3_4 _42283_ (.A(_11428_),
    .B(_11741_),
    .C(_11739_),
    .Y(_11744_));
 sky130_fd_sc_hd__nand2_4 _42284_ (.A(_11743_),
    .B(_11744_),
    .Y(_11745_));
 sky130_fd_sc_hd__a21boi_4 _42285_ (.A1(_11388_),
    .A2(_11383_),
    .B1_N(_11382_),
    .Y(_11746_));
 sky130_fd_sc_hd__nand2_4 _42286_ (.A(_11745_),
    .B(_11746_),
    .Y(_11747_));
 sky130_vsdinv _42287_ (.A(_11746_),
    .Y(_11748_));
 sky130_fd_sc_hd__nand3_4 _42288_ (.A(_11743_),
    .B(_11744_),
    .C(_11748_),
    .Y(_11749_));
 sky130_fd_sc_hd__nand2_4 _42289_ (.A(_11747_),
    .B(_11749_),
    .Y(_11750_));
 sky130_fd_sc_hd__a21oi_4 _42290_ (.A1(_11392_),
    .A2(_11394_),
    .B1(_11398_),
    .Y(_11751_));
 sky130_fd_sc_hd__o21ai_4 _42291_ (.A1(_11402_),
    .A2(_11751_),
    .B1(_11399_),
    .Y(_11752_));
 sky130_vsdinv _42292_ (.A(_11752_),
    .Y(_11753_));
 sky130_fd_sc_hd__nand2_4 _42293_ (.A(_11750_),
    .B(_11753_),
    .Y(_11754_));
 sky130_fd_sc_hd__nand3_4 _42294_ (.A(_11747_),
    .B(_11752_),
    .C(_11749_),
    .Y(_11755_));
 sky130_fd_sc_hd__nand2_4 _42295_ (.A(_11754_),
    .B(_11755_),
    .Y(_11756_));
 sky130_fd_sc_hd__a21boi_4 _42296_ (.A1(_11427_),
    .A2(_11407_),
    .B1_N(_11408_),
    .Y(_11757_));
 sky130_fd_sc_hd__xor2_4 _42297_ (.A(_11756_),
    .B(_11757_),
    .X(_01438_));
 sky130_fd_sc_hd__nand2_4 _42298_ (.A(_06384_),
    .B(_11433_),
    .Y(_11758_));
 sky130_fd_sc_hd__o21ai_4 _42299_ (.A1(_06133_),
    .A2(_11432_),
    .B1(_11758_),
    .Y(_11759_));
 sky130_fd_sc_hd__nand4_4 _42300_ (.A(_03254_),
    .B(_07196_),
    .C(_11438_),
    .D(_11107_),
    .Y(_11760_));
 sky130_fd_sc_hd__nand2_4 _42301_ (.A(_11759_),
    .B(_11760_),
    .Y(_11761_));
 sky130_fd_sc_hd__buf_1 _42302_ (.A(_10515_),
    .X(_11762_));
 sky130_fd_sc_hd__nand2_4 _42303_ (.A(_07365_),
    .B(_11762_),
    .Y(_11763_));
 sky130_fd_sc_hd__nand2_4 _42304_ (.A(_11761_),
    .B(_11763_),
    .Y(_11764_));
 sky130_vsdinv _42305_ (.A(_11763_),
    .Y(_11765_));
 sky130_fd_sc_hd__nand3_4 _42306_ (.A(_11759_),
    .B(_11765_),
    .C(_11760_),
    .Y(_11766_));
 sky130_fd_sc_hd__nand2_4 _42307_ (.A(_11764_),
    .B(_11766_),
    .Y(_11767_));
 sky130_fd_sc_hd__a21boi_4 _42308_ (.A1(_11435_),
    .A2(_11437_),
    .B1_N(_11439_),
    .Y(_11768_));
 sky130_fd_sc_hd__nand2_4 _42309_ (.A(_11767_),
    .B(_11768_),
    .Y(_11769_));
 sky130_fd_sc_hd__nand2_4 _42310_ (.A(_11440_),
    .B(_11439_),
    .Y(_11770_));
 sky130_fd_sc_hd__nand3_4 _42311_ (.A(_11770_),
    .B(_11766_),
    .C(_11764_),
    .Y(_11771_));
 sky130_fd_sc_hd__nand2_4 _42312_ (.A(_11769_),
    .B(_11771_),
    .Y(_11772_));
 sky130_fd_sc_hd__nand2_4 _42313_ (.A(_07938_),
    .B(_11447_),
    .Y(_11773_));
 sky130_fd_sc_hd__nand2_4 _42314_ (.A(_06163_),
    .B(_11449_),
    .Y(_11774_));
 sky130_fd_sc_hd__nand2_4 _42315_ (.A(_11773_),
    .B(_11774_),
    .Y(_11775_));
 sky130_fd_sc_hd__buf_1 _42316_ (.A(_10501_),
    .X(_11776_));
 sky130_fd_sc_hd__buf_1 _42317_ (.A(_03612_),
    .X(_11777_));
 sky130_fd_sc_hd__nand4_4 _42318_ (.A(_07526_),
    .B(_06163_),
    .C(_11776_),
    .D(_11777_),
    .Y(_11778_));
 sky130_fd_sc_hd__nand2_4 _42319_ (.A(_06155_),
    .B(_11125_),
    .Y(_11779_));
 sky130_vsdinv _42320_ (.A(_11779_),
    .Y(_11780_));
 sky130_fd_sc_hd__a21o_4 _42321_ (.A1(_11775_),
    .A2(_11778_),
    .B1(_11780_),
    .X(_11781_));
 sky130_fd_sc_hd__nand3_4 _42322_ (.A(_11775_),
    .B(_11778_),
    .C(_11780_),
    .Y(_11782_));
 sky130_fd_sc_hd__nand2_4 _42323_ (.A(_11781_),
    .B(_11782_),
    .Y(_11783_));
 sky130_fd_sc_hd__nand2_4 _42324_ (.A(_11772_),
    .B(_11783_),
    .Y(_11784_));
 sky130_vsdinv _42325_ (.A(_11783_),
    .Y(_11785_));
 sky130_fd_sc_hd__nand3_4 _42326_ (.A(_11769_),
    .B(_11785_),
    .C(_11771_),
    .Y(_11786_));
 sky130_fd_sc_hd__nand2_4 _42327_ (.A(_11784_),
    .B(_11786_),
    .Y(_11787_));
 sky130_fd_sc_hd__a21boi_4 _42328_ (.A1(_11459_),
    .A2(_11445_),
    .B1_N(_11443_),
    .Y(_11788_));
 sky130_fd_sc_hd__nand2_4 _42329_ (.A(_11787_),
    .B(_11788_),
    .Y(_11789_));
 sky130_fd_sc_hd__nand2_4 _42330_ (.A(_11460_),
    .B(_11443_),
    .Y(_11790_));
 sky130_fd_sc_hd__nand3_4 _42331_ (.A(_11790_),
    .B(_11784_),
    .C(_11786_),
    .Y(_11791_));
 sky130_fd_sc_hd__nand2_4 _42332_ (.A(_11789_),
    .B(_11791_),
    .Y(_11792_));
 sky130_fd_sc_hd__buf_1 _42333_ (.A(_09756_),
    .X(_11793_));
 sky130_fd_sc_hd__nand2_4 _42334_ (.A(_07762_),
    .B(_11793_),
    .Y(_11794_));
 sky130_fd_sc_hd__nand2_4 _42335_ (.A(_06451_),
    .B(_10922_),
    .Y(_11795_));
 sky130_fd_sc_hd__nand2_4 _42336_ (.A(_11794_),
    .B(_11795_),
    .Y(_11796_));
 sky130_fd_sc_hd__buf_1 _42337_ (.A(_09343_),
    .X(_11797_));
 sky130_fd_sc_hd__nand4_4 _42338_ (.A(_06550_),
    .B(_06564_),
    .C(_11797_),
    .D(_11142_),
    .Y(_11798_));
 sky130_fd_sc_hd__nand2_4 _42339_ (.A(_08394_),
    .B(_10927_),
    .Y(_11799_));
 sky130_vsdinv _42340_ (.A(_11799_),
    .Y(_11800_));
 sky130_fd_sc_hd__a21o_4 _42341_ (.A1(_11796_),
    .A2(_11798_),
    .B1(_11800_),
    .X(_11801_));
 sky130_fd_sc_hd__nand3_4 _42342_ (.A(_11796_),
    .B(_11798_),
    .C(_11800_),
    .Y(_11802_));
 sky130_fd_sc_hd__a21boi_4 _42343_ (.A1(_11451_),
    .A2(_11454_),
    .B1_N(_11452_),
    .Y(_11803_));
 sky130_fd_sc_hd__a21boi_4 _42344_ (.A1(_11801_),
    .A2(_11802_),
    .B1_N(_11803_),
    .Y(_11804_));
 sky130_vsdinv _42345_ (.A(_11804_),
    .Y(_11805_));
 sky130_vsdinv _42346_ (.A(_11803_),
    .Y(_11806_));
 sky130_fd_sc_hd__nand3_4 _42347_ (.A(_11806_),
    .B(_11801_),
    .C(_11802_),
    .Y(_11807_));
 sky130_fd_sc_hd__a21boi_4 _42348_ (.A1(_11471_),
    .A2(_11475_),
    .B1_N(_11472_),
    .Y(_11808_));
 sky130_vsdinv _42349_ (.A(_11808_),
    .Y(_11809_));
 sky130_fd_sc_hd__a21oi_4 _42350_ (.A1(_11805_),
    .A2(_11807_),
    .B1(_11809_),
    .Y(_11810_));
 sky130_fd_sc_hd__nand3_4 _42351_ (.A(_11805_),
    .B(_11809_),
    .C(_11807_),
    .Y(_11811_));
 sky130_vsdinv _42352_ (.A(_11811_),
    .Y(_11812_));
 sky130_fd_sc_hd__nor2_4 _42353_ (.A(_11810_),
    .B(_11812_),
    .Y(_11813_));
 sky130_vsdinv _42354_ (.A(_11813_),
    .Y(_11814_));
 sky130_fd_sc_hd__nand2_4 _42355_ (.A(_11792_),
    .B(_11814_),
    .Y(_11815_));
 sky130_fd_sc_hd__nand3_4 _42356_ (.A(_11813_),
    .B(_11789_),
    .C(_11791_),
    .Y(_11816_));
 sky130_fd_sc_hd__nand2_4 _42357_ (.A(_11815_),
    .B(_11816_),
    .Y(_11817_));
 sky130_fd_sc_hd__a21boi_4 _42358_ (.A1(_11458_),
    .A2(_11460_),
    .B1_N(_11463_),
    .Y(_11818_));
 sky130_fd_sc_hd__o21ai_4 _42359_ (.A1(_11487_),
    .A2(_11818_),
    .B1(_11466_),
    .Y(_11819_));
 sky130_vsdinv _42360_ (.A(_11819_),
    .Y(_11820_));
 sky130_fd_sc_hd__nand2_4 _42361_ (.A(_11817_),
    .B(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__nand3_4 _42362_ (.A(_11819_),
    .B(_11815_),
    .C(_11816_),
    .Y(_11822_));
 sky130_fd_sc_hd__nand2_4 _42363_ (.A(_11821_),
    .B(_11822_),
    .Y(_11823_));
 sky130_fd_sc_hd__buf_1 _42364_ (.A(_09313_),
    .X(_11824_));
 sky130_fd_sc_hd__nand2_4 _42365_ (.A(_10900_),
    .B(_11824_),
    .Y(_11825_));
 sky130_fd_sc_hd__buf_1 _42366_ (.A(_06711_),
    .X(_11826_));
 sky130_fd_sc_hd__nand2_4 _42367_ (.A(_11826_),
    .B(_08631_),
    .Y(_11827_));
 sky130_fd_sc_hd__nand2_4 _42368_ (.A(_11825_),
    .B(_11827_),
    .Y(_11828_));
 sky130_fd_sc_hd__buf_1 _42369_ (.A(_08630_),
    .X(_11829_));
 sky130_fd_sc_hd__nand4_4 _42370_ (.A(_07280_),
    .B(_11826_),
    .C(_11829_),
    .D(_11824_),
    .Y(_11830_));
 sky130_fd_sc_hd__nand2_4 _42371_ (.A(_07005_),
    .B(_10887_),
    .Y(_11831_));
 sky130_vsdinv _42372_ (.A(_11831_),
    .Y(_11832_));
 sky130_fd_sc_hd__a21o_4 _42373_ (.A1(_11828_),
    .A2(_11830_),
    .B1(_11832_),
    .X(_11833_));
 sky130_fd_sc_hd__nand3_4 _42374_ (.A(_11828_),
    .B(_11830_),
    .C(_11832_),
    .Y(_11834_));
 sky130_fd_sc_hd__nand2_4 _42375_ (.A(_11833_),
    .B(_11834_),
    .Y(_11835_));
 sky130_fd_sc_hd__a21o_4 _42376_ (.A1(_11504_),
    .A2(_11507_),
    .B1(_11835_),
    .X(_11836_));
 sky130_fd_sc_hd__nand3_4 _42377_ (.A(_11835_),
    .B(_11504_),
    .C(_11507_),
    .Y(_11837_));
 sky130_fd_sc_hd__nand2_4 _42378_ (.A(_11836_),
    .B(_11837_),
    .Y(_11838_));
 sky130_fd_sc_hd__nand2_4 _42379_ (.A(_11556_),
    .B(_03545_),
    .Y(_11839_));
 sky130_vsdinv _42380_ (.A(_11839_),
    .Y(_11840_));
 sky130_fd_sc_hd__nand2_4 _42381_ (.A(_07299_),
    .B(_11522_),
    .Y(_11841_));
 sky130_fd_sc_hd__buf_1 _42382_ (.A(_03552_),
    .X(_11842_));
 sky130_fd_sc_hd__nand2_4 _42383_ (.A(_07302_),
    .B(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__xnor2_4 _42384_ (.A(_11841_),
    .B(_11843_),
    .Y(_11844_));
 sky130_fd_sc_hd__xor2_4 _42385_ (.A(_11840_),
    .B(_11844_),
    .X(_11845_));
 sky130_fd_sc_hd__nand2_4 _42386_ (.A(_11838_),
    .B(_11845_),
    .Y(_11846_));
 sky130_fd_sc_hd__xor2_4 _42387_ (.A(_11839_),
    .B(_11844_),
    .X(_11847_));
 sky130_fd_sc_hd__nand3_4 _42388_ (.A(_11847_),
    .B(_11837_),
    .C(_11836_),
    .Y(_11848_));
 sky130_fd_sc_hd__a21oi_4 _42389_ (.A1(_11483_),
    .A2(_11482_),
    .B1(_11479_),
    .Y(_11849_));
 sky130_vsdinv _42390_ (.A(_11849_),
    .Y(_11850_));
 sky130_fd_sc_hd__a21o_4 _42391_ (.A1(_11846_),
    .A2(_11848_),
    .B1(_11850_),
    .X(_11851_));
 sky130_fd_sc_hd__nand3_4 _42392_ (.A(_11846_),
    .B(_11848_),
    .C(_11850_),
    .Y(_11852_));
 sky130_fd_sc_hd__a21boi_4 _42393_ (.A1(_11512_),
    .A2(_11526_),
    .B1_N(_11510_),
    .Y(_11853_));
 sky130_vsdinv _42394_ (.A(_11853_),
    .Y(_11854_));
 sky130_fd_sc_hd__a21o_4 _42395_ (.A1(_11851_),
    .A2(_11852_),
    .B1(_11854_),
    .X(_11855_));
 sky130_fd_sc_hd__nand3_4 _42396_ (.A(_11851_),
    .B(_11854_),
    .C(_11852_),
    .Y(_11856_));
 sky130_fd_sc_hd__nand2_4 _42397_ (.A(_11855_),
    .B(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__nand2_4 _42398_ (.A(_11823_),
    .B(_11857_),
    .Y(_11858_));
 sky130_fd_sc_hd__nand4_4 _42399_ (.A(_11856_),
    .B(_11821_),
    .C(_11855_),
    .D(_11822_),
    .Y(_11859_));
 sky130_fd_sc_hd__nand2_4 _42400_ (.A(_11858_),
    .B(_11859_),
    .Y(_11860_));
 sky130_fd_sc_hd__a21oi_4 _42401_ (.A1(_11488_),
    .A2(_11490_),
    .B1(_11493_),
    .Y(_11861_));
 sky130_fd_sc_hd__o21ai_4 _42402_ (.A1(_11540_),
    .A2(_11861_),
    .B1(_11496_),
    .Y(_11862_));
 sky130_vsdinv _42403_ (.A(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__nand2_4 _42404_ (.A(_11860_),
    .B(_11863_),
    .Y(_11864_));
 sky130_fd_sc_hd__nand3_4 _42405_ (.A(_11862_),
    .B(_11858_),
    .C(_11859_),
    .Y(_11865_));
 sky130_fd_sc_hd__nand2_4 _42406_ (.A(_11864_),
    .B(_11865_),
    .Y(_11866_));
 sky130_fd_sc_hd__maj3_4 _42407_ (.A(_11515_),
    .B(_11517_),
    .C(_11519_),
    .X(_11867_));
 sky130_fd_sc_hd__nand2_4 _42408_ (.A(_11014_),
    .B(_07557_),
    .Y(_11868_));
 sky130_fd_sc_hd__nand2_4 _42409_ (.A(_07630_),
    .B(_07554_),
    .Y(_11869_));
 sky130_fd_sc_hd__nand2_4 _42410_ (.A(_11868_),
    .B(_11869_),
    .Y(_11870_));
 sky130_fd_sc_hd__buf_1 _42411_ (.A(_08042_),
    .X(_11871_));
 sky130_fd_sc_hd__buf_1 _42412_ (.A(_08572_),
    .X(_11872_));
 sky130_fd_sc_hd__buf_1 _42413_ (.A(_07922_),
    .X(_11873_));
 sky130_fd_sc_hd__nand4_4 _42414_ (.A(_07627_),
    .B(_11871_),
    .C(_11872_),
    .D(_11873_),
    .Y(_11874_));
 sky130_fd_sc_hd__nand2_4 _42415_ (.A(_08307_),
    .B(_07563_),
    .Y(_11875_));
 sky130_vsdinv _42416_ (.A(_11875_),
    .Y(_11876_));
 sky130_fd_sc_hd__a21o_4 _42417_ (.A1(_11870_),
    .A2(_11874_),
    .B1(_11876_),
    .X(_11877_));
 sky130_fd_sc_hd__nand3_4 _42418_ (.A(_11870_),
    .B(_11874_),
    .C(_11876_),
    .Y(_11878_));
 sky130_fd_sc_hd__nand2_4 _42419_ (.A(_11877_),
    .B(_11878_),
    .Y(_11879_));
 sky130_fd_sc_hd__nor2_4 _42420_ (.A(_11867_),
    .B(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__nand2_4 _42421_ (.A(_11879_),
    .B(_11867_),
    .Y(_11881_));
 sky130_vsdinv _42422_ (.A(_11881_),
    .Y(_11882_));
 sky130_fd_sc_hd__a21boi_4 _42423_ (.A1(_11555_),
    .A2(_11561_),
    .B1_N(_11558_),
    .Y(_11883_));
 sky130_fd_sc_hd__o21ai_4 _42424_ (.A1(_11880_),
    .A2(_11882_),
    .B1(_11883_),
    .Y(_11884_));
 sky130_vsdinv _42425_ (.A(_11880_),
    .Y(_11885_));
 sky130_vsdinv _42426_ (.A(_11883_),
    .Y(_11886_));
 sky130_fd_sc_hd__nand3_4 _42427_ (.A(_11885_),
    .B(_11886_),
    .C(_11881_),
    .Y(_11887_));
 sky130_fd_sc_hd__a21oi_4 _42428_ (.A1(_11567_),
    .A2(_11569_),
    .B1(_11565_),
    .Y(_11888_));
 sky130_vsdinv _42429_ (.A(_11888_),
    .Y(_11889_));
 sky130_fd_sc_hd__a21o_4 _42430_ (.A1(_11884_),
    .A2(_11887_),
    .B1(_11889_),
    .X(_11890_));
 sky130_fd_sc_hd__nand3_4 _42431_ (.A(_11889_),
    .B(_11884_),
    .C(_11887_),
    .Y(_11891_));
 sky130_fd_sc_hd__nand2_4 _42432_ (.A(_11890_),
    .B(_11891_),
    .Y(_11892_));
 sky130_fd_sc_hd__buf_1 _42433_ (.A(_10703_),
    .X(_11893_));
 sky130_fd_sc_hd__nand2_4 _42434_ (.A(_11893_),
    .B(_06896_),
    .Y(_11894_));
 sky130_vsdinv _42435_ (.A(_11894_),
    .Y(_11895_));
 sky130_fd_sc_hd__nand2_4 _42436_ (.A(_10783_),
    .B(_07537_),
    .Y(_11896_));
 sky130_fd_sc_hd__nand2_4 _42437_ (.A(_11287_),
    .B(_06632_),
    .Y(_11897_));
 sky130_fd_sc_hd__nand2_4 _42438_ (.A(_11896_),
    .B(_11897_),
    .Y(_11898_));
 sky130_fd_sc_hd__nand4_4 _42439_ (.A(_10788_),
    .B(_10789_),
    .C(_07542_),
    .D(_07544_),
    .Y(_11899_));
 sky130_fd_sc_hd__nand2_4 _42440_ (.A(_11898_),
    .B(_11899_),
    .Y(_11900_));
 sky130_fd_sc_hd__xor2_4 _42441_ (.A(_11895_),
    .B(_11900_),
    .X(_11901_));
 sky130_fd_sc_hd__a21boi_4 _42442_ (.A1(_11581_),
    .A2(_11584_),
    .B1_N(_11582_),
    .Y(_11902_));
 sky130_vsdinv _42443_ (.A(_11902_),
    .Y(_11903_));
 sky130_fd_sc_hd__buf_8 _42444_ (.A(_10621_),
    .X(_11904_));
 sky130_fd_sc_hd__buf_1 _42445_ (.A(_07941_),
    .X(_11905_));
 sky130_fd_sc_hd__nand2_4 _42446_ (.A(_11904_),
    .B(_11905_),
    .Y(_11906_));
 sky130_fd_sc_hd__buf_8 _42447_ (.A(_03517_),
    .X(_11907_));
 sky130_fd_sc_hd__nand2_4 _42448_ (.A(_08749_),
    .B(_11907_),
    .Y(_11908_));
 sky130_fd_sc_hd__nand2_4 _42449_ (.A(_11906_),
    .B(_11908_),
    .Y(_11909_));
 sky130_fd_sc_hd__buf_1 _42450_ (.A(_11033_),
    .X(_11910_));
 sky130_fd_sc_hd__nand4_4 _42451_ (.A(_11910_),
    .B(_08754_),
    .C(_11907_),
    .D(_11905_),
    .Y(_11911_));
 sky130_fd_sc_hd__buf_1 _42452_ (.A(_10664_),
    .X(_11912_));
 sky130_fd_sc_hd__nand2_4 _42453_ (.A(_11912_),
    .B(_03513_),
    .Y(_11913_));
 sky130_fd_sc_hd__a21bo_4 _42454_ (.A1(_11909_),
    .A2(_11911_),
    .B1_N(_11913_),
    .X(_11914_));
 sky130_fd_sc_hd__buf_1 _42455_ (.A(_11912_),
    .X(_11915_));
 sky130_fd_sc_hd__nand4_4 _42456_ (.A(_11915_),
    .B(_11909_),
    .C(_11911_),
    .D(_03514_),
    .Y(_11916_));
 sky130_fd_sc_hd__nand2_4 _42457_ (.A(_11914_),
    .B(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__xor2_4 _42458_ (.A(_11903_),
    .B(_11917_),
    .X(_11918_));
 sky130_fd_sc_hd__xnor2_4 _42459_ (.A(_11901_),
    .B(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__nand2_4 _42460_ (.A(_11892_),
    .B(_11919_),
    .Y(_11920_));
 sky130_fd_sc_hd__xor2_4 _42461_ (.A(_11901_),
    .B(_11918_),
    .X(_11921_));
 sky130_fd_sc_hd__nand3_4 _42462_ (.A(_11921_),
    .B(_11890_),
    .C(_11891_),
    .Y(_11922_));
 sky130_fd_sc_hd__nand2_4 _42463_ (.A(_11920_),
    .B(_11922_),
    .Y(_11923_));
 sky130_fd_sc_hd__o21ai_4 _42464_ (.A1(_11535_),
    .A2(_11531_),
    .B1(_11532_),
    .Y(_11924_));
 sky130_vsdinv _42465_ (.A(_11924_),
    .Y(_11925_));
 sky130_fd_sc_hd__nand2_4 _42466_ (.A(_11923_),
    .B(_11925_),
    .Y(_11926_));
 sky130_fd_sc_hd__nand3_4 _42467_ (.A(_11920_),
    .B(_11922_),
    .C(_11924_),
    .Y(_11927_));
 sky130_fd_sc_hd__buf_1 _42468_ (.A(_11927_),
    .X(_11928_));
 sky130_fd_sc_hd__a21boi_4 _42469_ (.A1(_11574_),
    .A2(_11605_),
    .B1_N(_11576_),
    .Y(_11929_));
 sky130_vsdinv _42470_ (.A(_11929_),
    .Y(_11930_));
 sky130_fd_sc_hd__a21o_4 _42471_ (.A1(_11926_),
    .A2(_11928_),
    .B1(_11930_),
    .X(_11931_));
 sky130_fd_sc_hd__nand3_4 _42472_ (.A(_11926_),
    .B(_11930_),
    .C(_11927_),
    .Y(_11932_));
 sky130_fd_sc_hd__nand2_4 _42473_ (.A(_11931_),
    .B(_11932_),
    .Y(_11933_));
 sky130_fd_sc_hd__nand2_4 _42474_ (.A(_11866_),
    .B(_11933_),
    .Y(_11934_));
 sky130_fd_sc_hd__a21oi_4 _42475_ (.A1(_11926_),
    .A2(_11928_),
    .B1(_11930_),
    .Y(_11935_));
 sky130_vsdinv _42476_ (.A(_11932_),
    .Y(_11936_));
 sky130_fd_sc_hd__nor2_4 _42477_ (.A(_11935_),
    .B(_11936_),
    .Y(_11937_));
 sky130_fd_sc_hd__nand3_4 _42478_ (.A(_11937_),
    .B(_11865_),
    .C(_11864_),
    .Y(_11938_));
 sky130_fd_sc_hd__nand2_4 _42479_ (.A(_11934_),
    .B(_11938_),
    .Y(_11939_));
 sky130_fd_sc_hd__a21boi_4 _42480_ (.A1(_11623_),
    .A2(_11547_),
    .B1_N(_11549_),
    .Y(_11940_));
 sky130_fd_sc_hd__nand2_4 _42481_ (.A(_11939_),
    .B(_11940_),
    .Y(_11941_));
 sky130_fd_sc_hd__a21oi_4 _42482_ (.A1(_11541_),
    .A2(_11543_),
    .B1(_11548_),
    .Y(_11942_));
 sky130_fd_sc_hd__o21ai_4 _42483_ (.A1(_11619_),
    .A2(_11942_),
    .B1(_11549_),
    .Y(_11943_));
 sky130_fd_sc_hd__nand3_4 _42484_ (.A(_11943_),
    .B(_11938_),
    .C(_11934_),
    .Y(_11944_));
 sky130_fd_sc_hd__nand2_4 _42485_ (.A(_11941_),
    .B(_11944_),
    .Y(_11945_));
 sky130_fd_sc_hd__a21boi_4 _42486_ (.A1(_11655_),
    .A2(_11661_),
    .B1_N(_11657_),
    .Y(_11946_));
 sky130_vsdinv _42487_ (.A(_11946_),
    .Y(_11947_));
 sky130_fd_sc_hd__o21ai_4 _42488_ (.A1(_11589_),
    .A2(_11598_),
    .B1(_11602_),
    .Y(_11948_));
 sky130_fd_sc_hd__buf_1 _42489_ (.A(_10083_),
    .X(_11949_));
 sky130_fd_sc_hd__nand2_4 _42490_ (.A(_11949_),
    .B(_06794_),
    .Y(_11950_));
 sky130_fd_sc_hd__buf_1 _42491_ (.A(_10405_),
    .X(_11951_));
 sky130_fd_sc_hd__nand2_4 _42492_ (.A(_11951_),
    .B(_06377_),
    .Y(_11952_));
 sky130_fd_sc_hd__nand2_4 _42493_ (.A(_11950_),
    .B(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__buf_1 _42494_ (.A(_09847_),
    .X(_11954_));
 sky130_fd_sc_hd__buf_1 _42495_ (.A(_03383_),
    .X(_11955_));
 sky130_fd_sc_hd__nand4_4 _42496_ (.A(_11954_),
    .B(_11955_),
    .C(_03482_),
    .D(_06595_),
    .Y(_11956_));
 sky130_fd_sc_hd__buf_1 _42497_ (.A(_10406_),
    .X(_11957_));
 sky130_fd_sc_hd__nand2_4 _42498_ (.A(_11957_),
    .B(_06607_),
    .Y(_11958_));
 sky130_vsdinv _42499_ (.A(_11958_),
    .Y(_11959_));
 sky130_fd_sc_hd__a21o_4 _42500_ (.A1(_11953_),
    .A2(_11956_),
    .B1(_11959_),
    .X(_11960_));
 sky130_fd_sc_hd__nand3_4 _42501_ (.A(_11953_),
    .B(_11956_),
    .C(_11959_),
    .Y(_11961_));
 sky130_fd_sc_hd__nand2_4 _42502_ (.A(_11960_),
    .B(_11961_),
    .Y(_11962_));
 sky130_fd_sc_hd__nand2_4 _42503_ (.A(_11594_),
    .B(_11596_),
    .Y(_11963_));
 sky130_fd_sc_hd__nor2_4 _42504_ (.A(_11594_),
    .B(_11596_),
    .Y(_11964_));
 sky130_fd_sc_hd__a21oi_4 _42505_ (.A1(_11963_),
    .A2(_11592_),
    .B1(_11964_),
    .Y(_11965_));
 sky130_fd_sc_hd__nand2_4 _42506_ (.A(_11962_),
    .B(_11965_),
    .Y(_11966_));
 sky130_vsdinv _42507_ (.A(_11965_),
    .Y(_11967_));
 sky130_fd_sc_hd__nand3_4 _42508_ (.A(_11967_),
    .B(_11960_),
    .C(_11961_),
    .Y(_11968_));
 sky130_fd_sc_hd__a21boi_4 _42509_ (.A1(_11638_),
    .A2(_11644_),
    .B1_N(_11640_),
    .Y(_11969_));
 sky130_vsdinv _42510_ (.A(_11969_),
    .Y(_11970_));
 sky130_fd_sc_hd__nand3_4 _42511_ (.A(_11966_),
    .B(_11968_),
    .C(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__a21o_4 _42512_ (.A1(_11966_),
    .A2(_11968_),
    .B1(_11970_),
    .X(_11972_));
 sky130_fd_sc_hd__nand3_4 _42513_ (.A(_11948_),
    .B(_11971_),
    .C(_11972_),
    .Y(_11973_));
 sky130_fd_sc_hd__nand2_4 _42514_ (.A(_11972_),
    .B(_11971_),
    .Y(_11974_));
 sky130_fd_sc_hd__nand3_4 _42515_ (.A(_11974_),
    .B(_11602_),
    .C(_11603_),
    .Y(_11975_));
 sky130_fd_sc_hd__maj3_4 _42516_ (.A(_11649_),
    .B(_11647_),
    .C(_11633_),
    .X(_11976_));
 sky130_vsdinv _42517_ (.A(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__a21o_4 _42518_ (.A1(_11973_),
    .A2(_11975_),
    .B1(_11977_),
    .X(_11978_));
 sky130_fd_sc_hd__nand3_4 _42519_ (.A(_11973_),
    .B(_11975_),
    .C(_11977_),
    .Y(_11979_));
 sky130_fd_sc_hd__nand3_4 _42520_ (.A(_11947_),
    .B(_11978_),
    .C(_11979_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2_4 _42521_ (.A(_11978_),
    .B(_11979_),
    .Y(_11981_));
 sky130_fd_sc_hd__nand2_4 _42522_ (.A(_11981_),
    .B(_11946_),
    .Y(_11982_));
 sky130_fd_sc_hd__nand2_4 _42523_ (.A(_11980_),
    .B(_11982_),
    .Y(_11983_));
 sky130_fd_sc_hd__a21boi_4 _42524_ (.A1(_11672_),
    .A2(_11677_),
    .B1_N(_11674_),
    .Y(_11984_));
 sky130_fd_sc_hd__nand2_4 _42525_ (.A(_11673_),
    .B(_06229_),
    .Y(_11985_));
 sky130_fd_sc_hd__nand2_4 _42526_ (.A(_11675_),
    .B(_06228_),
    .Y(_11986_));
 sky130_fd_sc_hd__nand2_4 _42527_ (.A(_11985_),
    .B(_11986_),
    .Y(_11987_));
 sky130_fd_sc_hd__buf_1 _42528_ (.A(_10409_),
    .X(_11988_));
 sky130_fd_sc_hd__buf_1 _42529_ (.A(_10845_),
    .X(_11989_));
 sky130_fd_sc_hd__nand4_4 _42530_ (.A(_11988_),
    .B(_11989_),
    .C(_06321_),
    .D(_06323_),
    .Y(_11990_));
 sky130_fd_sc_hd__buf_1 _42531_ (.A(_11683_),
    .X(_11991_));
 sky130_fd_sc_hd__nand2_4 _42532_ (.A(_11991_),
    .B(_06551_),
    .Y(_11992_));
 sky130_vsdinv _42533_ (.A(_11992_),
    .Y(_11993_));
 sky130_fd_sc_hd__a21o_4 _42534_ (.A1(_11987_),
    .A2(_11990_),
    .B1(_11993_),
    .X(_11994_));
 sky130_fd_sc_hd__nand3_4 _42535_ (.A(_11987_),
    .B(_11990_),
    .C(_11993_),
    .Y(_11995_));
 sky130_fd_sc_hd__nand2_4 _42536_ (.A(_11994_),
    .B(_11995_),
    .Y(_11996_));
 sky130_fd_sc_hd__nor2_4 _42537_ (.A(_11984_),
    .B(_11996_),
    .Y(_11997_));
 sky130_vsdinv _42538_ (.A(_11997_),
    .Y(_11998_));
 sky130_fd_sc_hd__nand2_4 _42539_ (.A(_11996_),
    .B(_11984_),
    .Y(_11999_));
 sky130_fd_sc_hd__o21a_4 _42540_ (.A1(_03434_),
    .A2(_05938_),
    .B1(_11686_),
    .X(_12000_));
 sky130_fd_sc_hd__nand3_4 _42541_ (.A(_11691_),
    .B(_08047_),
    .C(_06080_),
    .Y(_12001_));
 sky130_fd_sc_hd__a21o_4 _42542_ (.A1(_12000_),
    .A2(_12001_),
    .B1(_11341_),
    .X(_12002_));
 sky130_fd_sc_hd__nand3_4 _42543_ (.A(_12000_),
    .B(_11341_),
    .C(_12001_),
    .Y(_12003_));
 sky130_fd_sc_hd__and2_4 _42544_ (.A(_12002_),
    .B(_12003_),
    .X(_12004_));
 sky130_fd_sc_hd__buf_1 _42545_ (.A(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__buf_1 _42546_ (.A(_12005_),
    .X(_12006_));
 sky130_fd_sc_hd__a21o_4 _42547_ (.A1(_11998_),
    .A2(_11999_),
    .B1(_12006_),
    .X(_12007_));
 sky130_fd_sc_hd__nand3_4 _42548_ (.A(_11998_),
    .B(_12006_),
    .C(_11999_),
    .Y(_12008_));
 sky130_fd_sc_hd__a21oi_4 _42549_ (.A1(_11698_),
    .A2(_11696_),
    .B1(_11681_),
    .Y(_12009_));
 sky130_vsdinv _42550_ (.A(_12009_),
    .Y(_12010_));
 sky130_fd_sc_hd__a21o_4 _42551_ (.A1(_12007_),
    .A2(_12008_),
    .B1(_12010_),
    .X(_12011_));
 sky130_fd_sc_hd__nand3_4 _42552_ (.A(_12010_),
    .B(_12007_),
    .C(_12008_),
    .Y(_12012_));
 sky130_fd_sc_hd__nand2_4 _42553_ (.A(_12011_),
    .B(_12012_),
    .Y(_12013_));
 sky130_fd_sc_hd__a21boi_4 _42554_ (.A1(_11689_),
    .A2(_11344_),
    .B1_N(_11693_),
    .Y(_12014_));
 sky130_fd_sc_hd__nand2_4 _42555_ (.A(_12013_),
    .B(_12014_),
    .Y(_12015_));
 sky130_vsdinv _42556_ (.A(_12014_),
    .Y(_12016_));
 sky130_fd_sc_hd__nand3_4 _42557_ (.A(_12011_),
    .B(_12016_),
    .C(_12012_),
    .Y(_12017_));
 sky130_fd_sc_hd__and2_4 _42558_ (.A(_12015_),
    .B(_12017_),
    .X(_12018_));
 sky130_vsdinv _42559_ (.A(_12018_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand2_4 _42560_ (.A(_11983_),
    .B(_12019_),
    .Y(_12020_));
 sky130_fd_sc_hd__nand3_4 _42561_ (.A(_12018_),
    .B(_11980_),
    .C(_11982_),
    .Y(_12021_));
 sky130_fd_sc_hd__nand2_4 _42562_ (.A(_12020_),
    .B(_12021_),
    .Y(_12022_));
 sky130_fd_sc_hd__a21oi_4 _42563_ (.A1(_11607_),
    .A2(_11608_),
    .B1(_11612_),
    .Y(_12023_));
 sky130_fd_sc_hd__o21ai_4 _42564_ (.A1(_11615_),
    .A2(_12023_),
    .B1(_11613_),
    .Y(_12024_));
 sky130_vsdinv _42565_ (.A(_12024_),
    .Y(_12025_));
 sky130_fd_sc_hd__nand2_4 _42566_ (.A(_12022_),
    .B(_12025_),
    .Y(_12026_));
 sky130_fd_sc_hd__nand3_4 _42567_ (.A(_12020_),
    .B(_12024_),
    .C(_12021_),
    .Y(_12027_));
 sky130_fd_sc_hd__buf_1 _42568_ (.A(_12027_),
    .X(_12028_));
 sky130_fd_sc_hd__nand2_4 _42569_ (.A(_12026_),
    .B(_12028_),
    .Y(_12029_));
 sky130_fd_sc_hd__a21boi_4 _42570_ (.A1(_11665_),
    .A2(_11711_),
    .B1_N(_11667_),
    .Y(_12030_));
 sky130_fd_sc_hd__nand2_4 _42571_ (.A(_12029_),
    .B(_12030_),
    .Y(_12031_));
 sky130_vsdinv _42572_ (.A(_12030_),
    .Y(_12032_));
 sky130_fd_sc_hd__nand3_4 _42573_ (.A(_12026_),
    .B(_12032_),
    .C(_12027_),
    .Y(_12033_));
 sky130_fd_sc_hd__nand2_4 _42574_ (.A(_12031_),
    .B(_12033_),
    .Y(_12034_));
 sky130_fd_sc_hd__nand2_4 _42575_ (.A(_11945_),
    .B(_12034_),
    .Y(_12035_));
 sky130_fd_sc_hd__a21oi_4 _42576_ (.A1(_12026_),
    .A2(_12028_),
    .B1(_12032_),
    .Y(_12036_));
 sky130_vsdinv _42577_ (.A(_12033_),
    .Y(_12037_));
 sky130_fd_sc_hd__nor2_4 _42578_ (.A(_12036_),
    .B(_12037_),
    .Y(_12038_));
 sky130_fd_sc_hd__nand3_4 _42579_ (.A(_12038_),
    .B(_11944_),
    .C(_11941_),
    .Y(_12039_));
 sky130_fd_sc_hd__nand2_4 _42580_ (.A(_12035_),
    .B(_12039_),
    .Y(_12040_));
 sky130_fd_sc_hd__a21oi_4 _42581_ (.A1(_11620_),
    .A2(_11624_),
    .B1(_11629_),
    .Y(_12041_));
 sky130_fd_sc_hd__o21a_4 _42582_ (.A1(_11725_),
    .A2(_12041_),
    .B1(_11630_),
    .X(_12042_));
 sky130_fd_sc_hd__nand2_4 _42583_ (.A(_12040_),
    .B(_12042_),
    .Y(_12043_));
 sky130_fd_sc_hd__o21ai_4 _42584_ (.A1(_11725_),
    .A2(_12041_),
    .B1(_11630_),
    .Y(_12044_));
 sky130_fd_sc_hd__nand3_4 _42585_ (.A(_12044_),
    .B(_12035_),
    .C(_12039_),
    .Y(_12045_));
 sky130_fd_sc_hd__nand2_4 _42586_ (.A(_12043_),
    .B(_12045_),
    .Y(_12046_));
 sky130_fd_sc_hd__maj3_4 _42587_ (.A(_11706_),
    .B(_11702_),
    .C(_11704_),
    .X(_12047_));
 sky130_fd_sc_hd__a21boi_4 _42588_ (.A1(_11717_),
    .A2(_11723_),
    .B1_N(_11719_),
    .Y(_12048_));
 sky130_fd_sc_hd__xnor2_4 _42589_ (.A(_12047_),
    .B(_12048_),
    .Y(_12049_));
 sky130_fd_sc_hd__nand2_4 _42590_ (.A(_12046_),
    .B(_12049_),
    .Y(_12050_));
 sky130_vsdinv _42591_ (.A(_12049_),
    .Y(_12051_));
 sky130_fd_sc_hd__nand3_4 _42592_ (.A(_12043_),
    .B(_12051_),
    .C(_12045_),
    .Y(_12052_));
 sky130_fd_sc_hd__nand2_4 _42593_ (.A(_12050_),
    .B(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__a21boi_4 _42594_ (.A1(_11732_),
    .A2(_11740_),
    .B1_N(_11734_),
    .Y(_12054_));
 sky130_fd_sc_hd__nand2_4 _42595_ (.A(_12053_),
    .B(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__nand2_4 _42596_ (.A(_11741_),
    .B(_11734_),
    .Y(_12056_));
 sky130_fd_sc_hd__nand3_4 _42597_ (.A(_12056_),
    .B(_12050_),
    .C(_12052_),
    .Y(_12057_));
 sky130_fd_sc_hd__nand2_4 _42598_ (.A(_12055_),
    .B(_12057_),
    .Y(_12058_));
 sky130_fd_sc_hd__a21oi_4 _42599_ (.A1(_11371_),
    .A2(_11367_),
    .B1(_11736_),
    .Y(_12059_));
 sky130_vsdinv _42600_ (.A(_12059_),
    .Y(_12060_));
 sky130_fd_sc_hd__nand2_4 _42601_ (.A(_12058_),
    .B(_12060_),
    .Y(_12061_));
 sky130_fd_sc_hd__nand3_4 _42602_ (.A(_12055_),
    .B(_12057_),
    .C(_12059_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_4 _42603_ (.A(_12061_),
    .B(_12062_),
    .Y(_12063_));
 sky130_fd_sc_hd__a21boi_4 _42604_ (.A1(_11743_),
    .A2(_11748_),
    .B1_N(_11744_),
    .Y(_12064_));
 sky130_fd_sc_hd__nand2_4 _42605_ (.A(_12063_),
    .B(_12064_),
    .Y(_12065_));
 sky130_fd_sc_hd__nand2_4 _42606_ (.A(_11749_),
    .B(_11744_),
    .Y(_12066_));
 sky130_fd_sc_hd__nand3_4 _42607_ (.A(_12066_),
    .B(_12062_),
    .C(_12061_),
    .Y(_12067_));
 sky130_fd_sc_hd__nand2_4 _42608_ (.A(_12065_),
    .B(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__nor2_4 _42609_ (.A(_11756_),
    .B(_11409_),
    .Y(_12069_));
 sky130_fd_sc_hd__nand2_4 _42610_ (.A(_11755_),
    .B(_11408_),
    .Y(_12070_));
 sky130_fd_sc_hd__nand2_4 _42611_ (.A(_12070_),
    .B(_11754_),
    .Y(_12071_));
 sky130_fd_sc_hd__a21boi_4 _42612_ (.A1(_11427_),
    .A2(_12069_),
    .B1_N(_12071_),
    .Y(_12072_));
 sky130_fd_sc_hd__xor2_4 _42613_ (.A(_12068_),
    .B(_12072_),
    .X(_01439_));
 sky130_fd_sc_hd__nand2_4 _42614_ (.A(_06010_),
    .B(_11102_),
    .Y(_12073_));
 sky130_fd_sc_hd__o21ai_4 _42615_ (.A1(_06008_),
    .A2(_03633_),
    .B1(_12073_),
    .Y(_12074_));
 sky130_fd_sc_hd__buf_1 _42616_ (.A(_03627_),
    .X(_12075_));
 sky130_fd_sc_hd__buf_1 _42617_ (.A(\pcpi_mul.rs2[32] ),
    .X(_12076_));
 sky130_fd_sc_hd__nand4_4 _42618_ (.A(_03257_),
    .B(_10480_),
    .C(_12075_),
    .D(_12076_),
    .Y(_12077_));
 sky130_fd_sc_hd__nand2_4 _42619_ (.A(_12074_),
    .B(_12077_),
    .Y(_12078_));
 sky130_fd_sc_hd__nand2_4 _42620_ (.A(_07736_),
    .B(_11762_),
    .Y(_12079_));
 sky130_fd_sc_hd__nand2_4 _42621_ (.A(_12078_),
    .B(_12079_),
    .Y(_12080_));
 sky130_vsdinv _42622_ (.A(_12079_),
    .Y(_12081_));
 sky130_fd_sc_hd__nand3_4 _42623_ (.A(_12074_),
    .B(_12081_),
    .C(_12077_),
    .Y(_12082_));
 sky130_fd_sc_hd__nand2_4 _42624_ (.A(_12080_),
    .B(_12082_),
    .Y(_12083_));
 sky130_fd_sc_hd__a21boi_4 _42625_ (.A1(_11759_),
    .A2(_11765_),
    .B1_N(_11760_),
    .Y(_12084_));
 sky130_fd_sc_hd__nand2_4 _42626_ (.A(_12083_),
    .B(_12084_),
    .Y(_12085_));
 sky130_fd_sc_hd__nand2_4 _42627_ (.A(_11766_),
    .B(_11760_),
    .Y(_12086_));
 sky130_fd_sc_hd__nand3_4 _42628_ (.A(_12086_),
    .B(_12082_),
    .C(_12080_),
    .Y(_12087_));
 sky130_fd_sc_hd__nand2_4 _42629_ (.A(_12085_),
    .B(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__nand2_4 _42630_ (.A(_06938_),
    .B(_03613_),
    .Y(_12089_));
 sky130_fd_sc_hd__nand2_4 _42631_ (.A(_06942_),
    .B(_03606_),
    .Y(_12090_));
 sky130_fd_sc_hd__nand2_4 _42632_ (.A(_12089_),
    .B(_12090_),
    .Y(_12091_));
 sky130_fd_sc_hd__buf_1 _42633_ (.A(_03605_),
    .X(_12092_));
 sky130_fd_sc_hd__buf_1 _42634_ (.A(_03612_),
    .X(_12093_));
 sky130_fd_sc_hd__nand4_4 _42635_ (.A(_06085_),
    .B(_06545_),
    .C(_12092_),
    .D(_12093_),
    .Y(_12094_));
 sky130_fd_sc_hd__buf_1 _42636_ (.A(_10035_),
    .X(_12095_));
 sky130_fd_sc_hd__nand2_4 _42637_ (.A(_06343_),
    .B(_12095_),
    .Y(_12096_));
 sky130_vsdinv _42638_ (.A(_12096_),
    .Y(_12097_));
 sky130_fd_sc_hd__a21o_4 _42639_ (.A1(_12091_),
    .A2(_12094_),
    .B1(_12097_),
    .X(_12098_));
 sky130_fd_sc_hd__nand3_4 _42640_ (.A(_12091_),
    .B(_12094_),
    .C(_12097_),
    .Y(_12099_));
 sky130_fd_sc_hd__and2_4 _42641_ (.A(_12098_),
    .B(_12099_),
    .X(_12100_));
 sky130_vsdinv _42642_ (.A(_12100_),
    .Y(_12101_));
 sky130_fd_sc_hd__nand2_4 _42643_ (.A(_12088_),
    .B(_12101_),
    .Y(_12102_));
 sky130_fd_sc_hd__nand3_4 _42644_ (.A(_12085_),
    .B(_12100_),
    .C(_12087_),
    .Y(_12103_));
 sky130_fd_sc_hd__nand2_4 _42645_ (.A(_12102_),
    .B(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__a21boi_4 _42646_ (.A1(_11769_),
    .A2(_11785_),
    .B1_N(_11771_),
    .Y(_12105_));
 sky130_fd_sc_hd__nand2_4 _42647_ (.A(_12104_),
    .B(_12105_),
    .Y(_12106_));
 sky130_fd_sc_hd__nand2_4 _42648_ (.A(_11786_),
    .B(_11771_),
    .Y(_12107_));
 sky130_fd_sc_hd__nand3_4 _42649_ (.A(_12107_),
    .B(_12103_),
    .C(_12102_),
    .Y(_12108_));
 sky130_fd_sc_hd__nand2_4 _42650_ (.A(_12106_),
    .B(_12108_),
    .Y(_12109_));
 sky130_fd_sc_hd__nand2_4 _42651_ (.A(_08168_),
    .B(_10925_),
    .Y(_12110_));
 sky130_fd_sc_hd__buf_1 _42652_ (.A(_09343_),
    .X(_12111_));
 sky130_fd_sc_hd__nand2_4 _42653_ (.A(_08169_),
    .B(_12111_),
    .Y(_12112_));
 sky130_fd_sc_hd__nand2_4 _42654_ (.A(_12110_),
    .B(_12112_),
    .Y(_12113_));
 sky130_fd_sc_hd__buf_1 _42655_ (.A(_10302_),
    .X(_12114_));
 sky130_fd_sc_hd__buf_1 _42656_ (.A(_10300_),
    .X(_12115_));
 sky130_fd_sc_hd__nand4_4 _42657_ (.A(_06980_),
    .B(_06833_),
    .C(_12114_),
    .D(_12115_),
    .Y(_12116_));
 sky130_fd_sc_hd__nand2_4 _42658_ (.A(_07130_),
    .B(_03582_),
    .Y(_12117_));
 sky130_vsdinv _42659_ (.A(_12117_),
    .Y(_12118_));
 sky130_fd_sc_hd__a21o_4 _42660_ (.A1(_12113_),
    .A2(_12116_),
    .B1(_12118_),
    .X(_12119_));
 sky130_fd_sc_hd__nand3_4 _42661_ (.A(_12113_),
    .B(_12116_),
    .C(_12118_),
    .Y(_12120_));
 sky130_fd_sc_hd__nand2_4 _42662_ (.A(_12119_),
    .B(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__a21boi_4 _42663_ (.A1(_11775_),
    .A2(_11780_),
    .B1_N(_11778_),
    .Y(_12122_));
 sky130_fd_sc_hd__nand2_4 _42664_ (.A(_12121_),
    .B(_12122_),
    .Y(_12123_));
 sky130_vsdinv _42665_ (.A(_12122_),
    .Y(_12124_));
 sky130_fd_sc_hd__nand3_4 _42666_ (.A(_12124_),
    .B(_12120_),
    .C(_12119_),
    .Y(_12125_));
 sky130_fd_sc_hd__a21boi_4 _42667_ (.A1(_11796_),
    .A2(_11800_),
    .B1_N(_11798_),
    .Y(_12126_));
 sky130_vsdinv _42668_ (.A(_12126_),
    .Y(_12127_));
 sky130_fd_sc_hd__a21o_4 _42669_ (.A1(_12123_),
    .A2(_12125_),
    .B1(_12127_),
    .X(_12128_));
 sky130_fd_sc_hd__nand3_4 _42670_ (.A(_12123_),
    .B(_12125_),
    .C(_12127_),
    .Y(_12129_));
 sky130_fd_sc_hd__and2_4 _42671_ (.A(_12128_),
    .B(_12129_),
    .X(_12130_));
 sky130_vsdinv _42672_ (.A(_12130_),
    .Y(_12131_));
 sky130_fd_sc_hd__nand2_4 _42673_ (.A(_12109_),
    .B(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__nand3_4 _42674_ (.A(_12106_),
    .B(_12130_),
    .C(_12108_),
    .Y(_12133_));
 sky130_fd_sc_hd__nand2_4 _42675_ (.A(_12132_),
    .B(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__a21boi_4 _42676_ (.A1(_11813_),
    .A2(_11789_),
    .B1_N(_11791_),
    .Y(_12135_));
 sky130_fd_sc_hd__nand2_4 _42677_ (.A(_12134_),
    .B(_12135_),
    .Y(_12136_));
 sky130_fd_sc_hd__nand2_4 _42678_ (.A(_11816_),
    .B(_11791_),
    .Y(_12137_));
 sky130_fd_sc_hd__nand3_4 _42679_ (.A(_12137_),
    .B(_12132_),
    .C(_12133_),
    .Y(_12138_));
 sky130_fd_sc_hd__nand2_4 _42680_ (.A(_12136_),
    .B(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__o21a_4 _42681_ (.A1(_11808_),
    .A2(_11804_),
    .B1(_11807_),
    .X(_12140_));
 sky130_vsdinv _42682_ (.A(_12140_),
    .Y(_12141_));
 sky130_fd_sc_hd__buf_1 _42683_ (.A(_03557_),
    .X(_12142_));
 sky130_fd_sc_hd__a2bb2o_4 _42684_ (.A1_N(_03326_),
    .A2_N(_03553_),
    .B1(_07158_),
    .B2(_12142_),
    .X(_12143_));
 sky130_fd_sc_hd__buf_1 _42685_ (.A(_08640_),
    .X(_12144_));
 sky130_fd_sc_hd__nand2_4 _42686_ (.A(_11557_),
    .B(_12144_),
    .Y(_12145_));
 sky130_vsdinv _42687_ (.A(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__nand4_4 _42688_ (.A(_07158_),
    .B(_11556_),
    .C(_11842_),
    .D(_12142_),
    .Y(_12147_));
 sky130_fd_sc_hd__nand3_4 _42689_ (.A(_12143_),
    .B(_12146_),
    .C(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__a21oi_4 _42690_ (.A1(_12143_),
    .A2(_12147_),
    .B1(_12146_),
    .Y(_12149_));
 sky130_vsdinv _42691_ (.A(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__a21boi_4 _42692_ (.A1(_11828_),
    .A2(_11832_),
    .B1_N(_11830_),
    .Y(_12151_));
 sky130_vsdinv _42693_ (.A(_12151_),
    .Y(_12152_));
 sky130_fd_sc_hd__nand2_4 _42694_ (.A(_06712_),
    .B(_10885_),
    .Y(_12153_));
 sky130_fd_sc_hd__nand2_4 _42695_ (.A(_08971_),
    .B(_10884_),
    .Y(_12154_));
 sky130_fd_sc_hd__nand2_4 _42696_ (.A(_12153_),
    .B(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__buf_1 _42697_ (.A(_10272_),
    .X(_12156_));
 sky130_fd_sc_hd__buf_1 _42698_ (.A(_10270_),
    .X(_12157_));
 sky130_fd_sc_hd__nand4_4 _42699_ (.A(_07416_),
    .B(_08971_),
    .C(_12156_),
    .D(_12157_),
    .Y(_12158_));
 sky130_fd_sc_hd__nand2_4 _42700_ (.A(_07422_),
    .B(_08635_),
    .Y(_12159_));
 sky130_vsdinv _42701_ (.A(_12159_),
    .Y(_12160_));
 sky130_fd_sc_hd__nand3_4 _42702_ (.A(_12155_),
    .B(_12158_),
    .C(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__a21o_4 _42703_ (.A1(_12155_),
    .A2(_12158_),
    .B1(_12160_),
    .X(_12162_));
 sky130_fd_sc_hd__nand3_4 _42704_ (.A(_12152_),
    .B(_12161_),
    .C(_12162_),
    .Y(_12163_));
 sky130_fd_sc_hd__nand2_4 _42705_ (.A(_12162_),
    .B(_12161_),
    .Y(_12164_));
 sky130_fd_sc_hd__nand2_4 _42706_ (.A(_12164_),
    .B(_12151_),
    .Y(_12165_));
 sky130_fd_sc_hd__nand4_4 _42707_ (.A(_12148_),
    .B(_12150_),
    .C(_12163_),
    .D(_12165_),
    .Y(_12166_));
 sky130_fd_sc_hd__nand2_4 _42708_ (.A(_12150_),
    .B(_12148_),
    .Y(_12167_));
 sky130_fd_sc_hd__nand2_4 _42709_ (.A(_12165_),
    .B(_12163_),
    .Y(_12168_));
 sky130_fd_sc_hd__nand2_4 _42710_ (.A(_12167_),
    .B(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__nand3_4 _42711_ (.A(_12141_),
    .B(_12166_),
    .C(_12169_),
    .Y(_12170_));
 sky130_fd_sc_hd__nand2_4 _42712_ (.A(_12169_),
    .B(_12166_),
    .Y(_12171_));
 sky130_fd_sc_hd__nand2_4 _42713_ (.A(_12171_),
    .B(_12140_),
    .Y(_12172_));
 sky130_fd_sc_hd__a21boi_4 _42714_ (.A1(_11847_),
    .A2(_11837_),
    .B1_N(_11836_),
    .Y(_12173_));
 sky130_vsdinv _42715_ (.A(_12173_),
    .Y(_12174_));
 sky130_fd_sc_hd__a21oi_4 _42716_ (.A1(_12170_),
    .A2(_12172_),
    .B1(_12174_),
    .Y(_12175_));
 sky130_fd_sc_hd__nand3_4 _42717_ (.A(_12170_),
    .B(_12172_),
    .C(_12174_),
    .Y(_12176_));
 sky130_vsdinv _42718_ (.A(_12176_),
    .Y(_12177_));
 sky130_fd_sc_hd__nor2_4 _42719_ (.A(_12175_),
    .B(_12177_),
    .Y(_12178_));
 sky130_vsdinv _42720_ (.A(_12178_),
    .Y(_12179_));
 sky130_fd_sc_hd__nand2_4 _42721_ (.A(_12139_),
    .B(_12179_),
    .Y(_12180_));
 sky130_fd_sc_hd__nand3_4 _42722_ (.A(_12136_),
    .B(_12178_),
    .C(_12138_),
    .Y(_12181_));
 sky130_fd_sc_hd__nand2_4 _42723_ (.A(_12180_),
    .B(_12181_),
    .Y(_12182_));
 sky130_fd_sc_hd__a21oi_4 _42724_ (.A1(_11815_),
    .A2(_11816_),
    .B1(_11819_),
    .Y(_12183_));
 sky130_fd_sc_hd__o21a_4 _42725_ (.A1(_12183_),
    .A2(_11857_),
    .B1(_11822_),
    .X(_12184_));
 sky130_fd_sc_hd__nand2_4 _42726_ (.A(_12182_),
    .B(_12184_),
    .Y(_12185_));
 sky130_fd_sc_hd__o21ai_4 _42727_ (.A1(_12183_),
    .A2(_11857_),
    .B1(_11822_),
    .Y(_12186_));
 sky130_fd_sc_hd__nand3_4 _42728_ (.A(_12186_),
    .B(_12180_),
    .C(_12181_),
    .Y(_12187_));
 sky130_fd_sc_hd__nand2_4 _42729_ (.A(_12185_),
    .B(_12187_),
    .Y(_12188_));
 sky130_fd_sc_hd__buf_1 _42730_ (.A(_08051_),
    .X(_12189_));
 sky130_fd_sc_hd__buf_1 _42731_ (.A(_08125_),
    .X(_12190_));
 sky130_fd_sc_hd__nand2_4 _42732_ (.A(_12189_),
    .B(_12190_),
    .Y(_12191_));
 sky130_fd_sc_hd__buf_1 _42733_ (.A(_07878_),
    .X(_12192_));
 sky130_fd_sc_hd__nand2_4 _42734_ (.A(_12192_),
    .B(_11872_),
    .Y(_12193_));
 sky130_fd_sc_hd__nand2_4 _42735_ (.A(_12191_),
    .B(_12193_),
    .Y(_12194_));
 sky130_fd_sc_hd__nand4_4 _42736_ (.A(_12189_),
    .B(_12192_),
    .C(_11872_),
    .D(_11873_),
    .Y(_12195_));
 sky130_fd_sc_hd__nand2_4 _42737_ (.A(_08526_),
    .B(_07337_),
    .Y(_12196_));
 sky130_vsdinv _42738_ (.A(_12196_),
    .Y(_12197_));
 sky130_fd_sc_hd__a21o_4 _42739_ (.A1(_12194_),
    .A2(_12195_),
    .B1(_12197_),
    .X(_12198_));
 sky130_fd_sc_hd__nand3_4 _42740_ (.A(_12194_),
    .B(_12195_),
    .C(_12197_),
    .Y(_12199_));
 sky130_fd_sc_hd__nand2_4 _42741_ (.A(_12198_),
    .B(_12199_),
    .Y(_12200_));
 sky130_fd_sc_hd__nand2_4 _42742_ (.A(_11841_),
    .B(_11843_),
    .Y(_12201_));
 sky130_fd_sc_hd__nor2_4 _42743_ (.A(_11841_),
    .B(_11843_),
    .Y(_12202_));
 sky130_fd_sc_hd__a21oi_4 _42744_ (.A1(_12201_),
    .A2(_11840_),
    .B1(_12202_),
    .Y(_12203_));
 sky130_fd_sc_hd__nand2_4 _42745_ (.A(_12200_),
    .B(_12203_),
    .Y(_12204_));
 sky130_vsdinv _42746_ (.A(_12203_),
    .Y(_12205_));
 sky130_fd_sc_hd__nand3_4 _42747_ (.A(_12205_),
    .B(_12199_),
    .C(_12198_),
    .Y(_12206_));
 sky130_fd_sc_hd__a21boi_4 _42748_ (.A1(_11870_),
    .A2(_11876_),
    .B1_N(_11874_),
    .Y(_12207_));
 sky130_vsdinv _42749_ (.A(_12207_),
    .Y(_12208_));
 sky130_fd_sc_hd__a21o_4 _42750_ (.A1(_12204_),
    .A2(_12206_),
    .B1(_12208_),
    .X(_12209_));
 sky130_fd_sc_hd__nand3_4 _42751_ (.A(_12204_),
    .B(_12206_),
    .C(_12208_),
    .Y(_12210_));
 sky130_fd_sc_hd__a21oi_4 _42752_ (.A1(_11881_),
    .A2(_11886_),
    .B1(_11880_),
    .Y(_12211_));
 sky130_vsdinv _42753_ (.A(_12211_),
    .Y(_12212_));
 sky130_fd_sc_hd__a21o_4 _42754_ (.A1(_12209_),
    .A2(_12210_),
    .B1(_12212_),
    .X(_12213_));
 sky130_fd_sc_hd__nand3_4 _42755_ (.A(_12212_),
    .B(_12210_),
    .C(_12209_),
    .Y(_12214_));
 sky130_fd_sc_hd__nand2_4 _42756_ (.A(_12213_),
    .B(_12214_),
    .Y(_12215_));
 sky130_fd_sc_hd__maj3_4 _42757_ (.A(_11906_),
    .B(_11913_),
    .C(_11908_),
    .X(_12216_));
 sky130_fd_sc_hd__nand2_4 _42758_ (.A(_08315_),
    .B(_07523_),
    .Y(_12217_));
 sky130_fd_sc_hd__nand2_4 _42759_ (.A(_08531_),
    .B(_07192_),
    .Y(_12218_));
 sky130_fd_sc_hd__nand2_4 _42760_ (.A(_12217_),
    .B(_12218_),
    .Y(_12219_));
 sky130_fd_sc_hd__buf_1 _42761_ (.A(_08748_),
    .X(_12220_));
 sky130_fd_sc_hd__buf_1 _42762_ (.A(_07362_),
    .X(_12221_));
 sky130_fd_sc_hd__nand4_4 _42763_ (.A(_12220_),
    .B(_03358_),
    .C(_03518_),
    .D(_12221_),
    .Y(_12222_));
 sky130_fd_sc_hd__nand2_4 _42764_ (.A(_08760_),
    .B(_06881_),
    .Y(_12223_));
 sky130_fd_sc_hd__a21bo_4 _42765_ (.A1(_12219_),
    .A2(_12222_),
    .B1_N(_12223_),
    .X(_12224_));
 sky130_fd_sc_hd__buf_1 _42766_ (.A(_09565_),
    .X(_12225_));
 sky130_fd_sc_hd__buf_1 _42767_ (.A(_12225_),
    .X(_12226_));
 sky130_fd_sc_hd__nand4_4 _42768_ (.A(_12226_),
    .B(_12219_),
    .C(_12222_),
    .D(_11023_),
    .Y(_12227_));
 sky130_fd_sc_hd__nand2_4 _42769_ (.A(_12224_),
    .B(_12227_),
    .Y(_12228_));
 sky130_fd_sc_hd__nor2_4 _42770_ (.A(_12216_),
    .B(_12228_),
    .Y(_12229_));
 sky130_fd_sc_hd__a21boi_4 _42771_ (.A1(_12227_),
    .A2(_12224_),
    .B1_N(_12216_),
    .Y(_12230_));
 sky130_fd_sc_hd__buf_1 _42772_ (.A(_09574_),
    .X(_12231_));
 sky130_fd_sc_hd__a2bb2o_4 _42773_ (.A1_N(_03377_),
    .A2_N(_03502_),
    .B1(_12231_),
    .B2(_07669_),
    .X(_12232_));
 sky130_fd_sc_hd__buf_1 _42774_ (.A(_11635_),
    .X(_12233_));
 sky130_fd_sc_hd__nand4_4 _42775_ (.A(_12231_),
    .B(_12233_),
    .C(_06892_),
    .D(_07038_),
    .Y(_12234_));
 sky130_fd_sc_hd__nand2_4 _42776_ (.A(_11954_),
    .B(_06896_),
    .Y(_12235_));
 sky130_vsdinv _42777_ (.A(_12235_),
    .Y(_12236_));
 sky130_fd_sc_hd__a21o_4 _42778_ (.A1(_12232_),
    .A2(_12234_),
    .B1(_12236_),
    .X(_12237_));
 sky130_fd_sc_hd__nand3_4 _42779_ (.A(_12232_),
    .B(_12236_),
    .C(_12234_),
    .Y(_12238_));
 sky130_fd_sc_hd__nand2_4 _42780_ (.A(_12237_),
    .B(_12238_),
    .Y(_12239_));
 sky130_fd_sc_hd__or3_4 _42781_ (.A(_12229_),
    .B(_12230_),
    .C(_12239_),
    .X(_12240_));
 sky130_fd_sc_hd__o21a_4 _42782_ (.A1(_12229_),
    .A2(_12230_),
    .B1(_12239_),
    .X(_12241_));
 sky130_vsdinv _42783_ (.A(_12241_),
    .Y(_12242_));
 sky130_fd_sc_hd__nand2_4 _42784_ (.A(_12240_),
    .B(_12242_),
    .Y(_12243_));
 sky130_fd_sc_hd__nand2_4 _42785_ (.A(_12215_),
    .B(_12243_),
    .Y(_12244_));
 sky130_fd_sc_hd__nand4_4 _42786_ (.A(_12240_),
    .B(_12213_),
    .C(_12242_),
    .D(_12214_),
    .Y(_12245_));
 sky130_fd_sc_hd__nand2_4 _42787_ (.A(_12244_),
    .B(_12245_),
    .Y(_12246_));
 sky130_fd_sc_hd__a21oi_4 _42788_ (.A1(_11846_),
    .A2(_11848_),
    .B1(_11850_),
    .Y(_12247_));
 sky130_fd_sc_hd__o21ai_4 _42789_ (.A1(_11853_),
    .A2(_12247_),
    .B1(_11852_),
    .Y(_12248_));
 sky130_vsdinv _42790_ (.A(_12248_),
    .Y(_12249_));
 sky130_fd_sc_hd__nand2_4 _42791_ (.A(_12246_),
    .B(_12249_),
    .Y(_12250_));
 sky130_fd_sc_hd__nand3_4 _42792_ (.A(_12248_),
    .B(_12244_),
    .C(_12245_),
    .Y(_12251_));
 sky130_fd_sc_hd__a21boi_4 _42793_ (.A1(_11921_),
    .A2(_11890_),
    .B1_N(_11891_),
    .Y(_12252_));
 sky130_vsdinv _42794_ (.A(_12252_),
    .Y(_12253_));
 sky130_fd_sc_hd__a21oi_4 _42795_ (.A1(_12250_),
    .A2(_12251_),
    .B1(_12253_),
    .Y(_12254_));
 sky130_vsdinv _42796_ (.A(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__nand3_4 _42797_ (.A(_12250_),
    .B(_12253_),
    .C(_12251_),
    .Y(_12256_));
 sky130_fd_sc_hd__nand2_4 _42798_ (.A(_12255_),
    .B(_12256_),
    .Y(_12257_));
 sky130_fd_sc_hd__nand2_4 _42799_ (.A(_12188_),
    .B(_12257_),
    .Y(_12258_));
 sky130_vsdinv _42800_ (.A(_12256_),
    .Y(_12259_));
 sky130_fd_sc_hd__nor2_4 _42801_ (.A(_12254_),
    .B(_12259_),
    .Y(_12260_));
 sky130_fd_sc_hd__nand3_4 _42802_ (.A(_12260_),
    .B(_12185_),
    .C(_12187_),
    .Y(_12261_));
 sky130_fd_sc_hd__nand2_4 _42803_ (.A(_12258_),
    .B(_12261_),
    .Y(_12262_));
 sky130_fd_sc_hd__a21boi_4 _42804_ (.A1(_11937_),
    .A2(_11864_),
    .B1_N(_11865_),
    .Y(_12263_));
 sky130_fd_sc_hd__nand2_4 _42805_ (.A(_12262_),
    .B(_12263_),
    .Y(_12264_));
 sky130_fd_sc_hd__a21oi_4 _42806_ (.A1(_11858_),
    .A2(_11859_),
    .B1(_11862_),
    .Y(_12265_));
 sky130_fd_sc_hd__o21ai_4 _42807_ (.A1(_12265_),
    .A2(_11933_),
    .B1(_11865_),
    .Y(_12266_));
 sky130_fd_sc_hd__nand3_4 _42808_ (.A(_12266_),
    .B(_12258_),
    .C(_12261_),
    .Y(_12267_));
 sky130_fd_sc_hd__nand2_4 _42809_ (.A(_12264_),
    .B(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__a21boi_4 _42810_ (.A1(_11914_),
    .A2(_11916_),
    .B1_N(_11902_),
    .Y(_12269_));
 sky130_fd_sc_hd__nand3_4 _42811_ (.A(_11903_),
    .B(_11914_),
    .C(_11916_),
    .Y(_12270_));
 sky130_fd_sc_hd__o21a_4 _42812_ (.A1(_11901_),
    .A2(_12269_),
    .B1(_12270_),
    .X(_12271_));
 sky130_vsdinv _42813_ (.A(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__buf_1 _42814_ (.A(_10405_),
    .X(_12273_));
 sky130_fd_sc_hd__nand2_4 _42815_ (.A(_12273_),
    .B(_06483_),
    .Y(_12274_));
 sky130_fd_sc_hd__nand2_4 _42816_ (.A(_11957_),
    .B(_07097_),
    .Y(_12275_));
 sky130_fd_sc_hd__nand2_4 _42817_ (.A(_12274_),
    .B(_12275_),
    .Y(_12276_));
 sky130_fd_sc_hd__buf_1 _42818_ (.A(_11317_),
    .X(_12277_));
 sky130_fd_sc_hd__buf_1 _42819_ (.A(_03387_),
    .X(_12278_));
 sky130_fd_sc_hd__buf_1 _42820_ (.A(_12278_),
    .X(_12279_));
 sky130_fd_sc_hd__nand4_4 _42821_ (.A(_12277_),
    .B(_12279_),
    .C(_06601_),
    .D(_06595_),
    .Y(_12280_));
 sky130_fd_sc_hd__nand2_4 _42822_ (.A(_10840_),
    .B(_06607_),
    .Y(_12281_));
 sky130_vsdinv _42823_ (.A(_12281_),
    .Y(_12282_));
 sky130_fd_sc_hd__a21o_4 _42824_ (.A1(_12276_),
    .A2(_12280_),
    .B1(_12282_),
    .X(_12283_));
 sky130_fd_sc_hd__nand3_4 _42825_ (.A(_12276_),
    .B(_12280_),
    .C(_12282_),
    .Y(_12284_));
 sky130_fd_sc_hd__nand2_4 _42826_ (.A(_12283_),
    .B(_12284_),
    .Y(_12285_));
 sky130_fd_sc_hd__a21boi_4 _42827_ (.A1(_11898_),
    .A2(_11895_),
    .B1_N(_11899_),
    .Y(_12286_));
 sky130_fd_sc_hd__nand2_4 _42828_ (.A(_12285_),
    .B(_12286_),
    .Y(_12287_));
 sky130_vsdinv _42829_ (.A(_12286_),
    .Y(_12288_));
 sky130_fd_sc_hd__nand3_4 _42830_ (.A(_12288_),
    .B(_12283_),
    .C(_12284_),
    .Y(_12289_));
 sky130_fd_sc_hd__a21boi_4 _42831_ (.A1(_11953_),
    .A2(_11959_),
    .B1_N(_11956_),
    .Y(_12290_));
 sky130_vsdinv _42832_ (.A(_12290_),
    .Y(_12291_));
 sky130_fd_sc_hd__nand3_4 _42833_ (.A(_12287_),
    .B(_12289_),
    .C(_12291_),
    .Y(_12292_));
 sky130_fd_sc_hd__a21o_4 _42834_ (.A1(_12287_),
    .A2(_12289_),
    .B1(_12291_),
    .X(_12293_));
 sky130_fd_sc_hd__nand3_4 _42835_ (.A(_12272_),
    .B(_12292_),
    .C(_12293_),
    .Y(_12294_));
 sky130_fd_sc_hd__nand2_4 _42836_ (.A(_12293_),
    .B(_12292_),
    .Y(_12295_));
 sky130_fd_sc_hd__nand2_4 _42837_ (.A(_12295_),
    .B(_12271_),
    .Y(_12296_));
 sky130_fd_sc_hd__a21boi_4 _42838_ (.A1(_11966_),
    .A2(_11970_),
    .B1_N(_11968_),
    .Y(_12297_));
 sky130_vsdinv _42839_ (.A(_12297_),
    .Y(_12298_));
 sky130_fd_sc_hd__a21o_4 _42840_ (.A1(_12294_),
    .A2(_12296_),
    .B1(_12298_),
    .X(_12299_));
 sky130_fd_sc_hd__nand3_4 _42841_ (.A(_12294_),
    .B(_12296_),
    .C(_12298_),
    .Y(_12300_));
 sky130_fd_sc_hd__nand2_4 _42842_ (.A(_12299_),
    .B(_12300_),
    .Y(_12301_));
 sky130_fd_sc_hd__a21boi_4 _42843_ (.A1(_11977_),
    .A2(_11975_),
    .B1_N(_11973_),
    .Y(_12302_));
 sky130_fd_sc_hd__nand2_4 _42844_ (.A(_12301_),
    .B(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__nand2_4 _42845_ (.A(_11979_),
    .B(_11973_),
    .Y(_12304_));
 sky130_fd_sc_hd__nand3_4 _42846_ (.A(_12304_),
    .B(_12299_),
    .C(_12300_),
    .Y(_12305_));
 sky130_fd_sc_hd__nand2_4 _42847_ (.A(_12303_),
    .B(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__a21boi_4 _42848_ (.A1(_11987_),
    .A2(_11993_),
    .B1_N(_11990_),
    .Y(_12307_));
 sky130_fd_sc_hd__buf_1 _42849_ (.A(_11333_),
    .X(_12308_));
 sky130_fd_sc_hd__nand2_4 _42850_ (.A(_12308_),
    .B(_06128_),
    .Y(_12309_));
 sky130_fd_sc_hd__buf_1 _42851_ (.A(_11683_),
    .X(_12310_));
 sky130_fd_sc_hd__nand2_4 _42852_ (.A(_12310_),
    .B(_06130_),
    .Y(_12311_));
 sky130_fd_sc_hd__nand2_4 _42853_ (.A(_12309_),
    .B(_12311_),
    .Y(_12312_));
 sky130_fd_sc_hd__buf_1 _42854_ (.A(_11683_),
    .X(_12313_));
 sky130_fd_sc_hd__nand4_4 _42855_ (.A(_10846_),
    .B(_12313_),
    .C(_07132_),
    .D(_07128_),
    .Y(_12314_));
 sky130_fd_sc_hd__buf_1 _42856_ (.A(\pcpi_mul.rs1[32] ),
    .X(_12315_));
 sky130_fd_sc_hd__nand2_4 _42857_ (.A(_12315_),
    .B(_06231_),
    .Y(_12316_));
 sky130_vsdinv _42858_ (.A(_12316_),
    .Y(_12317_));
 sky130_fd_sc_hd__buf_1 _42859_ (.A(_12317_),
    .X(_12318_));
 sky130_fd_sc_hd__a21o_4 _42860_ (.A1(_12312_),
    .A2(_12314_),
    .B1(_12318_),
    .X(_12319_));
 sky130_fd_sc_hd__nand3_4 _42861_ (.A(_12312_),
    .B(_12314_),
    .C(_12318_),
    .Y(_12320_));
 sky130_fd_sc_hd__nand2_4 _42862_ (.A(_12319_),
    .B(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__nor2_4 _42863_ (.A(_12307_),
    .B(_12321_),
    .Y(_12322_));
 sky130_vsdinv _42864_ (.A(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__nand2_4 _42865_ (.A(_12321_),
    .B(_12307_),
    .Y(_12324_));
 sky130_fd_sc_hd__buf_1 _42866_ (.A(_12005_),
    .X(_12325_));
 sky130_fd_sc_hd__a21o_4 _42867_ (.A1(_12323_),
    .A2(_12324_),
    .B1(_12325_),
    .X(_12326_));
 sky130_fd_sc_hd__nand3_4 _42868_ (.A(_12323_),
    .B(_12325_),
    .C(_12324_),
    .Y(_12327_));
 sky130_fd_sc_hd__nand2_4 _42869_ (.A(_12326_),
    .B(_12327_),
    .Y(_12328_));
 sky130_fd_sc_hd__a21oi_4 _42870_ (.A1(_12325_),
    .A2(_11999_),
    .B1(_11997_),
    .Y(_12329_));
 sky130_fd_sc_hd__nand2_4 _42871_ (.A(_12328_),
    .B(_12329_),
    .Y(_12330_));
 sky130_vsdinv _42872_ (.A(_12329_),
    .Y(_12331_));
 sky130_fd_sc_hd__nand3_4 _42873_ (.A(_12326_),
    .B(_12327_),
    .C(_12331_),
    .Y(_12332_));
 sky130_fd_sc_hd__a21boi_4 _42874_ (.A1(_12000_),
    .A2(_11344_),
    .B1_N(_12001_),
    .Y(_12333_));
 sky130_vsdinv _42875_ (.A(_12333_),
    .Y(_12334_));
 sky130_fd_sc_hd__buf_1 _42876_ (.A(_12334_),
    .X(_12335_));
 sky130_fd_sc_hd__a21oi_4 _42877_ (.A1(_12330_),
    .A2(_12332_),
    .B1(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__buf_1 _42878_ (.A(_12334_),
    .X(_12337_));
 sky130_fd_sc_hd__nand3_4 _42879_ (.A(_12330_),
    .B(_12337_),
    .C(_12332_),
    .Y(_12338_));
 sky130_vsdinv _42880_ (.A(_12338_),
    .Y(_12339_));
 sky130_fd_sc_hd__nor2_4 _42881_ (.A(_12336_),
    .B(_12339_),
    .Y(_12340_));
 sky130_vsdinv _42882_ (.A(_12340_),
    .Y(_12341_));
 sky130_fd_sc_hd__nand2_4 _42883_ (.A(_12306_),
    .B(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__nand3_4 _42884_ (.A(_12303_),
    .B(_12340_),
    .C(_12305_),
    .Y(_12343_));
 sky130_fd_sc_hd__nand2_4 _42885_ (.A(_12342_),
    .B(_12343_),
    .Y(_12344_));
 sky130_fd_sc_hd__a21boi_4 _42886_ (.A1(_11926_),
    .A2(_11930_),
    .B1_N(_11928_),
    .Y(_12345_));
 sky130_fd_sc_hd__nand2_4 _42887_ (.A(_12344_),
    .B(_12345_),
    .Y(_12346_));
 sky130_fd_sc_hd__a21oi_4 _42888_ (.A1(_11920_),
    .A2(_11922_),
    .B1(_11924_),
    .Y(_12347_));
 sky130_fd_sc_hd__o21ai_4 _42889_ (.A1(_11929_),
    .A2(_12347_),
    .B1(_11928_),
    .Y(_12348_));
 sky130_fd_sc_hd__nand3_4 _42890_ (.A(_12348_),
    .B(_12342_),
    .C(_12343_),
    .Y(_12349_));
 sky130_fd_sc_hd__a21boi_4 _42891_ (.A1(_12018_),
    .A2(_11982_),
    .B1_N(_11980_),
    .Y(_12350_));
 sky130_vsdinv _42892_ (.A(_12350_),
    .Y(_12351_));
 sky130_fd_sc_hd__a21oi_4 _42893_ (.A1(_12346_),
    .A2(_12349_),
    .B1(_12351_),
    .Y(_12352_));
 sky130_vsdinv _42894_ (.A(_12352_),
    .Y(_12353_));
 sky130_fd_sc_hd__nand3_4 _42895_ (.A(_12346_),
    .B(_12351_),
    .C(_12349_),
    .Y(_12354_));
 sky130_fd_sc_hd__nand2_4 _42896_ (.A(_12353_),
    .B(_12354_),
    .Y(_12355_));
 sky130_fd_sc_hd__nand2_4 _42897_ (.A(_12268_),
    .B(_12355_),
    .Y(_12356_));
 sky130_vsdinv _42898_ (.A(_12354_),
    .Y(_12357_));
 sky130_fd_sc_hd__nor2_4 _42899_ (.A(_12352_),
    .B(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__nand3_4 _42900_ (.A(_12358_),
    .B(_12264_),
    .C(_12267_),
    .Y(_12359_));
 sky130_fd_sc_hd__nand2_4 _42901_ (.A(_12356_),
    .B(_12359_),
    .Y(_12360_));
 sky130_fd_sc_hd__a21boi_4 _42902_ (.A1(_12038_),
    .A2(_11941_),
    .B1_N(_11944_),
    .Y(_12361_));
 sky130_fd_sc_hd__nand2_4 _42903_ (.A(_12360_),
    .B(_12361_),
    .Y(_12362_));
 sky130_fd_sc_hd__a21oi_4 _42904_ (.A1(_11934_),
    .A2(_11938_),
    .B1(_11943_),
    .Y(_12363_));
 sky130_fd_sc_hd__o21ai_4 _42905_ (.A1(_12034_),
    .A2(_12363_),
    .B1(_11944_),
    .Y(_12364_));
 sky130_fd_sc_hd__nand3_4 _42906_ (.A(_12364_),
    .B(_12356_),
    .C(_12359_),
    .Y(_12365_));
 sky130_fd_sc_hd__nand2_4 _42907_ (.A(_12362_),
    .B(_12365_),
    .Y(_12366_));
 sky130_fd_sc_hd__a21boi_4 _42908_ (.A1(_12011_),
    .A2(_12016_),
    .B1_N(_12012_),
    .Y(_12367_));
 sky130_fd_sc_hd__a21boi_4 _42909_ (.A1(_12026_),
    .A2(_12032_),
    .B1_N(_12028_),
    .Y(_12368_));
 sky130_fd_sc_hd__xnor2_4 _42910_ (.A(_12367_),
    .B(_12368_),
    .Y(_12369_));
 sky130_fd_sc_hd__nand2_4 _42911_ (.A(_12366_),
    .B(_12369_),
    .Y(_12370_));
 sky130_vsdinv _42912_ (.A(_12369_),
    .Y(_12371_));
 sky130_fd_sc_hd__nand3_4 _42913_ (.A(_12362_),
    .B(_12365_),
    .C(_12371_),
    .Y(_12372_));
 sky130_fd_sc_hd__nand2_4 _42914_ (.A(_12370_),
    .B(_12372_),
    .Y(_12373_));
 sky130_fd_sc_hd__a21boi_4 _42915_ (.A1(_12043_),
    .A2(_12051_),
    .B1_N(_12045_),
    .Y(_12374_));
 sky130_fd_sc_hd__nand2_4 _42916_ (.A(_12373_),
    .B(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__nand2_4 _42917_ (.A(_12052_),
    .B(_12045_),
    .Y(_12376_));
 sky130_fd_sc_hd__nand3_4 _42918_ (.A(_12376_),
    .B(_12370_),
    .C(_12372_),
    .Y(_12377_));
 sky130_fd_sc_hd__nand2_4 _42919_ (.A(_12375_),
    .B(_12377_),
    .Y(_12378_));
 sky130_fd_sc_hd__a21oi_4 _42920_ (.A1(_11724_),
    .A2(_11719_),
    .B1(_12047_),
    .Y(_12379_));
 sky130_vsdinv _42921_ (.A(_12379_),
    .Y(_12380_));
 sky130_fd_sc_hd__nand2_4 _42922_ (.A(_12378_),
    .B(_12380_),
    .Y(_12381_));
 sky130_fd_sc_hd__nand3_4 _42923_ (.A(_12375_),
    .B(_12377_),
    .C(_12379_),
    .Y(_12382_));
 sky130_fd_sc_hd__nand2_4 _42924_ (.A(_12381_),
    .B(_12382_),
    .Y(_12383_));
 sky130_fd_sc_hd__a21boi_4 _42925_ (.A1(_12055_),
    .A2(_12059_),
    .B1_N(_12057_),
    .Y(_12384_));
 sky130_fd_sc_hd__nand2_4 _42926_ (.A(_12383_),
    .B(_12384_),
    .Y(_12385_));
 sky130_fd_sc_hd__nand2_4 _42927_ (.A(_12062_),
    .B(_12057_),
    .Y(_12386_));
 sky130_fd_sc_hd__nand3_4 _42928_ (.A(_12386_),
    .B(_12382_),
    .C(_12381_),
    .Y(_12387_));
 sky130_fd_sc_hd__nand2_4 _42929_ (.A(_12385_),
    .B(_12387_),
    .Y(_12388_));
 sky130_fd_sc_hd__o21ai_4 _42930_ (.A1(_12068_),
    .A2(_12072_),
    .B1(_12067_),
    .Y(_12389_));
 sky130_fd_sc_hd__xnor2_4 _42931_ (.A(_12388_),
    .B(_12389_),
    .Y(_01440_));
 sky130_fd_sc_hd__buf_1 _42932_ (.A(\pcpi_mul.rs2[31] ),
    .X(_12390_));
 sky130_fd_sc_hd__nand2_4 _42933_ (.A(_07736_),
    .B(_12390_),
    .Y(_12391_));
 sky130_fd_sc_hd__o21ai_4 _42934_ (.A1(_06142_),
    .A2(_11101_),
    .B1(_12391_),
    .Y(_12392_));
 sky130_fd_sc_hd__buf_1 _42935_ (.A(\pcpi_mul.rs2[32] ),
    .X(_12393_));
 sky130_fd_sc_hd__nand4_4 _42936_ (.A(_03262_),
    .B(_07736_),
    .C(_03628_),
    .D(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__nand2_4 _42937_ (.A(_12392_),
    .B(_12394_),
    .Y(_12395_));
 sky130_fd_sc_hd__nand2_4 _42938_ (.A(_06169_),
    .B(_03619_),
    .Y(_12396_));
 sky130_fd_sc_hd__nand2_4 _42939_ (.A(_12395_),
    .B(_12396_),
    .Y(_12397_));
 sky130_vsdinv _42940_ (.A(_12396_),
    .Y(_12398_));
 sky130_fd_sc_hd__nand3_4 _42941_ (.A(_12392_),
    .B(_12398_),
    .C(_12394_),
    .Y(_12399_));
 sky130_fd_sc_hd__nand2_4 _42942_ (.A(_12082_),
    .B(_12077_),
    .Y(_12400_));
 sky130_fd_sc_hd__a21o_4 _42943_ (.A1(_12397_),
    .A2(_12399_),
    .B1(_12400_),
    .X(_12401_));
 sky130_fd_sc_hd__nand3_4 _42944_ (.A(_12400_),
    .B(_12399_),
    .C(_12397_),
    .Y(_12402_));
 sky130_fd_sc_hd__nand2_4 _42945_ (.A(_12401_),
    .B(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__buf_1 _42946_ (.A(_10324_),
    .X(_12404_));
 sky130_fd_sc_hd__nand2_4 _42947_ (.A(_06945_),
    .B(_12404_),
    .Y(_12405_));
 sky130_fd_sc_hd__buf_1 _42948_ (.A(_10322_),
    .X(_12406_));
 sky130_fd_sc_hd__nand2_4 _42949_ (.A(_06550_),
    .B(_12406_),
    .Y(_12407_));
 sky130_fd_sc_hd__nand2_4 _42950_ (.A(_12405_),
    .B(_12407_),
    .Y(_12408_));
 sky130_fd_sc_hd__buf_1 _42951_ (.A(_10946_),
    .X(_12409_));
 sky130_fd_sc_hd__buf_1 _42952_ (.A(_10947_),
    .X(_12410_));
 sky130_fd_sc_hd__nand4_4 _42953_ (.A(_06252_),
    .B(_06444_),
    .C(_12409_),
    .D(_12410_),
    .Y(_12411_));
 sky130_fd_sc_hd__nand2_4 _42954_ (.A(_06980_),
    .B(_10512_),
    .Y(_12412_));
 sky130_vsdinv _42955_ (.A(_12412_),
    .Y(_12413_));
 sky130_fd_sc_hd__a21o_4 _42956_ (.A1(_12408_),
    .A2(_12411_),
    .B1(_12413_),
    .X(_12414_));
 sky130_fd_sc_hd__nand3_4 _42957_ (.A(_12408_),
    .B(_12411_),
    .C(_12413_),
    .Y(_12415_));
 sky130_fd_sc_hd__nand2_4 _42958_ (.A(_12414_),
    .B(_12415_),
    .Y(_12416_));
 sky130_fd_sc_hd__nand2_4 _42959_ (.A(_12403_),
    .B(_12416_),
    .Y(_12417_));
 sky130_vsdinv _42960_ (.A(_12416_),
    .Y(_12418_));
 sky130_fd_sc_hd__nand3_4 _42961_ (.A(_12401_),
    .B(_12418_),
    .C(_12402_),
    .Y(_12419_));
 sky130_fd_sc_hd__nand2_4 _42962_ (.A(_12417_),
    .B(_12419_),
    .Y(_12420_));
 sky130_fd_sc_hd__a21boi_4 _42963_ (.A1(_12085_),
    .A2(_12100_),
    .B1_N(_12087_),
    .Y(_12421_));
 sky130_fd_sc_hd__nand2_4 _42964_ (.A(_12420_),
    .B(_12421_),
    .Y(_12422_));
 sky130_vsdinv _42965_ (.A(_12421_),
    .Y(_12423_));
 sky130_fd_sc_hd__nand3_4 _42966_ (.A(_12423_),
    .B(_12419_),
    .C(_12417_),
    .Y(_12424_));
 sky130_fd_sc_hd__nand2_4 _42967_ (.A(_12422_),
    .B(_12424_),
    .Y(_12425_));
 sky130_fd_sc_hd__nand2_4 _42968_ (.A(_08169_),
    .B(_03596_),
    .Y(_12426_));
 sky130_fd_sc_hd__buf_1 _42969_ (.A(_09760_),
    .X(_12427_));
 sky130_fd_sc_hd__nand2_4 _42970_ (.A(_10900_),
    .B(_12427_),
    .Y(_12428_));
 sky130_fd_sc_hd__nand2_4 _42971_ (.A(_12426_),
    .B(_12428_),
    .Y(_12429_));
 sky130_fd_sc_hd__buf_1 _42972_ (.A(_10302_),
    .X(_12430_));
 sky130_fd_sc_hd__buf_1 _42973_ (.A(_10476_),
    .X(_12431_));
 sky130_fd_sc_hd__nand4_4 _42974_ (.A(_06833_),
    .B(_07284_),
    .C(_12430_),
    .D(_12431_),
    .Y(_12432_));
 sky130_fd_sc_hd__nand2_4 _42975_ (.A(_08835_),
    .B(_09347_),
    .Y(_12433_));
 sky130_vsdinv _42976_ (.A(_12433_),
    .Y(_12434_));
 sky130_fd_sc_hd__a21o_4 _42977_ (.A1(_12429_),
    .A2(_12432_),
    .B1(_12434_),
    .X(_12435_));
 sky130_fd_sc_hd__nand3_4 _42978_ (.A(_12429_),
    .B(_12432_),
    .C(_12434_),
    .Y(_12436_));
 sky130_fd_sc_hd__nand2_4 _42979_ (.A(_12435_),
    .B(_12436_),
    .Y(_12437_));
 sky130_fd_sc_hd__a21o_4 _42980_ (.A1(_12094_),
    .A2(_12099_),
    .B1(_12437_),
    .X(_12438_));
 sky130_fd_sc_hd__a21boi_4 _42981_ (.A1(_12091_),
    .A2(_12097_),
    .B1_N(_12094_),
    .Y(_12439_));
 sky130_fd_sc_hd__nand2_4 _42982_ (.A(_12437_),
    .B(_12439_),
    .Y(_12440_));
 sky130_fd_sc_hd__nand2_4 _42983_ (.A(_12438_),
    .B(_12440_),
    .Y(_12441_));
 sky130_fd_sc_hd__a21boi_4 _42984_ (.A1(_12113_),
    .A2(_12118_),
    .B1_N(_12116_),
    .Y(_12442_));
 sky130_fd_sc_hd__nand2_4 _42985_ (.A(_12441_),
    .B(_12442_),
    .Y(_12443_));
 sky130_vsdinv _42986_ (.A(_12442_),
    .Y(_12444_));
 sky130_fd_sc_hd__nand3_4 _42987_ (.A(_12438_),
    .B(_12444_),
    .C(_12440_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand2_4 _42988_ (.A(_12443_),
    .B(_12445_),
    .Y(_12446_));
 sky130_fd_sc_hd__nand2_4 _42989_ (.A(_12425_),
    .B(_12446_),
    .Y(_12447_));
 sky130_vsdinv _42990_ (.A(_12446_),
    .Y(_12448_));
 sky130_fd_sc_hd__nand3_4 _42991_ (.A(_12448_),
    .B(_12424_),
    .C(_12422_),
    .Y(_12449_));
 sky130_fd_sc_hd__nand2_4 _42992_ (.A(_12447_),
    .B(_12449_),
    .Y(_12450_));
 sky130_fd_sc_hd__a21boi_4 _42993_ (.A1(_12106_),
    .A2(_12130_),
    .B1_N(_12108_),
    .Y(_12451_));
 sky130_fd_sc_hd__nand2_4 _42994_ (.A(_12450_),
    .B(_12451_),
    .Y(_12452_));
 sky130_vsdinv _42995_ (.A(_12451_),
    .Y(_12453_));
 sky130_fd_sc_hd__nand3_4 _42996_ (.A(_12453_),
    .B(_12447_),
    .C(_12449_),
    .Y(_12454_));
 sky130_fd_sc_hd__nand2_4 _42997_ (.A(_12452_),
    .B(_12454_),
    .Y(_12455_));
 sky130_fd_sc_hd__buf_1 _42998_ (.A(_07979_),
    .X(_12456_));
 sky130_fd_sc_hd__nand2_4 _42999_ (.A(_11015_),
    .B(_12456_),
    .Y(_12457_));
 sky130_fd_sc_hd__buf_1 _43000_ (.A(_07620_),
    .X(_12458_));
 sky130_fd_sc_hd__nand2_4 _43001_ (.A(_12458_),
    .B(_12142_),
    .Y(_12459_));
 sky130_fd_sc_hd__nand2_4 _43002_ (.A(_11014_),
    .B(_07977_),
    .Y(_12460_));
 sky130_fd_sc_hd__xnor2_4 _43003_ (.A(_12459_),
    .B(_12460_),
    .Y(_12461_));
 sky130_fd_sc_hd__xor2_4 _43004_ (.A(_12457_),
    .B(_12461_),
    .X(_12462_));
 sky130_fd_sc_hd__nand2_4 _43005_ (.A(_07147_),
    .B(_11503_),
    .Y(_12463_));
 sky130_fd_sc_hd__nand2_4 _43006_ (.A(_07605_),
    .B(_11502_),
    .Y(_12464_));
 sky130_fd_sc_hd__nand2_4 _43007_ (.A(_12463_),
    .B(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__buf_1 _43008_ (.A(_03569_),
    .X(_12466_));
 sky130_fd_sc_hd__buf_1 _43009_ (.A(_10275_),
    .X(_12467_));
 sky130_fd_sc_hd__nand4_4 _43010_ (.A(_07151_),
    .B(_07153_),
    .C(_12466_),
    .D(_12467_),
    .Y(_12468_));
 sky130_fd_sc_hd__nand2_4 _43011_ (.A(_07858_),
    .B(_11175_),
    .Y(_12469_));
 sky130_vsdinv _43012_ (.A(_12469_),
    .Y(_12470_));
 sky130_fd_sc_hd__nand3_4 _43013_ (.A(_12465_),
    .B(_12468_),
    .C(_12470_),
    .Y(_12471_));
 sky130_fd_sc_hd__a21o_4 _43014_ (.A1(_12465_),
    .A2(_12468_),
    .B1(_12470_),
    .X(_12472_));
 sky130_fd_sc_hd__a21boi_4 _43015_ (.A1(_12155_),
    .A2(_12160_),
    .B1_N(_12158_),
    .Y(_12473_));
 sky130_vsdinv _43016_ (.A(_12473_),
    .Y(_12474_));
 sky130_fd_sc_hd__a21o_4 _43017_ (.A1(_12471_),
    .A2(_12472_),
    .B1(_12474_),
    .X(_12475_));
 sky130_fd_sc_hd__nand3_4 _43018_ (.A(_12474_),
    .B(_12472_),
    .C(_12471_),
    .Y(_12476_));
 sky130_fd_sc_hd__nand3_4 _43019_ (.A(_12462_),
    .B(_12475_),
    .C(_12476_),
    .Y(_12477_));
 sky130_fd_sc_hd__nand2_4 _43020_ (.A(_12475_),
    .B(_12476_),
    .Y(_12478_));
 sky130_vsdinv _43021_ (.A(_12457_),
    .Y(_12479_));
 sky130_fd_sc_hd__xor2_4 _43022_ (.A(_12479_),
    .B(_12461_),
    .X(_12480_));
 sky130_fd_sc_hd__nand2_4 _43023_ (.A(_12478_),
    .B(_12480_),
    .Y(_12481_));
 sky130_fd_sc_hd__a21boi_4 _43024_ (.A1(_12123_),
    .A2(_12127_),
    .B1_N(_12125_),
    .Y(_12482_));
 sky130_vsdinv _43025_ (.A(_12482_),
    .Y(_12483_));
 sky130_fd_sc_hd__a21o_4 _43026_ (.A1(_12477_),
    .A2(_12481_),
    .B1(_12483_),
    .X(_12484_));
 sky130_fd_sc_hd__nand3_4 _43027_ (.A(_12483_),
    .B(_12477_),
    .C(_12481_),
    .Y(_12485_));
 sky130_fd_sc_hd__nand2_4 _43028_ (.A(_12484_),
    .B(_12485_),
    .Y(_12486_));
 sky130_fd_sc_hd__o21a_4 _43029_ (.A1(_12168_),
    .A2(_12167_),
    .B1(_12163_),
    .X(_12487_));
 sky130_fd_sc_hd__nand2_4 _43030_ (.A(_12486_),
    .B(_12487_),
    .Y(_12488_));
 sky130_vsdinv _43031_ (.A(_12487_),
    .Y(_12489_));
 sky130_fd_sc_hd__nand3_4 _43032_ (.A(_12484_),
    .B(_12489_),
    .C(_12485_),
    .Y(_12490_));
 sky130_fd_sc_hd__nand2_4 _43033_ (.A(_12488_),
    .B(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__nand2_4 _43034_ (.A(_12455_),
    .B(_12491_),
    .Y(_12492_));
 sky130_vsdinv _43035_ (.A(_12491_),
    .Y(_12493_));
 sky130_fd_sc_hd__nand3_4 _43036_ (.A(_12493_),
    .B(_12452_),
    .C(_12454_),
    .Y(_12494_));
 sky130_fd_sc_hd__nand2_4 _43037_ (.A(_12492_),
    .B(_12494_),
    .Y(_12495_));
 sky130_fd_sc_hd__a21boi_4 _43038_ (.A1(_12136_),
    .A2(_12178_),
    .B1_N(_12138_),
    .Y(_12496_));
 sky130_fd_sc_hd__nand2_4 _43039_ (.A(_12495_),
    .B(_12496_),
    .Y(_12497_));
 sky130_vsdinv _43040_ (.A(_12496_),
    .Y(_12498_));
 sky130_fd_sc_hd__nand3_4 _43041_ (.A(_12498_),
    .B(_12492_),
    .C(_12494_),
    .Y(_12499_));
 sky130_fd_sc_hd__nand2_4 _43042_ (.A(_12497_),
    .B(_12499_),
    .Y(_12500_));
 sky130_fd_sc_hd__nand2_4 _43043_ (.A(_07878_),
    .B(_07922_),
    .Y(_12501_));
 sky130_fd_sc_hd__nand2_4 _43044_ (.A(_08308_),
    .B(_07713_),
    .Y(_12502_));
 sky130_fd_sc_hd__nand2_4 _43045_ (.A(_12501_),
    .B(_12502_),
    .Y(_12503_));
 sky130_fd_sc_hd__nand4_4 _43046_ (.A(_11019_),
    .B(_10621_),
    .C(_10990_),
    .D(_03541_),
    .Y(_12504_));
 sky130_fd_sc_hd__nand2_4 _43047_ (.A(_11030_),
    .B(_03530_),
    .Y(_12505_));
 sky130_vsdinv _43048_ (.A(_12505_),
    .Y(_12506_));
 sky130_fd_sc_hd__a21o_4 _43049_ (.A1(_12503_),
    .A2(_12504_),
    .B1(_12506_),
    .X(_12507_));
 sky130_fd_sc_hd__nand3_4 _43050_ (.A(_12503_),
    .B(_12504_),
    .C(_12506_),
    .Y(_12508_));
 sky130_fd_sc_hd__nand2_4 _43051_ (.A(_12507_),
    .B(_12508_),
    .Y(_12509_));
 sky130_fd_sc_hd__a21o_4 _43052_ (.A1(_12148_),
    .A2(_12147_),
    .B1(_12509_),
    .X(_12510_));
 sky130_fd_sc_hd__nand3_4 _43053_ (.A(_12509_),
    .B(_12148_),
    .C(_12147_),
    .Y(_12511_));
 sky130_fd_sc_hd__a21boi_4 _43054_ (.A1(_12194_),
    .A2(_12197_),
    .B1_N(_12195_),
    .Y(_12512_));
 sky130_vsdinv _43055_ (.A(_12512_),
    .Y(_12513_));
 sky130_fd_sc_hd__a21o_4 _43056_ (.A1(_12510_),
    .A2(_12511_),
    .B1(_12513_),
    .X(_12514_));
 sky130_fd_sc_hd__nand3_4 _43057_ (.A(_12510_),
    .B(_12513_),
    .C(_12511_),
    .Y(_12515_));
 sky130_fd_sc_hd__nand2_4 _43058_ (.A(_12514_),
    .B(_12515_),
    .Y(_12516_));
 sky130_fd_sc_hd__a21boi_4 _43059_ (.A1(_12204_),
    .A2(_12208_),
    .B1_N(_12206_),
    .Y(_12517_));
 sky130_fd_sc_hd__nand2_4 _43060_ (.A(_12516_),
    .B(_12517_),
    .Y(_12518_));
 sky130_vsdinv _43061_ (.A(_12517_),
    .Y(_12519_));
 sky130_fd_sc_hd__nand3_4 _43062_ (.A(_12514_),
    .B(_12519_),
    .C(_12515_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand2_4 _43063_ (.A(_12518_),
    .B(_12520_),
    .Y(_12521_));
 sky130_fd_sc_hd__maj3_4 _43064_ (.A(_12223_),
    .B(_12217_),
    .C(_12218_),
    .X(_12522_));
 sky130_fd_sc_hd__buf_1 _43065_ (.A(_07193_),
    .X(_12523_));
 sky130_fd_sc_hd__nand2_4 _43066_ (.A(_08755_),
    .B(_12523_),
    .Y(_12524_));
 sky130_fd_sc_hd__nand2_4 _43067_ (.A(_09831_),
    .B(_07059_),
    .Y(_12525_));
 sky130_fd_sc_hd__nand2_4 _43068_ (.A(_12524_),
    .B(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__buf_1 _43069_ (.A(_07356_),
    .X(_12527_));
 sky130_fd_sc_hd__buf_1 _43070_ (.A(_07353_),
    .X(_12528_));
 sky130_fd_sc_hd__nand4_4 _43071_ (.A(_03358_),
    .B(_12225_),
    .C(_12527_),
    .D(_12528_),
    .Y(_12529_));
 sky130_fd_sc_hd__buf_1 _43072_ (.A(_09212_),
    .X(_12530_));
 sky130_fd_sc_hd__nand2_4 _43073_ (.A(_12530_),
    .B(_06881_),
    .Y(_12531_));
 sky130_fd_sc_hd__a21bo_4 _43074_ (.A1(_12526_),
    .A2(_12529_),
    .B1_N(_12531_),
    .X(_12532_));
 sky130_fd_sc_hd__buf_1 _43075_ (.A(_10785_),
    .X(_12533_));
 sky130_fd_sc_hd__nand4_4 _43076_ (.A(_12533_),
    .B(_12526_),
    .C(_12529_),
    .D(_07747_),
    .Y(_12534_));
 sky130_fd_sc_hd__nand2_4 _43077_ (.A(_12532_),
    .B(_12534_),
    .Y(_12535_));
 sky130_fd_sc_hd__nor2_4 _43078_ (.A(_12522_),
    .B(_12535_),
    .Y(_12536_));
 sky130_fd_sc_hd__a21boi_4 _43079_ (.A1(_12534_),
    .A2(_12532_),
    .B1_N(_12522_),
    .Y(_12537_));
 sky130_fd_sc_hd__nand2_4 _43080_ (.A(_10822_),
    .B(_07205_),
    .Y(_12538_));
 sky130_vsdinv _43081_ (.A(_12538_),
    .Y(_12539_));
 sky130_fd_sc_hd__nand2_4 _43082_ (.A(_09846_),
    .B(_07668_),
    .Y(_12540_));
 sky130_fd_sc_hd__nand2_4 _43083_ (.A(_09847_),
    .B(_06891_),
    .Y(_12541_));
 sky130_fd_sc_hd__xnor2_4 _43084_ (.A(_12540_),
    .B(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__xor2_4 _43085_ (.A(_12539_),
    .B(_12542_),
    .X(_12543_));
 sky130_fd_sc_hd__o21a_4 _43086_ (.A1(_12536_),
    .A2(_12537_),
    .B1(_12543_),
    .X(_12544_));
 sky130_vsdinv _43087_ (.A(_12543_),
    .Y(_12545_));
 sky130_vsdinv _43088_ (.A(_12537_),
    .Y(_12546_));
 sky130_vsdinv _43089_ (.A(_12536_),
    .Y(_12547_));
 sky130_fd_sc_hd__nand3_4 _43090_ (.A(_12545_),
    .B(_12546_),
    .C(_12547_),
    .Y(_12548_));
 sky130_vsdinv _43091_ (.A(_12548_),
    .Y(_12549_));
 sky130_fd_sc_hd__nor2_4 _43092_ (.A(_12544_),
    .B(_12549_),
    .Y(_12550_));
 sky130_vsdinv _43093_ (.A(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__nand2_4 _43094_ (.A(_12521_),
    .B(_12551_),
    .Y(_12552_));
 sky130_fd_sc_hd__nand3_4 _43095_ (.A(_12550_),
    .B(_12518_),
    .C(_12520_),
    .Y(_12553_));
 sky130_fd_sc_hd__nand2_4 _43096_ (.A(_12552_),
    .B(_12553_),
    .Y(_12554_));
 sky130_fd_sc_hd__a21boi_4 _43097_ (.A1(_12174_),
    .A2(_12172_),
    .B1_N(_12170_),
    .Y(_12555_));
 sky130_fd_sc_hd__nand2_4 _43098_ (.A(_12554_),
    .B(_12555_),
    .Y(_12556_));
 sky130_vsdinv _43099_ (.A(_12555_),
    .Y(_12557_));
 sky130_fd_sc_hd__nand3_4 _43100_ (.A(_12552_),
    .B(_12557_),
    .C(_12553_),
    .Y(_12558_));
 sky130_fd_sc_hd__nand2_4 _43101_ (.A(_12556_),
    .B(_12558_),
    .Y(_12559_));
 sky130_fd_sc_hd__o21a_4 _43102_ (.A1(_12243_),
    .A2(_12215_),
    .B1(_12214_),
    .X(_12560_));
 sky130_fd_sc_hd__nand2_4 _43103_ (.A(_12559_),
    .B(_12560_),
    .Y(_12561_));
 sky130_vsdinv _43104_ (.A(_12560_),
    .Y(_12562_));
 sky130_fd_sc_hd__nand3_4 _43105_ (.A(_12556_),
    .B(_12562_),
    .C(_12558_),
    .Y(_12563_));
 sky130_fd_sc_hd__nand2_4 _43106_ (.A(_12561_),
    .B(_12563_),
    .Y(_12564_));
 sky130_fd_sc_hd__nand2_4 _43107_ (.A(_12500_),
    .B(_12564_),
    .Y(_12565_));
 sky130_fd_sc_hd__a21oi_4 _43108_ (.A1(_12556_),
    .A2(_12558_),
    .B1(_12562_),
    .Y(_12566_));
 sky130_vsdinv _43109_ (.A(_12563_),
    .Y(_12567_));
 sky130_fd_sc_hd__nor2_4 _43110_ (.A(_12566_),
    .B(_12567_),
    .Y(_12568_));
 sky130_fd_sc_hd__nand3_4 _43111_ (.A(_12568_),
    .B(_12497_),
    .C(_12499_),
    .Y(_12569_));
 sky130_fd_sc_hd__nand2_4 _43112_ (.A(_12565_),
    .B(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__a21boi_4 _43113_ (.A1(_12260_),
    .A2(_12185_),
    .B1_N(_12187_),
    .Y(_12571_));
 sky130_fd_sc_hd__nand2_4 _43114_ (.A(_12570_),
    .B(_12571_),
    .Y(_12572_));
 sky130_vsdinv _43115_ (.A(_12571_),
    .Y(_12573_));
 sky130_fd_sc_hd__nand3_4 _43116_ (.A(_12573_),
    .B(_12565_),
    .C(_12569_),
    .Y(_12574_));
 sky130_fd_sc_hd__nand2_4 _43117_ (.A(_12572_),
    .B(_12574_),
    .Y(_12575_));
 sky130_vsdinv _43118_ (.A(_12229_),
    .Y(_12576_));
 sky130_fd_sc_hd__o21a_4 _43119_ (.A1(_12230_),
    .A2(_12239_),
    .B1(_12576_),
    .X(_12577_));
 sky130_vsdinv _43120_ (.A(_12577_),
    .Y(_12578_));
 sky130_fd_sc_hd__nand2_4 _43121_ (.A(_10826_),
    .B(_03491_),
    .Y(_12579_));
 sky130_fd_sc_hd__nand2_4 _43122_ (.A(_03393_),
    .B(_06477_),
    .Y(_12580_));
 sky130_fd_sc_hd__nand2_4 _43123_ (.A(_12579_),
    .B(_12580_),
    .Y(_12581_));
 sky130_fd_sc_hd__nand4_4 _43124_ (.A(_12278_),
    .B(_10409_),
    .C(_07096_),
    .D(_08082_),
    .Y(_12582_));
 sky130_fd_sc_hd__nand2_4 _43125_ (.A(_12581_),
    .B(_12582_),
    .Y(_12583_));
 sky130_fd_sc_hd__nand2_4 _43126_ (.A(_11333_),
    .B(_06796_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand2_4 _43127_ (.A(_12583_),
    .B(_12584_),
    .Y(_12585_));
 sky130_vsdinv _43128_ (.A(_12584_),
    .Y(_12586_));
 sky130_fd_sc_hd__nand3_4 _43129_ (.A(_12581_),
    .B(_12582_),
    .C(_12586_),
    .Y(_12587_));
 sky130_fd_sc_hd__and2_4 _43130_ (.A(_12585_),
    .B(_12587_),
    .X(_12588_));
 sky130_vsdinv _43131_ (.A(_12588_),
    .Y(_12589_));
 sky130_fd_sc_hd__a21boi_4 _43132_ (.A1(_12232_),
    .A2(_12236_),
    .B1_N(_12234_),
    .Y(_12590_));
 sky130_fd_sc_hd__nand2_4 _43133_ (.A(_12589_),
    .B(_12590_),
    .Y(_12591_));
 sky130_fd_sc_hd__nand2_4 _43134_ (.A(_12238_),
    .B(_12234_),
    .Y(_12592_));
 sky130_fd_sc_hd__nand2_4 _43135_ (.A(_12592_),
    .B(_12588_),
    .Y(_12593_));
 sky130_fd_sc_hd__a21boi_4 _43136_ (.A1(_12276_),
    .A2(_12282_),
    .B1_N(_12280_),
    .Y(_12594_));
 sky130_vsdinv _43137_ (.A(_12594_),
    .Y(_12595_));
 sky130_fd_sc_hd__nand3_4 _43138_ (.A(_12591_),
    .B(_12593_),
    .C(_12595_),
    .Y(_12596_));
 sky130_fd_sc_hd__nand2_4 _43139_ (.A(_12591_),
    .B(_12593_),
    .Y(_12597_));
 sky130_fd_sc_hd__nand2_4 _43140_ (.A(_12597_),
    .B(_12594_),
    .Y(_12598_));
 sky130_fd_sc_hd__nand3_4 _43141_ (.A(_12578_),
    .B(_12596_),
    .C(_12598_),
    .Y(_12599_));
 sky130_fd_sc_hd__nand2_4 _43142_ (.A(_12598_),
    .B(_12596_),
    .Y(_12600_));
 sky130_fd_sc_hd__nand2_4 _43143_ (.A(_12600_),
    .B(_12577_),
    .Y(_12601_));
 sky130_fd_sc_hd__nand2_4 _43144_ (.A(_12599_),
    .B(_12601_),
    .Y(_12602_));
 sky130_fd_sc_hd__a21boi_4 _43145_ (.A1(_12287_),
    .A2(_12291_),
    .B1_N(_12289_),
    .Y(_12603_));
 sky130_fd_sc_hd__nand2_4 _43146_ (.A(_12602_),
    .B(_12603_),
    .Y(_12604_));
 sky130_vsdinv _43147_ (.A(_12603_),
    .Y(_12605_));
 sky130_fd_sc_hd__nand3_4 _43148_ (.A(_12599_),
    .B(_12601_),
    .C(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__a21boi_4 _43149_ (.A1(_12298_),
    .A2(_12296_),
    .B1_N(_12294_),
    .Y(_12607_));
 sky130_vsdinv _43150_ (.A(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__a21o_4 _43151_ (.A1(_12604_),
    .A2(_12606_),
    .B1(_12608_),
    .X(_12609_));
 sky130_fd_sc_hd__nand3_4 _43152_ (.A(_12608_),
    .B(_12604_),
    .C(_12606_),
    .Y(_12610_));
 sky130_fd_sc_hd__nand2_4 _43153_ (.A(_12609_),
    .B(_12610_),
    .Y(_12611_));
 sky130_fd_sc_hd__buf_1 _43154_ (.A(_12317_),
    .X(_12612_));
 sky130_fd_sc_hd__a21boi_4 _43155_ (.A1(_12312_),
    .A2(_12612_),
    .B1_N(_12314_),
    .Y(_12613_));
 sky130_fd_sc_hd__nand2_4 _43156_ (.A(_12313_),
    .B(_06229_),
    .Y(_12614_));
 sky130_fd_sc_hd__nand2_4 _43157_ (.A(_11687_),
    .B(_06228_),
    .Y(_12615_));
 sky130_fd_sc_hd__nand2_4 _43158_ (.A(_12614_),
    .B(_12615_),
    .Y(_12616_));
 sky130_fd_sc_hd__nand4_4 _43159_ (.A(_11337_),
    .B(_11692_),
    .C(_06427_),
    .D(_06696_),
    .Y(_12617_));
 sky130_fd_sc_hd__a21o_4 _43160_ (.A1(_12616_),
    .A2(_12617_),
    .B1(_12318_),
    .X(_12618_));
 sky130_fd_sc_hd__nand3_4 _43161_ (.A(_12616_),
    .B(_12617_),
    .C(_12612_),
    .Y(_12619_));
 sky130_fd_sc_hd__nand2_4 _43162_ (.A(_12618_),
    .B(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__nor2_4 _43163_ (.A(_12613_),
    .B(_12620_),
    .Y(_12621_));
 sky130_vsdinv _43164_ (.A(_12621_),
    .Y(_12622_));
 sky130_fd_sc_hd__nand2_4 _43165_ (.A(_12620_),
    .B(_12613_),
    .Y(_12623_));
 sky130_fd_sc_hd__a21o_4 _43166_ (.A1(_12622_),
    .A2(_12623_),
    .B1(_12006_),
    .X(_12624_));
 sky130_fd_sc_hd__nand3_4 _43167_ (.A(_12622_),
    .B(_12006_),
    .C(_12623_),
    .Y(_12625_));
 sky130_fd_sc_hd__a21oi_4 _43168_ (.A1(_12325_),
    .A2(_12324_),
    .B1(_12322_),
    .Y(_12626_));
 sky130_vsdinv _43169_ (.A(_12626_),
    .Y(_12627_));
 sky130_fd_sc_hd__a21o_4 _43170_ (.A1(_12624_),
    .A2(_12625_),
    .B1(_12627_),
    .X(_12628_));
 sky130_fd_sc_hd__nand3_4 _43171_ (.A(_12624_),
    .B(_12625_),
    .C(_12627_),
    .Y(_12629_));
 sky130_fd_sc_hd__a21o_4 _43172_ (.A1(_12628_),
    .A2(_12629_),
    .B1(_12337_),
    .X(_12630_));
 sky130_fd_sc_hd__nand3_4 _43173_ (.A(_12628_),
    .B(_12335_),
    .C(_12629_),
    .Y(_12631_));
 sky130_fd_sc_hd__and2_4 _43174_ (.A(_12630_),
    .B(_12631_),
    .X(_12632_));
 sky130_vsdinv _43175_ (.A(_12632_),
    .Y(_12633_));
 sky130_fd_sc_hd__nand2_4 _43176_ (.A(_12611_),
    .B(_12633_),
    .Y(_12634_));
 sky130_fd_sc_hd__nand3_4 _43177_ (.A(_12632_),
    .B(_12609_),
    .C(_12610_),
    .Y(_12635_));
 sky130_fd_sc_hd__nand2_4 _43178_ (.A(_12634_),
    .B(_12635_),
    .Y(_12636_));
 sky130_fd_sc_hd__a21boi_4 _43179_ (.A1(_12250_),
    .A2(_12253_),
    .B1_N(_12251_),
    .Y(_12637_));
 sky130_fd_sc_hd__nand2_4 _43180_ (.A(_12636_),
    .B(_12637_),
    .Y(_12638_));
 sky130_vsdinv _43181_ (.A(_12637_),
    .Y(_12639_));
 sky130_fd_sc_hd__nand3_4 _43182_ (.A(_12634_),
    .B(_12639_),
    .C(_12635_),
    .Y(_12640_));
 sky130_fd_sc_hd__buf_1 _43183_ (.A(_12640_),
    .X(_12641_));
 sky130_fd_sc_hd__a21boi_4 _43184_ (.A1(_12303_),
    .A2(_12340_),
    .B1_N(_12305_),
    .Y(_12642_));
 sky130_vsdinv _43185_ (.A(_12642_),
    .Y(_12643_));
 sky130_fd_sc_hd__a21o_4 _43186_ (.A1(_12638_),
    .A2(_12641_),
    .B1(_12643_),
    .X(_12644_));
 sky130_fd_sc_hd__nand3_4 _43187_ (.A(_12638_),
    .B(_12643_),
    .C(_12640_),
    .Y(_12645_));
 sky130_fd_sc_hd__nand2_4 _43188_ (.A(_12644_),
    .B(_12645_),
    .Y(_12646_));
 sky130_fd_sc_hd__nand2_4 _43189_ (.A(_12575_),
    .B(_12646_),
    .Y(_12647_));
 sky130_fd_sc_hd__a21oi_4 _43190_ (.A1(_12638_),
    .A2(_12641_),
    .B1(_12643_),
    .Y(_12648_));
 sky130_vsdinv _43191_ (.A(_12645_),
    .Y(_12649_));
 sky130_fd_sc_hd__nor2_4 _43192_ (.A(_12648_),
    .B(_12649_),
    .Y(_12650_));
 sky130_fd_sc_hd__nand3_4 _43193_ (.A(_12650_),
    .B(_12572_),
    .C(_12574_),
    .Y(_12651_));
 sky130_fd_sc_hd__nand2_4 _43194_ (.A(_12647_),
    .B(_12651_),
    .Y(_12652_));
 sky130_fd_sc_hd__a21boi_4 _43195_ (.A1(_12358_),
    .A2(_12264_),
    .B1_N(_12267_),
    .Y(_12653_));
 sky130_fd_sc_hd__nand2_4 _43196_ (.A(_12652_),
    .B(_12653_),
    .Y(_12654_));
 sky130_vsdinv _43197_ (.A(_12653_),
    .Y(_12655_));
 sky130_fd_sc_hd__nand3_4 _43198_ (.A(_12655_),
    .B(_12647_),
    .C(_12651_),
    .Y(_12656_));
 sky130_fd_sc_hd__nand2_4 _43199_ (.A(_12654_),
    .B(_12656_),
    .Y(_12657_));
 sky130_fd_sc_hd__buf_1 _43200_ (.A(_12335_),
    .X(_12658_));
 sky130_fd_sc_hd__a21boi_4 _43201_ (.A1(_12330_),
    .A2(_12658_),
    .B1_N(_12332_),
    .Y(_12659_));
 sky130_fd_sc_hd__a21boi_4 _43202_ (.A1(_12346_),
    .A2(_12351_),
    .B1_N(_12349_),
    .Y(_12660_));
 sky130_fd_sc_hd__xnor2_4 _43203_ (.A(_12659_),
    .B(_12660_),
    .Y(_12661_));
 sky130_fd_sc_hd__nand2_4 _43204_ (.A(_12657_),
    .B(_12661_),
    .Y(_12662_));
 sky130_vsdinv _43205_ (.A(_12661_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand3_4 _43206_ (.A(_12654_),
    .B(_12656_),
    .C(_12663_),
    .Y(_12664_));
 sky130_fd_sc_hd__nand2_4 _43207_ (.A(_12662_),
    .B(_12664_),
    .Y(_12665_));
 sky130_fd_sc_hd__a21boi_4 _43208_ (.A1(_12362_),
    .A2(_12371_),
    .B1_N(_12365_),
    .Y(_12666_));
 sky130_fd_sc_hd__nand2_4 _43209_ (.A(_12665_),
    .B(_12666_),
    .Y(_12667_));
 sky130_vsdinv _43210_ (.A(_12666_),
    .Y(_12668_));
 sky130_fd_sc_hd__nand3_4 _43211_ (.A(_12668_),
    .B(_12662_),
    .C(_12664_),
    .Y(_12669_));
 sky130_fd_sc_hd__nand2_4 _43212_ (.A(_12667_),
    .B(_12669_),
    .Y(_12670_));
 sky130_fd_sc_hd__a21oi_4 _43213_ (.A1(_12033_),
    .A2(_12028_),
    .B1(_12367_),
    .Y(_12671_));
 sky130_vsdinv _43214_ (.A(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__nand2_4 _43215_ (.A(_12670_),
    .B(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__nand3_4 _43216_ (.A(_12667_),
    .B(_12671_),
    .C(_12669_),
    .Y(_12674_));
 sky130_fd_sc_hd__nand2_4 _43217_ (.A(_12673_),
    .B(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__a21boi_4 _43218_ (.A1(_12375_),
    .A2(_12379_),
    .B1_N(_12377_),
    .Y(_12676_));
 sky130_fd_sc_hd__nand2_4 _43219_ (.A(_12675_),
    .B(_12676_),
    .Y(_12677_));
 sky130_vsdinv _43220_ (.A(_12676_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand3_4 _43221_ (.A(_12678_),
    .B(_12674_),
    .C(_12673_),
    .Y(_12679_));
 sky130_fd_sc_hd__nand2_4 _43222_ (.A(_12677_),
    .B(_12679_),
    .Y(_12680_));
 sky130_fd_sc_hd__nand4_4 _43223_ (.A(_12067_),
    .B(_12065_),
    .C(_12385_),
    .D(_12387_),
    .Y(_12681_));
 sky130_fd_sc_hd__nor3_4 _43224_ (.A(_11409_),
    .B(_11756_),
    .C(_12681_),
    .Y(_12682_));
 sky130_vsdinv _43225_ (.A(_12067_),
    .Y(_12683_));
 sky130_fd_sc_hd__a21boi_4 _43226_ (.A1(_12683_),
    .A2(_12385_),
    .B1_N(_12387_),
    .Y(_12684_));
 sky130_fd_sc_hd__o21ai_4 _43227_ (.A1(_12071_),
    .A2(_12681_),
    .B1(_12684_),
    .Y(_12685_));
 sky130_fd_sc_hd__a21oi_4 _43228_ (.A1(_11427_),
    .A2(_12682_),
    .B1(_12685_),
    .Y(_12686_));
 sky130_fd_sc_hd__xor2_4 _43229_ (.A(_12680_),
    .B(_12686_),
    .X(_01441_));
 sky130_fd_sc_hd__a21boi_4 _43230_ (.A1(_12392_),
    .A2(_12398_),
    .B1_N(_12394_),
    .Y(_12687_));
 sky130_vsdinv _43231_ (.A(_12687_),
    .Y(_12688_));
 sky130_fd_sc_hd__nand2_4 _43232_ (.A(_06084_),
    .B(_12390_),
    .Y(_12689_));
 sky130_fd_sc_hd__o21ai_4 _43233_ (.A1(_07938_),
    .A2(_11101_),
    .B1(_12689_),
    .Y(_12690_));
 sky130_fd_sc_hd__nand2_4 _43234_ (.A(_06544_),
    .B(_10515_),
    .Y(_12691_));
 sky130_vsdinv _43235_ (.A(_12691_),
    .Y(_12692_));
 sky130_fd_sc_hd__nand4_4 _43236_ (.A(_03269_),
    .B(_06325_),
    .C(_12390_),
    .D(_11106_),
    .Y(_12693_));
 sky130_fd_sc_hd__nand3_4 _43237_ (.A(_12690_),
    .B(_12692_),
    .C(_12693_),
    .Y(_12694_));
 sky130_fd_sc_hd__nand2_4 _43238_ (.A(_12690_),
    .B(_12693_),
    .Y(_12695_));
 sky130_fd_sc_hd__nand2_4 _43239_ (.A(_12695_),
    .B(_12691_),
    .Y(_12696_));
 sky130_fd_sc_hd__nand3_4 _43240_ (.A(_12688_),
    .B(_12694_),
    .C(_12696_),
    .Y(_12697_));
 sky130_fd_sc_hd__nand2_4 _43241_ (.A(_12696_),
    .B(_12694_),
    .Y(_12698_));
 sky130_fd_sc_hd__nand2_4 _43242_ (.A(_12698_),
    .B(_12687_),
    .Y(_12699_));
 sky130_fd_sc_hd__nand2_4 _43243_ (.A(_12697_),
    .B(_12699_),
    .Y(_12700_));
 sky130_fd_sc_hd__nand2_4 _43244_ (.A(_06255_),
    .B(_10947_),
    .Y(_12701_));
 sky130_fd_sc_hd__nand2_4 _43245_ (.A(_06446_),
    .B(_10946_),
    .Y(_12702_));
 sky130_fd_sc_hd__nand2_4 _43246_ (.A(_12701_),
    .B(_12702_),
    .Y(_12703_));
 sky130_fd_sc_hd__nand4_4 _43247_ (.A(_06255_),
    .B(_06446_),
    .C(_10946_),
    .D(_10947_),
    .Y(_12704_));
 sky130_fd_sc_hd__nand2_4 _43248_ (.A(_03294_),
    .B(_10508_),
    .Y(_12705_));
 sky130_vsdinv _43249_ (.A(_12705_),
    .Y(_12706_));
 sky130_fd_sc_hd__a21o_4 _43250_ (.A1(_12703_),
    .A2(_12704_),
    .B1(_12706_),
    .X(_12707_));
 sky130_fd_sc_hd__nand3_4 _43251_ (.A(_12703_),
    .B(_12704_),
    .C(_12706_),
    .Y(_12708_));
 sky130_fd_sc_hd__nand2_4 _43252_ (.A(_12707_),
    .B(_12708_),
    .Y(_12709_));
 sky130_fd_sc_hd__nand2_4 _43253_ (.A(_12700_),
    .B(_12709_),
    .Y(_12710_));
 sky130_fd_sc_hd__nand4_4 _43254_ (.A(_12708_),
    .B(_12697_),
    .C(_12699_),
    .D(_12707_),
    .Y(_12711_));
 sky130_fd_sc_hd__nand2_4 _43255_ (.A(_12710_),
    .B(_12711_),
    .Y(_12712_));
 sky130_vsdinv _43256_ (.A(_12402_),
    .Y(_12713_));
 sky130_fd_sc_hd__a21oi_4 _43257_ (.A1(_12401_),
    .A2(_12418_),
    .B1(_12713_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand2_4 _43258_ (.A(_12712_),
    .B(_12714_),
    .Y(_12715_));
 sky130_fd_sc_hd__a21o_4 _43259_ (.A1(_12401_),
    .A2(_12418_),
    .B1(_12713_),
    .X(_12716_));
 sky130_fd_sc_hd__nand3_4 _43260_ (.A(_12716_),
    .B(_12711_),
    .C(_12710_),
    .Y(_12717_));
 sky130_fd_sc_hd__nand2_4 _43261_ (.A(_12715_),
    .B(_12717_),
    .Y(_12718_));
 sky130_fd_sc_hd__buf_1 _43262_ (.A(_10300_),
    .X(_12719_));
 sky130_fd_sc_hd__nand2_4 _43263_ (.A(_06983_),
    .B(_12719_),
    .Y(_12720_));
 sky130_fd_sc_hd__buf_1 _43264_ (.A(_10481_),
    .X(_12721_));
 sky130_fd_sc_hd__nand2_4 _43265_ (.A(_06996_),
    .B(_12721_),
    .Y(_12722_));
 sky130_fd_sc_hd__nand2_4 _43266_ (.A(_12720_),
    .B(_12722_),
    .Y(_12723_));
 sky130_fd_sc_hd__nand4_4 _43267_ (.A(_06983_),
    .B(_06996_),
    .C(_03588_),
    .D(_12719_),
    .Y(_12724_));
 sky130_fd_sc_hd__nand2_4 _43268_ (.A(_07151_),
    .B(_03582_),
    .Y(_12725_));
 sky130_vsdinv _43269_ (.A(_12725_),
    .Y(_12726_));
 sky130_fd_sc_hd__nand3_4 _43270_ (.A(_12723_),
    .B(_12724_),
    .C(_12726_),
    .Y(_12727_));
 sky130_fd_sc_hd__a21o_4 _43271_ (.A1(_12723_),
    .A2(_12724_),
    .B1(_12726_),
    .X(_12728_));
 sky130_fd_sc_hd__a21boi_4 _43272_ (.A1(_12408_),
    .A2(_12413_),
    .B1_N(_12411_),
    .Y(_12729_));
 sky130_vsdinv _43273_ (.A(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__a21o_4 _43274_ (.A1(_12727_),
    .A2(_12728_),
    .B1(_12730_),
    .X(_12731_));
 sky130_fd_sc_hd__nand3_4 _43275_ (.A(_12730_),
    .B(_12728_),
    .C(_12727_),
    .Y(_12732_));
 sky130_fd_sc_hd__a21boi_4 _43276_ (.A1(_12429_),
    .A2(_12434_),
    .B1_N(_12432_),
    .Y(_12733_));
 sky130_vsdinv _43277_ (.A(_12733_),
    .Y(_12734_));
 sky130_fd_sc_hd__a21o_4 _43278_ (.A1(_12731_),
    .A2(_12732_),
    .B1(_12734_),
    .X(_12735_));
 sky130_fd_sc_hd__nand3_4 _43279_ (.A(_12731_),
    .B(_12732_),
    .C(_12734_),
    .Y(_12736_));
 sky130_fd_sc_hd__nand2_4 _43280_ (.A(_12735_),
    .B(_12736_),
    .Y(_12737_));
 sky130_fd_sc_hd__nand2_4 _43281_ (.A(_12718_),
    .B(_12737_),
    .Y(_12738_));
 sky130_fd_sc_hd__nand4_4 _43282_ (.A(_12736_),
    .B(_12715_),
    .C(_12735_),
    .D(_12717_),
    .Y(_12739_));
 sky130_fd_sc_hd__nand2_4 _43283_ (.A(_12738_),
    .B(_12739_),
    .Y(_12740_));
 sky130_fd_sc_hd__a21boi_4 _43284_ (.A1(_12417_),
    .A2(_12419_),
    .B1_N(_12421_),
    .Y(_12741_));
 sky130_fd_sc_hd__o21ai_4 _43285_ (.A1(_12446_),
    .A2(_12741_),
    .B1(_12424_),
    .Y(_12742_));
 sky130_vsdinv _43286_ (.A(_12742_),
    .Y(_12743_));
 sky130_fd_sc_hd__nand2_4 _43287_ (.A(_12740_),
    .B(_12743_),
    .Y(_12744_));
 sky130_fd_sc_hd__nand3_4 _43288_ (.A(_12742_),
    .B(_12738_),
    .C(_12739_),
    .Y(_12745_));
 sky130_fd_sc_hd__nand2_4 _43289_ (.A(_12744_),
    .B(_12745_),
    .Y(_12746_));
 sky130_fd_sc_hd__a21boi_4 _43290_ (.A1(_12465_),
    .A2(_12470_),
    .B1_N(_12468_),
    .Y(_12747_));
 sky130_fd_sc_hd__nand2_4 _43291_ (.A(_06992_),
    .B(_10537_),
    .Y(_12748_));
 sky130_fd_sc_hd__nand2_4 _43292_ (.A(_08026_),
    .B(_10536_),
    .Y(_12749_));
 sky130_fd_sc_hd__nand2_4 _43293_ (.A(_12748_),
    .B(_12749_),
    .Y(_12750_));
 sky130_fd_sc_hd__nand4_4 _43294_ (.A(_07422_),
    .B(_03318_),
    .C(_10884_),
    .D(_10885_),
    .Y(_12751_));
 sky130_fd_sc_hd__nand2_4 _43295_ (.A(_07621_),
    .B(_11175_),
    .Y(_12752_));
 sky130_fd_sc_hd__a21bo_4 _43296_ (.A1(_12750_),
    .A2(_12751_),
    .B1_N(_12752_),
    .X(_12753_));
 sky130_fd_sc_hd__buf_1 _43297_ (.A(_08635_),
    .X(_12754_));
 sky130_fd_sc_hd__nand4_4 _43298_ (.A(_07295_),
    .B(_12750_),
    .C(_12751_),
    .D(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__nand2_4 _43299_ (.A(_12753_),
    .B(_12755_),
    .Y(_12756_));
 sky130_fd_sc_hd__nor2_4 _43300_ (.A(_12747_),
    .B(_12756_),
    .Y(_12757_));
 sky130_vsdinv _43301_ (.A(_12757_),
    .Y(_12758_));
 sky130_fd_sc_hd__nand2_4 _43302_ (.A(_12756_),
    .B(_12747_),
    .Y(_12759_));
 sky130_fd_sc_hd__nand2_4 _43303_ (.A(_10212_),
    .B(_09416_),
    .Y(_12760_));
 sky130_fd_sc_hd__o21ai_4 _43304_ (.A1(_03333_),
    .A2(_03558_),
    .B1(_12760_),
    .Y(_12761_));
 sky130_fd_sc_hd__buf_1 _43305_ (.A(_08643_),
    .X(_12762_));
 sky130_fd_sc_hd__nand4_4 _43306_ (.A(_11557_),
    .B(_11559_),
    .C(_12762_),
    .D(_08198_),
    .Y(_12763_));
 sky130_fd_sc_hd__nand2_4 _43307_ (.A(_11019_),
    .B(_12144_),
    .Y(_12764_));
 sky130_vsdinv _43308_ (.A(_12764_),
    .Y(_12765_));
 sky130_fd_sc_hd__a21o_4 _43309_ (.A1(_12761_),
    .A2(_12763_),
    .B1(_12765_),
    .X(_12766_));
 sky130_fd_sc_hd__nand3_4 _43310_ (.A(_12761_),
    .B(_12763_),
    .C(_12765_),
    .Y(_12767_));
 sky130_fd_sc_hd__and2_4 _43311_ (.A(_12766_),
    .B(_12767_),
    .X(_12768_));
 sky130_fd_sc_hd__buf_1 _43312_ (.A(_12768_),
    .X(_12769_));
 sky130_fd_sc_hd__a21o_4 _43313_ (.A1(_12758_),
    .A2(_12759_),
    .B1(_12769_),
    .X(_12770_));
 sky130_fd_sc_hd__nand3_4 _43314_ (.A(_12758_),
    .B(_12769_),
    .C(_12759_),
    .Y(_12771_));
 sky130_fd_sc_hd__nand2_4 _43315_ (.A(_12770_),
    .B(_12771_),
    .Y(_12772_));
 sky130_fd_sc_hd__maj3_4 _43316_ (.A(_12442_),
    .B(_12437_),
    .C(_12439_),
    .X(_12773_));
 sky130_fd_sc_hd__nand2_4 _43317_ (.A(_12772_),
    .B(_12773_),
    .Y(_12774_));
 sky130_vsdinv _43318_ (.A(_12773_),
    .Y(_12775_));
 sky130_fd_sc_hd__nand3_4 _43319_ (.A(_12770_),
    .B(_12775_),
    .C(_12771_),
    .Y(_12776_));
 sky130_fd_sc_hd__a21boi_4 _43320_ (.A1(_12462_),
    .A2(_12475_),
    .B1_N(_12476_),
    .Y(_12777_));
 sky130_vsdinv _43321_ (.A(_12777_),
    .Y(_12778_));
 sky130_fd_sc_hd__a21oi_4 _43322_ (.A1(_12774_),
    .A2(_12776_),
    .B1(_12778_),
    .Y(_12779_));
 sky130_vsdinv _43323_ (.A(_12779_),
    .Y(_12780_));
 sky130_fd_sc_hd__nand3_4 _43324_ (.A(_12774_),
    .B(_12778_),
    .C(_12776_),
    .Y(_12781_));
 sky130_fd_sc_hd__nand2_4 _43325_ (.A(_12780_),
    .B(_12781_),
    .Y(_12782_));
 sky130_fd_sc_hd__nand2_4 _43326_ (.A(_12746_),
    .B(_12782_),
    .Y(_12783_));
 sky130_fd_sc_hd__nand4_4 _43327_ (.A(_12781_),
    .B(_12744_),
    .C(_12780_),
    .D(_12745_),
    .Y(_12784_));
 sky130_fd_sc_hd__nand2_4 _43328_ (.A(_12783_),
    .B(_12784_),
    .Y(_12785_));
 sky130_fd_sc_hd__a21boi_4 _43329_ (.A1(_12493_),
    .A2(_12452_),
    .B1_N(_12454_),
    .Y(_12786_));
 sky130_fd_sc_hd__nand2_4 _43330_ (.A(_12785_),
    .B(_12786_),
    .Y(_12787_));
 sky130_fd_sc_hd__a21boi_4 _43331_ (.A1(_12447_),
    .A2(_12449_),
    .B1_N(_12451_),
    .Y(_12788_));
 sky130_fd_sc_hd__o21ai_4 _43332_ (.A1(_12491_),
    .A2(_12788_),
    .B1(_12454_),
    .Y(_12789_));
 sky130_fd_sc_hd__nand3_4 _43333_ (.A(_12789_),
    .B(_12783_),
    .C(_12784_),
    .Y(_12790_));
 sky130_fd_sc_hd__nand2_4 _43334_ (.A(_12787_),
    .B(_12790_),
    .Y(_12791_));
 sky130_fd_sc_hd__nand2_4 _43335_ (.A(_12515_),
    .B(_12510_),
    .Y(_12792_));
 sky130_vsdinv _43336_ (.A(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__maj3_4 _43337_ (.A(_12457_),
    .B(_12459_),
    .C(_12460_),
    .X(_12794_));
 sky130_fd_sc_hd__nand2_4 _43338_ (.A(_10621_),
    .B(_08125_),
    .Y(_12795_));
 sky130_fd_sc_hd__nand2_4 _43339_ (.A(_08748_),
    .B(_08572_),
    .Y(_12796_));
 sky130_fd_sc_hd__nand2_4 _43340_ (.A(_12795_),
    .B(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__nand4_4 _43341_ (.A(_10625_),
    .B(_08753_),
    .C(_08357_),
    .D(_08358_),
    .Y(_12798_));
 sky130_fd_sc_hd__nand2_4 _43342_ (.A(_10664_),
    .B(_03530_),
    .Y(_12799_));
 sky130_vsdinv _43343_ (.A(_12799_),
    .Y(_12800_));
 sky130_fd_sc_hd__a21o_4 _43344_ (.A1(_12797_),
    .A2(_12798_),
    .B1(_12800_),
    .X(_12801_));
 sky130_fd_sc_hd__nand3_4 _43345_ (.A(_12797_),
    .B(_12798_),
    .C(_12800_),
    .Y(_12802_));
 sky130_fd_sc_hd__nand2_4 _43346_ (.A(_12801_),
    .B(_12802_),
    .Y(_12803_));
 sky130_fd_sc_hd__or2_4 _43347_ (.A(_12794_),
    .B(_12803_),
    .X(_12804_));
 sky130_fd_sc_hd__nand2_4 _43348_ (.A(_12803_),
    .B(_12794_),
    .Y(_12805_));
 sky130_fd_sc_hd__nand2_4 _43349_ (.A(_12804_),
    .B(_12805_),
    .Y(_12806_));
 sky130_fd_sc_hd__a21boi_4 _43350_ (.A1(_12503_),
    .A2(_12506_),
    .B1_N(_12504_),
    .Y(_12807_));
 sky130_fd_sc_hd__nand2_4 _43351_ (.A(_12806_),
    .B(_12807_),
    .Y(_12808_));
 sky130_vsdinv _43352_ (.A(_12807_),
    .Y(_12809_));
 sky130_fd_sc_hd__nand3_4 _43353_ (.A(_12804_),
    .B(_12809_),
    .C(_12805_),
    .Y(_12810_));
 sky130_fd_sc_hd__nand2_4 _43354_ (.A(_12808_),
    .B(_12810_),
    .Y(_12811_));
 sky130_fd_sc_hd__nand2_4 _43355_ (.A(_12793_),
    .B(_12811_),
    .Y(_12812_));
 sky130_fd_sc_hd__nand3_4 _43356_ (.A(_12792_),
    .B(_12810_),
    .C(_12808_),
    .Y(_12813_));
 sky130_fd_sc_hd__nand2_4 _43357_ (.A(_12812_),
    .B(_12813_),
    .Y(_12814_));
 sky130_fd_sc_hd__maj3_4 _43358_ (.A(_12531_),
    .B(_12524_),
    .C(_12525_),
    .X(_12815_));
 sky130_fd_sc_hd__nand2_4 _43359_ (.A(_12225_),
    .B(_07194_),
    .Y(_12816_));
 sky130_fd_sc_hd__buf_1 _43360_ (.A(_03365_),
    .X(_12817_));
 sky130_fd_sc_hd__nand2_4 _43361_ (.A(_12817_),
    .B(_07192_),
    .Y(_12818_));
 sky130_fd_sc_hd__nand2_4 _43362_ (.A(_12816_),
    .B(_12818_),
    .Y(_12819_));
 sky130_fd_sc_hd__nand4_4 _43363_ (.A(_08760_),
    .B(_09577_),
    .C(_03518_),
    .D(_12221_),
    .Y(_12820_));
 sky130_fd_sc_hd__buf_1 _43364_ (.A(_10703_),
    .X(_12821_));
 sky130_fd_sc_hd__nand2_4 _43365_ (.A(_12821_),
    .B(_03513_),
    .Y(_12822_));
 sky130_fd_sc_hd__a21bo_4 _43366_ (.A1(_12819_),
    .A2(_12820_),
    .B1_N(_12822_),
    .X(_12823_));
 sky130_fd_sc_hd__buf_1 _43367_ (.A(_10791_),
    .X(_12824_));
 sky130_fd_sc_hd__nand4_4 _43368_ (.A(_12824_),
    .B(_12819_),
    .C(_12820_),
    .D(_11023_),
    .Y(_12825_));
 sky130_fd_sc_hd__nand2_4 _43369_ (.A(_12823_),
    .B(_12825_),
    .Y(_12826_));
 sky130_fd_sc_hd__nor2_4 _43370_ (.A(_12815_),
    .B(_12826_),
    .Y(_12827_));
 sky130_fd_sc_hd__a21boi_4 _43371_ (.A1(_12825_),
    .A2(_12823_),
    .B1_N(_12815_),
    .Y(_12828_));
 sky130_fd_sc_hd__nand2_4 _43372_ (.A(_11957_),
    .B(_11590_),
    .Y(_12829_));
 sky130_fd_sc_hd__buf_1 _43373_ (.A(_10393_),
    .X(_12830_));
 sky130_fd_sc_hd__nand2_4 _43374_ (.A(_12830_),
    .B(_07215_),
    .Y(_12831_));
 sky130_fd_sc_hd__buf_1 _43375_ (.A(_09849_),
    .X(_12832_));
 sky130_fd_sc_hd__nand2_4 _43376_ (.A(_12832_),
    .B(_07213_),
    .Y(_12833_));
 sky130_fd_sc_hd__nand2_4 _43377_ (.A(_12831_),
    .B(_12833_),
    .Y(_12834_));
 sky130_fd_sc_hd__nand4_4 _43378_ (.A(_11954_),
    .B(_12273_),
    .C(_06888_),
    .D(_06894_),
    .Y(_12835_));
 sky130_fd_sc_hd__nand2_4 _43379_ (.A(_12834_),
    .B(_12835_),
    .Y(_12836_));
 sky130_fd_sc_hd__xor2_4 _43380_ (.A(_12829_),
    .B(_12836_),
    .X(_12837_));
 sky130_vsdinv _43381_ (.A(_12837_),
    .Y(_12838_));
 sky130_fd_sc_hd__o21a_4 _43382_ (.A1(_12827_),
    .A2(_12828_),
    .B1(_12838_),
    .X(_12839_));
 sky130_fd_sc_hd__nor2_4 _43383_ (.A(_12827_),
    .B(_12828_),
    .Y(_12840_));
 sky130_fd_sc_hd__nand2_4 _43384_ (.A(_12840_),
    .B(_12837_),
    .Y(_12841_));
 sky130_vsdinv _43385_ (.A(_12841_),
    .Y(_12842_));
 sky130_fd_sc_hd__nor2_4 _43386_ (.A(_12839_),
    .B(_12842_),
    .Y(_12843_));
 sky130_vsdinv _43387_ (.A(_12843_),
    .Y(_12844_));
 sky130_fd_sc_hd__nand2_4 _43388_ (.A(_12814_),
    .B(_12844_),
    .Y(_12845_));
 sky130_fd_sc_hd__nand3_4 _43389_ (.A(_12812_),
    .B(_12843_),
    .C(_12813_),
    .Y(_12846_));
 sky130_fd_sc_hd__nand2_4 _43390_ (.A(_12845_),
    .B(_12846_),
    .Y(_12847_));
 sky130_fd_sc_hd__a21boi_4 _43391_ (.A1(_12484_),
    .A2(_12489_),
    .B1_N(_12485_),
    .Y(_12848_));
 sky130_fd_sc_hd__nand2_4 _43392_ (.A(_12847_),
    .B(_12848_),
    .Y(_12849_));
 sky130_vsdinv _43393_ (.A(_12848_),
    .Y(_12850_));
 sky130_fd_sc_hd__nand3_4 _43394_ (.A(_12850_),
    .B(_12845_),
    .C(_12846_),
    .Y(_12851_));
 sky130_fd_sc_hd__a21boi_4 _43395_ (.A1(_12550_),
    .A2(_12518_),
    .B1_N(_12520_),
    .Y(_12852_));
 sky130_vsdinv _43396_ (.A(_12852_),
    .Y(_12853_));
 sky130_fd_sc_hd__a21oi_4 _43397_ (.A1(_12849_),
    .A2(_12851_),
    .B1(_12853_),
    .Y(_12854_));
 sky130_vsdinv _43398_ (.A(_12854_),
    .Y(_12855_));
 sky130_fd_sc_hd__nand3_4 _43399_ (.A(_12849_),
    .B(_12851_),
    .C(_12853_),
    .Y(_12856_));
 sky130_fd_sc_hd__nand2_4 _43400_ (.A(_12855_),
    .B(_12856_),
    .Y(_12857_));
 sky130_fd_sc_hd__nand2_4 _43401_ (.A(_12791_),
    .B(_12857_),
    .Y(_12858_));
 sky130_vsdinv _43402_ (.A(_12856_),
    .Y(_12859_));
 sky130_fd_sc_hd__nor2_4 _43403_ (.A(_12854_),
    .B(_12859_),
    .Y(_12860_));
 sky130_fd_sc_hd__nand3_4 _43404_ (.A(_12860_),
    .B(_12790_),
    .C(_12787_),
    .Y(_12861_));
 sky130_fd_sc_hd__nand2_4 _43405_ (.A(_12858_),
    .B(_12861_),
    .Y(_12862_));
 sky130_fd_sc_hd__a21boi_4 _43406_ (.A1(_12568_),
    .A2(_12497_),
    .B1_N(_12499_),
    .Y(_12863_));
 sky130_fd_sc_hd__nand2_4 _43407_ (.A(_12862_),
    .B(_12863_),
    .Y(_12864_));
 sky130_fd_sc_hd__a21boi_4 _43408_ (.A1(_12492_),
    .A2(_12494_),
    .B1_N(_12496_),
    .Y(_12865_));
 sky130_fd_sc_hd__o21ai_4 _43409_ (.A1(_12564_),
    .A2(_12865_),
    .B1(_12499_),
    .Y(_12866_));
 sky130_fd_sc_hd__nand3_4 _43410_ (.A(_12866_),
    .B(_12861_),
    .C(_12858_),
    .Y(_12867_));
 sky130_fd_sc_hd__nand2_4 _43411_ (.A(_12864_),
    .B(_12867_),
    .Y(_12868_));
 sky130_fd_sc_hd__a21oi_4 _43412_ (.A1(_12552_),
    .A2(_12553_),
    .B1(_12557_),
    .Y(_12869_));
 sky130_fd_sc_hd__o21ai_4 _43413_ (.A1(_12560_),
    .A2(_12869_),
    .B1(_12558_),
    .Y(_12870_));
 sky130_vsdinv _43414_ (.A(_12870_),
    .Y(_12871_));
 sky130_fd_sc_hd__o21ai_4 _43415_ (.A1(_12537_),
    .A2(_12543_),
    .B1(_12547_),
    .Y(_12872_));
 sky130_vsdinv _43416_ (.A(_12872_),
    .Y(_12873_));
 sky130_fd_sc_hd__maj3_4 _43417_ (.A(_12538_),
    .B(_12540_),
    .C(_12541_),
    .X(_12874_));
 sky130_fd_sc_hd__nand2_4 _43418_ (.A(_10409_),
    .B(_06788_),
    .Y(_12875_));
 sky130_fd_sc_hd__nand2_4 _43419_ (.A(_10845_),
    .B(_06946_),
    .Y(_12876_));
 sky130_fd_sc_hd__nand2_4 _43420_ (.A(_12875_),
    .B(_12876_),
    .Y(_12877_));
 sky130_fd_sc_hd__buf_1 _43421_ (.A(_10408_),
    .X(_12878_));
 sky130_fd_sc_hd__nand4_4 _43422_ (.A(_12878_),
    .B(_03396_),
    .C(_06376_),
    .D(_08082_),
    .Y(_12879_));
 sky130_fd_sc_hd__nand2_4 _43423_ (.A(_10836_),
    .B(_03476_),
    .Y(_12880_));
 sky130_vsdinv _43424_ (.A(_12880_),
    .Y(_12881_));
 sky130_fd_sc_hd__a21o_4 _43425_ (.A1(_12877_),
    .A2(_12879_),
    .B1(_12881_),
    .X(_12882_));
 sky130_fd_sc_hd__nand3_4 _43426_ (.A(_12877_),
    .B(_12879_),
    .C(_12881_),
    .Y(_12883_));
 sky130_fd_sc_hd__nand2_4 _43427_ (.A(_12882_),
    .B(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__nor2_4 _43428_ (.A(_12874_),
    .B(_12884_),
    .Y(_12885_));
 sky130_vsdinv _43429_ (.A(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__nand2_4 _43430_ (.A(_12884_),
    .B(_12874_),
    .Y(_12887_));
 sky130_fd_sc_hd__nand2_4 _43431_ (.A(_12886_),
    .B(_12887_),
    .Y(_12888_));
 sky130_fd_sc_hd__a21boi_4 _43432_ (.A1(_12581_),
    .A2(_12586_),
    .B1_N(_12582_),
    .Y(_12889_));
 sky130_fd_sc_hd__nand2_4 _43433_ (.A(_12888_),
    .B(_12889_),
    .Y(_12890_));
 sky130_vsdinv _43434_ (.A(_12889_),
    .Y(_12891_));
 sky130_fd_sc_hd__nand3_4 _43435_ (.A(_12886_),
    .B(_12891_),
    .C(_12887_),
    .Y(_12892_));
 sky130_fd_sc_hd__nand2_4 _43436_ (.A(_12890_),
    .B(_12892_),
    .Y(_12893_));
 sky130_fd_sc_hd__nand2_4 _43437_ (.A(_12873_),
    .B(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__nand3_4 _43438_ (.A(_12872_),
    .B(_12892_),
    .C(_12890_),
    .Y(_12895_));
 sky130_fd_sc_hd__nand2_4 _43439_ (.A(_12894_),
    .B(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__a21boi_4 _43440_ (.A1(_12591_),
    .A2(_12595_),
    .B1_N(_12593_),
    .Y(_12897_));
 sky130_fd_sc_hd__nand2_4 _43441_ (.A(_12896_),
    .B(_12897_),
    .Y(_12898_));
 sky130_vsdinv _43442_ (.A(_12897_),
    .Y(_12899_));
 sky130_fd_sc_hd__nand3_4 _43443_ (.A(_12894_),
    .B(_12899_),
    .C(_12895_),
    .Y(_12900_));
 sky130_fd_sc_hd__nand2_4 _43444_ (.A(_12898_),
    .B(_12900_),
    .Y(_12901_));
 sky130_fd_sc_hd__a21boi_4 _43445_ (.A1(_12605_),
    .A2(_12601_),
    .B1_N(_12599_),
    .Y(_12902_));
 sky130_fd_sc_hd__nand2_4 _43446_ (.A(_12901_),
    .B(_12902_),
    .Y(_12903_));
 sky130_fd_sc_hd__nand2_4 _43447_ (.A(_12606_),
    .B(_12599_),
    .Y(_12904_));
 sky130_fd_sc_hd__nand3_4 _43448_ (.A(_12904_),
    .B(_12900_),
    .C(_12898_),
    .Y(_12905_));
 sky130_fd_sc_hd__nand2_4 _43449_ (.A(_12903_),
    .B(_12905_),
    .Y(_12906_));
 sky130_fd_sc_hd__buf_1 _43450_ (.A(_11687_),
    .X(_12907_));
 sky130_fd_sc_hd__o21a_4 _43451_ (.A1(_03466_),
    .A2(_03473_),
    .B1(_12907_),
    .X(_12908_));
 sky130_fd_sc_hd__buf_1 _43452_ (.A(_11686_),
    .X(_12909_));
 sky130_fd_sc_hd__buf_1 _43453_ (.A(_12909_),
    .X(_12910_));
 sky130_fd_sc_hd__nand3_4 _43454_ (.A(_12910_),
    .B(_03466_),
    .C(_03473_),
    .Y(_12911_));
 sky130_fd_sc_hd__a21o_4 _43455_ (.A1(_12908_),
    .A2(_12911_),
    .B1(_12316_),
    .X(_12912_));
 sky130_fd_sc_hd__nand3_4 _43456_ (.A(_12908_),
    .B(_12316_),
    .C(_12911_),
    .Y(_12913_));
 sky130_fd_sc_hd__a21boi_4 _43457_ (.A1(_12616_),
    .A2(_12318_),
    .B1_N(_12617_),
    .Y(_12914_));
 sky130_vsdinv _43458_ (.A(_12914_),
    .Y(_12915_));
 sky130_fd_sc_hd__a21o_4 _43459_ (.A1(_12912_),
    .A2(_12913_),
    .B1(_12915_),
    .X(_12916_));
 sky130_fd_sc_hd__nand3_4 _43460_ (.A(_12915_),
    .B(_12912_),
    .C(_12913_),
    .Y(_12917_));
 sky130_vsdinv _43461_ (.A(_12004_),
    .Y(_12918_));
 sky130_fd_sc_hd__a21o_4 _43462_ (.A1(_12916_),
    .A2(_12917_),
    .B1(_12918_),
    .X(_12919_));
 sky130_fd_sc_hd__buf_1 _43463_ (.A(_12918_),
    .X(_12920_));
 sky130_fd_sc_hd__nand3_4 _43464_ (.A(_12920_),
    .B(_12916_),
    .C(_12917_),
    .Y(_12921_));
 sky130_fd_sc_hd__a21oi_4 _43465_ (.A1(_12005_),
    .A2(_12623_),
    .B1(_12621_),
    .Y(_12922_));
 sky130_vsdinv _43466_ (.A(_12922_),
    .Y(_12923_));
 sky130_fd_sc_hd__a21o_4 _43467_ (.A1(_12919_),
    .A2(_12921_),
    .B1(_12923_),
    .X(_12924_));
 sky130_fd_sc_hd__nand3_4 _43468_ (.A(_12923_),
    .B(_12919_),
    .C(_12921_),
    .Y(_12925_));
 sky130_fd_sc_hd__a21o_4 _43469_ (.A1(_12924_),
    .A2(_12925_),
    .B1(_12334_),
    .X(_12926_));
 sky130_fd_sc_hd__nand3_4 _43470_ (.A(_12924_),
    .B(_12925_),
    .C(_12337_),
    .Y(_12927_));
 sky130_fd_sc_hd__and2_4 _43471_ (.A(_12926_),
    .B(_12927_),
    .X(_12928_));
 sky130_vsdinv _43472_ (.A(_12928_),
    .Y(_12929_));
 sky130_fd_sc_hd__nand2_4 _43473_ (.A(_12906_),
    .B(_12929_),
    .Y(_12930_));
 sky130_fd_sc_hd__nand3_4 _43474_ (.A(_12928_),
    .B(_12903_),
    .C(_12905_),
    .Y(_12931_));
 sky130_fd_sc_hd__nand2_4 _43475_ (.A(_12930_),
    .B(_12931_),
    .Y(_12932_));
 sky130_fd_sc_hd__nand2_4 _43476_ (.A(_12871_),
    .B(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__nand3_4 _43477_ (.A(_12870_),
    .B(_12930_),
    .C(_12931_),
    .Y(_12934_));
 sky130_fd_sc_hd__a21boi_4 _43478_ (.A1(_12632_),
    .A2(_12609_),
    .B1_N(_12610_),
    .Y(_12935_));
 sky130_vsdinv _43479_ (.A(_12935_),
    .Y(_12936_));
 sky130_fd_sc_hd__a21oi_4 _43480_ (.A1(_12933_),
    .A2(_12934_),
    .B1(_12936_),
    .Y(_12937_));
 sky130_vsdinv _43481_ (.A(_12937_),
    .Y(_12938_));
 sky130_fd_sc_hd__nand3_4 _43482_ (.A(_12933_),
    .B(_12936_),
    .C(_12934_),
    .Y(_12939_));
 sky130_fd_sc_hd__nand2_4 _43483_ (.A(_12938_),
    .B(_12939_),
    .Y(_12940_));
 sky130_fd_sc_hd__nand2_4 _43484_ (.A(_12868_),
    .B(_12940_),
    .Y(_12941_));
 sky130_vsdinv _43485_ (.A(_12939_),
    .Y(_12942_));
 sky130_fd_sc_hd__nor2_4 _43486_ (.A(_12937_),
    .B(_12942_),
    .Y(_12943_));
 sky130_fd_sc_hd__nand3_4 _43487_ (.A(_12943_),
    .B(_12867_),
    .C(_12864_),
    .Y(_12944_));
 sky130_fd_sc_hd__nand2_4 _43488_ (.A(_12941_),
    .B(_12944_),
    .Y(_12945_));
 sky130_fd_sc_hd__a21boi_4 _43489_ (.A1(_12650_),
    .A2(_12572_),
    .B1_N(_12574_),
    .Y(_12946_));
 sky130_fd_sc_hd__nand2_4 _43490_ (.A(_12945_),
    .B(_12946_),
    .Y(_12947_));
 sky130_fd_sc_hd__a21boi_4 _43491_ (.A1(_12565_),
    .A2(_12569_),
    .B1_N(_12571_),
    .Y(_12948_));
 sky130_fd_sc_hd__o21ai_4 _43492_ (.A1(_12948_),
    .A2(_12646_),
    .B1(_12574_),
    .Y(_12949_));
 sky130_fd_sc_hd__nand3_4 _43493_ (.A(_12949_),
    .B(_12944_),
    .C(_12941_),
    .Y(_12950_));
 sky130_fd_sc_hd__nand2_4 _43494_ (.A(_12947_),
    .B(_12950_),
    .Y(_12951_));
 sky130_fd_sc_hd__a21boi_4 _43495_ (.A1(_12628_),
    .A2(_12658_),
    .B1_N(_12629_),
    .Y(_12952_));
 sky130_fd_sc_hd__a21boi_4 _43496_ (.A1(_12638_),
    .A2(_12643_),
    .B1_N(_12641_),
    .Y(_12953_));
 sky130_fd_sc_hd__xnor2_4 _43497_ (.A(_12952_),
    .B(_12953_),
    .Y(_12954_));
 sky130_fd_sc_hd__nand2_4 _43498_ (.A(_12951_),
    .B(_12954_),
    .Y(_12955_));
 sky130_vsdinv _43499_ (.A(_12954_),
    .Y(_12956_));
 sky130_fd_sc_hd__nand3_4 _43500_ (.A(_12947_),
    .B(_12950_),
    .C(_12956_),
    .Y(_12957_));
 sky130_fd_sc_hd__nand2_4 _43501_ (.A(_12955_),
    .B(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__a21boi_4 _43502_ (.A1(_12654_),
    .A2(_12663_),
    .B1_N(_12656_),
    .Y(_12959_));
 sky130_fd_sc_hd__nand2_4 _43503_ (.A(_12958_),
    .B(_12959_),
    .Y(_12960_));
 sky130_fd_sc_hd__a21boi_4 _43504_ (.A1(_12647_),
    .A2(_12651_),
    .B1_N(_12653_),
    .Y(_12961_));
 sky130_fd_sc_hd__o21ai_4 _43505_ (.A1(_12661_),
    .A2(_12961_),
    .B1(_12656_),
    .Y(_12962_));
 sky130_fd_sc_hd__nand3_4 _43506_ (.A(_12962_),
    .B(_12955_),
    .C(_12957_),
    .Y(_12963_));
 sky130_fd_sc_hd__nand2_4 _43507_ (.A(_12960_),
    .B(_12963_),
    .Y(_12964_));
 sky130_fd_sc_hd__a21oi_4 _43508_ (.A1(_12354_),
    .A2(_12349_),
    .B1(_12659_),
    .Y(_12965_));
 sky130_vsdinv _43509_ (.A(_12965_),
    .Y(_12966_));
 sky130_fd_sc_hd__nand2_4 _43510_ (.A(_12964_),
    .B(_12966_),
    .Y(_12967_));
 sky130_fd_sc_hd__nand3_4 _43511_ (.A(_12960_),
    .B(_12965_),
    .C(_12963_),
    .Y(_12968_));
 sky130_fd_sc_hd__nand2_4 _43512_ (.A(_12967_),
    .B(_12968_),
    .Y(_12969_));
 sky130_fd_sc_hd__a21boi_4 _43513_ (.A1(_12667_),
    .A2(_12671_),
    .B1_N(_12669_),
    .Y(_12970_));
 sky130_fd_sc_hd__nand2_4 _43514_ (.A(_12969_),
    .B(_12970_),
    .Y(_12971_));
 sky130_fd_sc_hd__nand2_4 _43515_ (.A(_12674_),
    .B(_12669_),
    .Y(_12972_));
 sky130_fd_sc_hd__nand3_4 _43516_ (.A(_12972_),
    .B(_12967_),
    .C(_12968_),
    .Y(_12973_));
 sky130_fd_sc_hd__nand2_4 _43517_ (.A(_12971_),
    .B(_12973_),
    .Y(_12974_));
 sky130_fd_sc_hd__o21ai_4 _43518_ (.A1(_12680_),
    .A2(_12686_),
    .B1(_12679_),
    .Y(_12975_));
 sky130_fd_sc_hd__xnor2_4 _43519_ (.A(_12974_),
    .B(_12975_),
    .Y(_01442_));
 sky130_fd_sc_hd__a21boi_4 _43520_ (.A1(_12690_),
    .A2(_12692_),
    .B1_N(_12693_),
    .Y(_12976_));
 sky130_vsdinv _43521_ (.A(_12976_),
    .Y(_12977_));
 sky130_fd_sc_hd__nand2_4 _43522_ (.A(_06247_),
    .B(_12390_),
    .Y(_12978_));
 sky130_fd_sc_hd__o21ai_4 _43523_ (.A1(_07939_),
    .A2(_11101_),
    .B1(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__nand2_4 _43524_ (.A(_03280_),
    .B(_03619_),
    .Y(_12980_));
 sky130_vsdinv _43525_ (.A(_12980_),
    .Y(_12981_));
 sky130_fd_sc_hd__nand4_4 _43526_ (.A(_03272_),
    .B(_08381_),
    .C(_11433_),
    .D(_12393_),
    .Y(_12982_));
 sky130_fd_sc_hd__nand3_4 _43527_ (.A(_12979_),
    .B(_12981_),
    .C(_12982_),
    .Y(_12983_));
 sky130_fd_sc_hd__nand2_4 _43528_ (.A(_12979_),
    .B(_12982_),
    .Y(_12984_));
 sky130_fd_sc_hd__nand2_4 _43529_ (.A(_12984_),
    .B(_12980_),
    .Y(_12985_));
 sky130_fd_sc_hd__nand3_4 _43530_ (.A(_12977_),
    .B(_12983_),
    .C(_12985_),
    .Y(_12986_));
 sky130_fd_sc_hd__nand2_4 _43531_ (.A(_12985_),
    .B(_12983_),
    .Y(_12987_));
 sky130_fd_sc_hd__nand2_4 _43532_ (.A(_12987_),
    .B(_12976_),
    .Y(_12988_));
 sky130_fd_sc_hd__nand2_4 _43533_ (.A(_12986_),
    .B(_12988_),
    .Y(_12989_));
 sky130_fd_sc_hd__nand2_4 _43534_ (.A(_10265_),
    .B(_11777_),
    .Y(_12990_));
 sky130_fd_sc_hd__nand2_4 _43535_ (.A(_07654_),
    .B(_10502_),
    .Y(_12991_));
 sky130_fd_sc_hd__nand2_4 _43536_ (.A(_12990_),
    .B(_12991_),
    .Y(_12992_));
 sky130_fd_sc_hd__nand4_4 _43537_ (.A(_08168_),
    .B(_08169_),
    .C(_12092_),
    .D(_12093_),
    .Y(_12993_));
 sky130_fd_sc_hd__nand2_4 _43538_ (.A(_07822_),
    .B(_11125_),
    .Y(_12994_));
 sky130_vsdinv _43539_ (.A(_12994_),
    .Y(_12995_));
 sky130_fd_sc_hd__a21oi_4 _43540_ (.A1(_12992_),
    .A2(_12993_),
    .B1(_12995_),
    .Y(_12996_));
 sky130_fd_sc_hd__nand3_4 _43541_ (.A(_12992_),
    .B(_12993_),
    .C(_12995_),
    .Y(_12997_));
 sky130_vsdinv _43542_ (.A(_12997_),
    .Y(_12998_));
 sky130_fd_sc_hd__nor2_4 _43543_ (.A(_12996_),
    .B(_12998_),
    .Y(_12999_));
 sky130_vsdinv _43544_ (.A(_12999_),
    .Y(_13000_));
 sky130_fd_sc_hd__nand2_4 _43545_ (.A(_12989_),
    .B(_13000_),
    .Y(_13001_));
 sky130_fd_sc_hd__nand3_4 _43546_ (.A(_12986_),
    .B(_12988_),
    .C(_12999_),
    .Y(_13002_));
 sky130_fd_sc_hd__nand2_4 _43547_ (.A(_13001_),
    .B(_13002_),
    .Y(_13003_));
 sky130_fd_sc_hd__nand3_4 _43548_ (.A(_13003_),
    .B(_12697_),
    .C(_12711_),
    .Y(_13004_));
 sky130_fd_sc_hd__nand2_4 _43549_ (.A(_12711_),
    .B(_12697_),
    .Y(_13005_));
 sky130_fd_sc_hd__nand3_4 _43550_ (.A(_13005_),
    .B(_13002_),
    .C(_13001_),
    .Y(_13006_));
 sky130_fd_sc_hd__nand2_4 _43551_ (.A(_13004_),
    .B(_13006_),
    .Y(_13007_));
 sky130_fd_sc_hd__nand2_4 _43552_ (.A(_07819_),
    .B(_10300_),
    .Y(_13008_));
 sky130_fd_sc_hd__nand2_4 _43553_ (.A(_07824_),
    .B(_10481_),
    .Y(_13009_));
 sky130_fd_sc_hd__nand2_4 _43554_ (.A(_13008_),
    .B(_13009_),
    .Y(_13010_));
 sky130_fd_sc_hd__buf_1 _43555_ (.A(_09760_),
    .X(_13011_));
 sky130_fd_sc_hd__nand4_4 _43556_ (.A(_11826_),
    .B(_10584_),
    .C(_13011_),
    .D(_11793_),
    .Y(_13012_));
 sky130_fd_sc_hd__nand2_4 _43557_ (.A(_03314_),
    .B(_03581_),
    .Y(_13013_));
 sky130_vsdinv _43558_ (.A(_13013_),
    .Y(_13014_));
 sky130_fd_sc_hd__a21o_4 _43559_ (.A1(_13010_),
    .A2(_13012_),
    .B1(_13014_),
    .X(_13015_));
 sky130_fd_sc_hd__nand3_4 _43560_ (.A(_13010_),
    .B(_13012_),
    .C(_13014_),
    .Y(_13016_));
 sky130_fd_sc_hd__a21boi_4 _43561_ (.A1(_12703_),
    .A2(_12706_),
    .B1_N(_12704_),
    .Y(_13017_));
 sky130_fd_sc_hd__a21boi_4 _43562_ (.A1(_13015_),
    .A2(_13016_),
    .B1_N(_13017_),
    .Y(_13018_));
 sky130_vsdinv _43563_ (.A(_13018_),
    .Y(_13019_));
 sky130_vsdinv _43564_ (.A(_13017_),
    .Y(_13020_));
 sky130_fd_sc_hd__nand3_4 _43565_ (.A(_13020_),
    .B(_13016_),
    .C(_13015_),
    .Y(_13021_));
 sky130_fd_sc_hd__a21boi_4 _43566_ (.A1(_12723_),
    .A2(_12726_),
    .B1_N(_12724_),
    .Y(_13022_));
 sky130_vsdinv _43567_ (.A(_13022_),
    .Y(_13023_));
 sky130_fd_sc_hd__a21oi_4 _43568_ (.A1(_13019_),
    .A2(_13021_),
    .B1(_13023_),
    .Y(_13024_));
 sky130_vsdinv _43569_ (.A(_13024_),
    .Y(_13025_));
 sky130_fd_sc_hd__nand3_4 _43570_ (.A(_13019_),
    .B(_13023_),
    .C(_13021_),
    .Y(_13026_));
 sky130_fd_sc_hd__nand2_4 _43571_ (.A(_13025_),
    .B(_13026_),
    .Y(_13027_));
 sky130_fd_sc_hd__nand2_4 _43572_ (.A(_13007_),
    .B(_13027_),
    .Y(_13028_));
 sky130_vsdinv _43573_ (.A(_13027_),
    .Y(_13029_));
 sky130_fd_sc_hd__nand3_4 _43574_ (.A(_13029_),
    .B(_13006_),
    .C(_13004_),
    .Y(_13030_));
 sky130_fd_sc_hd__nand2_4 _43575_ (.A(_13028_),
    .B(_13030_),
    .Y(_13031_));
 sky130_fd_sc_hd__maj3_4 _43576_ (.A(_12712_),
    .B(_12737_),
    .C(_12714_),
    .X(_13032_));
 sky130_fd_sc_hd__nand2_4 _43577_ (.A(_13031_),
    .B(_13032_),
    .Y(_13033_));
 sky130_fd_sc_hd__nand2_4 _43578_ (.A(_12739_),
    .B(_12717_),
    .Y(_13034_));
 sky130_fd_sc_hd__nand3_4 _43579_ (.A(_13034_),
    .B(_13030_),
    .C(_13028_),
    .Y(_13035_));
 sky130_fd_sc_hd__nand2_4 _43580_ (.A(_13033_),
    .B(_13035_),
    .Y(_13036_));
 sky130_fd_sc_hd__maj3_4 _43581_ (.A(_12748_),
    .B(_12752_),
    .C(_12749_),
    .X(_13037_));
 sky130_fd_sc_hd__nand2_4 _43582_ (.A(_07158_),
    .B(_11503_),
    .Y(_13038_));
 sky130_fd_sc_hd__nand2_4 _43583_ (.A(_07621_),
    .B(_11169_),
    .Y(_13039_));
 sky130_fd_sc_hd__nand2_4 _43584_ (.A(_13038_),
    .B(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__nand4_4 _43585_ (.A(_07858_),
    .B(_12458_),
    .C(_03570_),
    .D(_11503_),
    .Y(_13041_));
 sky130_fd_sc_hd__buf_1 _43586_ (.A(_11010_),
    .X(_13042_));
 sky130_fd_sc_hd__nand2_4 _43587_ (.A(_13042_),
    .B(_12754_),
    .Y(_13043_));
 sky130_fd_sc_hd__a21bo_4 _43588_ (.A1(_13040_),
    .A2(_13041_),
    .B1_N(_13043_),
    .X(_13044_));
 sky130_fd_sc_hd__nand4_4 _43589_ (.A(_13042_),
    .B(_13040_),
    .C(_13041_),
    .D(_03565_),
    .Y(_13045_));
 sky130_fd_sc_hd__nand2_4 _43590_ (.A(_13044_),
    .B(_13045_),
    .Y(_13046_));
 sky130_fd_sc_hd__nor2_4 _43591_ (.A(_13037_),
    .B(_13046_),
    .Y(_13047_));
 sky130_vsdinv _43592_ (.A(_13047_),
    .Y(_13048_));
 sky130_fd_sc_hd__nand2_4 _43593_ (.A(_13046_),
    .B(_13037_),
    .Y(_13049_));
 sky130_fd_sc_hd__nand2_4 _43594_ (.A(_08309_),
    .B(_12456_),
    .Y(_13050_));
 sky130_fd_sc_hd__buf_1 _43595_ (.A(_10619_),
    .X(_13051_));
 sky130_fd_sc_hd__nand2_4 _43596_ (.A(_13051_),
    .B(_11521_),
    .Y(_13052_));
 sky130_fd_sc_hd__o21ai_4 _43597_ (.A1(_03338_),
    .A2(_03559_),
    .B1(_13052_),
    .Y(_13053_));
 sky130_fd_sc_hd__buf_1 _43598_ (.A(_07630_),
    .X(_13054_));
 sky130_fd_sc_hd__buf_1 _43599_ (.A(_08194_),
    .X(_13055_));
 sky130_fd_sc_hd__nand4_4 _43600_ (.A(_13054_),
    .B(_13051_),
    .C(_11521_),
    .D(_13055_),
    .Y(_13056_));
 sky130_fd_sc_hd__nand2_4 _43601_ (.A(_13053_),
    .B(_13056_),
    .Y(_13057_));
 sky130_fd_sc_hd__xor2_4 _43602_ (.A(_13050_),
    .B(_13057_),
    .X(_13058_));
 sky130_fd_sc_hd__a21o_4 _43603_ (.A1(_13048_),
    .A2(_13049_),
    .B1(_13058_),
    .X(_13059_));
 sky130_fd_sc_hd__nand3_4 _43604_ (.A(_13048_),
    .B(_13058_),
    .C(_13049_),
    .Y(_13060_));
 sky130_fd_sc_hd__a21boi_4 _43605_ (.A1(_12731_),
    .A2(_12734_),
    .B1_N(_12732_),
    .Y(_13061_));
 sky130_vsdinv _43606_ (.A(_13061_),
    .Y(_13062_));
 sky130_fd_sc_hd__a21oi_4 _43607_ (.A1(_13059_),
    .A2(_13060_),
    .B1(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__nand3_4 _43608_ (.A(_13059_),
    .B(_13062_),
    .C(_13060_),
    .Y(_13064_));
 sky130_vsdinv _43609_ (.A(_13064_),
    .Y(_13065_));
 sky130_fd_sc_hd__a21oi_4 _43610_ (.A1(_12769_),
    .A2(_12759_),
    .B1(_12757_),
    .Y(_13066_));
 sky130_fd_sc_hd__o21ai_4 _43611_ (.A1(_13063_),
    .A2(_13065_),
    .B1(_13066_),
    .Y(_13067_));
 sky130_fd_sc_hd__a21o_4 _43612_ (.A1(_13059_),
    .A2(_13060_),
    .B1(_13062_),
    .X(_13068_));
 sky130_vsdinv _43613_ (.A(_13066_),
    .Y(_13069_));
 sky130_fd_sc_hd__nand3_4 _43614_ (.A(_13068_),
    .B(_13069_),
    .C(_13064_),
    .Y(_13070_));
 sky130_fd_sc_hd__nand2_4 _43615_ (.A(_13067_),
    .B(_13070_),
    .Y(_13071_));
 sky130_fd_sc_hd__nand2_4 _43616_ (.A(_13036_),
    .B(_13071_),
    .Y(_13072_));
 sky130_fd_sc_hd__nand4_4 _43617_ (.A(_13070_),
    .B(_13033_),
    .C(_13035_),
    .D(_13067_),
    .Y(_13073_));
 sky130_fd_sc_hd__nand2_4 _43618_ (.A(_13072_),
    .B(_13073_),
    .Y(_13074_));
 sky130_vsdinv _43619_ (.A(_12781_),
    .Y(_13075_));
 sky130_fd_sc_hd__nor2_4 _43620_ (.A(_12779_),
    .B(_13075_),
    .Y(_13076_));
 sky130_vsdinv _43621_ (.A(_12745_),
    .Y(_13077_));
 sky130_fd_sc_hd__a21oi_4 _43622_ (.A1(_13076_),
    .A2(_12744_),
    .B1(_13077_),
    .Y(_13078_));
 sky130_fd_sc_hd__nand2_4 _43623_ (.A(_13074_),
    .B(_13078_),
    .Y(_13079_));
 sky130_fd_sc_hd__a21o_4 _43624_ (.A1(_13076_),
    .A2(_12744_),
    .B1(_13077_),
    .X(_13080_));
 sky130_fd_sc_hd__nand3_4 _43625_ (.A(_13080_),
    .B(_13072_),
    .C(_13073_),
    .Y(_13081_));
 sky130_fd_sc_hd__nand2_4 _43626_ (.A(_13079_),
    .B(_13081_),
    .Y(_13082_));
 sky130_fd_sc_hd__nand2_4 _43627_ (.A(_12220_),
    .B(_07923_),
    .Y(_13083_));
 sky130_fd_sc_hd__buf_1 _43628_ (.A(_09087_),
    .X(_13084_));
 sky130_fd_sc_hd__nand2_4 _43629_ (.A(_13084_),
    .B(_07920_),
    .Y(_13085_));
 sky130_fd_sc_hd__nand2_4 _43630_ (.A(_13083_),
    .B(_13085_),
    .Y(_13086_));
 sky130_fd_sc_hd__buf_1 _43631_ (.A(_11030_),
    .X(_13087_));
 sky130_fd_sc_hd__buf_1 _43632_ (.A(_09830_),
    .X(_13088_));
 sky130_fd_sc_hd__buf_1 _43633_ (.A(_10990_),
    .X(_13089_));
 sky130_fd_sc_hd__nand4_4 _43634_ (.A(_13087_),
    .B(_13088_),
    .C(_13089_),
    .D(_03542_),
    .Y(_13090_));
 sky130_fd_sc_hd__nand2_4 _43635_ (.A(_10788_),
    .B(_03531_),
    .Y(_13091_));
 sky130_vsdinv _43636_ (.A(_13091_),
    .Y(_13092_));
 sky130_fd_sc_hd__a21o_4 _43637_ (.A1(_13086_),
    .A2(_13090_),
    .B1(_13092_),
    .X(_13093_));
 sky130_fd_sc_hd__nand3_4 _43638_ (.A(_13086_),
    .B(_13090_),
    .C(_13092_),
    .Y(_13094_));
 sky130_fd_sc_hd__nand2_4 _43639_ (.A(_13093_),
    .B(_13094_),
    .Y(_13095_));
 sky130_fd_sc_hd__a21o_4 _43640_ (.A1(_12763_),
    .A2(_12767_),
    .B1(_13095_),
    .X(_13096_));
 sky130_fd_sc_hd__a21boi_4 _43641_ (.A1(_12761_),
    .A2(_12765_),
    .B1_N(_12763_),
    .Y(_13097_));
 sky130_fd_sc_hd__nand2_4 _43642_ (.A(_13095_),
    .B(_13097_),
    .Y(_13098_));
 sky130_fd_sc_hd__a21boi_4 _43643_ (.A1(_12797_),
    .A2(_12800_),
    .B1_N(_12798_),
    .Y(_13099_));
 sky130_vsdinv _43644_ (.A(_13099_),
    .Y(_13100_));
 sky130_fd_sc_hd__a21o_4 _43645_ (.A1(_13096_),
    .A2(_13098_),
    .B1(_13100_),
    .X(_13101_));
 sky130_fd_sc_hd__nand3_4 _43646_ (.A(_13096_),
    .B(_13100_),
    .C(_13098_),
    .Y(_13102_));
 sky130_fd_sc_hd__maj3_4 _43647_ (.A(_12807_),
    .B(_12803_),
    .C(_12794_),
    .X(_13103_));
 sky130_vsdinv _43648_ (.A(_13103_),
    .Y(_13104_));
 sky130_fd_sc_hd__a21o_4 _43649_ (.A1(_13101_),
    .A2(_13102_),
    .B1(_13104_),
    .X(_13105_));
 sky130_fd_sc_hd__nand3_4 _43650_ (.A(_13104_),
    .B(_13101_),
    .C(_13102_),
    .Y(_13106_));
 sky130_fd_sc_hd__nand2_4 _43651_ (.A(_13105_),
    .B(_13106_),
    .Y(_13107_));
 sky130_fd_sc_hd__maj3_4 _43652_ (.A(_12822_),
    .B(_12816_),
    .C(_12818_),
    .X(_13108_));
 sky130_fd_sc_hd__nand2_4 _43653_ (.A(_12817_),
    .B(_12523_),
    .Y(_13109_));
 sky130_fd_sc_hd__nand2_4 _43654_ (.A(_09846_),
    .B(_07051_),
    .Y(_13110_));
 sky130_fd_sc_hd__nand2_4 _43655_ (.A(_13109_),
    .B(_13110_),
    .Y(_13111_));
 sky130_fd_sc_hd__buf_1 _43656_ (.A(_09843_),
    .X(_13112_));
 sky130_fd_sc_hd__nand4_4 _43657_ (.A(_12530_),
    .B(_13112_),
    .C(_11016_),
    .D(_11017_),
    .Y(_13113_));
 sky130_fd_sc_hd__buf_1 _43658_ (.A(_10083_),
    .X(_13114_));
 sky130_fd_sc_hd__nand2_4 _43659_ (.A(_13114_),
    .B(_03513_),
    .Y(_13115_));
 sky130_fd_sc_hd__a21bo_4 _43660_ (.A1(_13111_),
    .A2(_13113_),
    .B1_N(_13115_),
    .X(_13116_));
 sky130_fd_sc_hd__buf_1 _43661_ (.A(_12830_),
    .X(_13117_));
 sky130_fd_sc_hd__nand4_4 _43662_ (.A(_13117_),
    .B(_13111_),
    .C(_13113_),
    .D(_07747_),
    .Y(_13118_));
 sky130_fd_sc_hd__nand2_4 _43663_ (.A(_13116_),
    .B(_13118_),
    .Y(_13119_));
 sky130_fd_sc_hd__nor2_4 _43664_ (.A(_13108_),
    .B(_13119_),
    .Y(_13120_));
 sky130_fd_sc_hd__a21boi_4 _43665_ (.A1(_13118_),
    .A2(_13116_),
    .B1_N(_13108_),
    .Y(_13121_));
 sky130_fd_sc_hd__nand2_4 _43666_ (.A(_11988_),
    .B(_11590_),
    .Y(_13122_));
 sky130_fd_sc_hd__nand2_4 _43667_ (.A(_12832_),
    .B(_07537_),
    .Y(_13123_));
 sky130_fd_sc_hd__buf_1 _43668_ (.A(_10826_),
    .X(_13124_));
 sky130_fd_sc_hd__nand2_4 _43669_ (.A(_13124_),
    .B(_06506_),
    .Y(_13125_));
 sky130_fd_sc_hd__nand2_4 _43670_ (.A(_13123_),
    .B(_13125_),
    .Y(_13126_));
 sky130_fd_sc_hd__buf_1 _43671_ (.A(_10405_),
    .X(_13127_));
 sky130_fd_sc_hd__buf_1 _43672_ (.A(_10826_),
    .X(_13128_));
 sky130_fd_sc_hd__nand4_4 _43673_ (.A(_13127_),
    .B(_13128_),
    .C(_07542_),
    .D(_07544_),
    .Y(_13129_));
 sky130_fd_sc_hd__nand2_4 _43674_ (.A(_13126_),
    .B(_13129_),
    .Y(_13130_));
 sky130_fd_sc_hd__xor2_4 _43675_ (.A(_13122_),
    .B(_13130_),
    .X(_13131_));
 sky130_vsdinv _43676_ (.A(_13131_),
    .Y(_13132_));
 sky130_fd_sc_hd__o21a_4 _43677_ (.A1(_13120_),
    .A2(_13121_),
    .B1(_13132_),
    .X(_13133_));
 sky130_fd_sc_hd__nor2_4 _43678_ (.A(_13120_),
    .B(_13121_),
    .Y(_13134_));
 sky130_fd_sc_hd__nand2_4 _43679_ (.A(_13134_),
    .B(_13131_),
    .Y(_13135_));
 sky130_vsdinv _43680_ (.A(_13135_),
    .Y(_13136_));
 sky130_fd_sc_hd__nor2_4 _43681_ (.A(_13133_),
    .B(_13136_),
    .Y(_13137_));
 sky130_vsdinv _43682_ (.A(_13137_),
    .Y(_13138_));
 sky130_fd_sc_hd__nand2_4 _43683_ (.A(_13107_),
    .B(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__nand3_4 _43684_ (.A(_13105_),
    .B(_13137_),
    .C(_13106_),
    .Y(_13140_));
 sky130_fd_sc_hd__nand2_4 _43685_ (.A(_12781_),
    .B(_12776_),
    .Y(_13141_));
 sky130_fd_sc_hd__a21oi_4 _43686_ (.A1(_13139_),
    .A2(_13140_),
    .B1(_13141_),
    .Y(_13142_));
 sky130_fd_sc_hd__nand3_4 _43687_ (.A(_13141_),
    .B(_13139_),
    .C(_13140_),
    .Y(_13143_));
 sky130_vsdinv _43688_ (.A(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__a21boi_4 _43689_ (.A1(_12812_),
    .A2(_12843_),
    .B1_N(_12813_),
    .Y(_13145_));
 sky130_fd_sc_hd__o21ai_4 _43690_ (.A1(_13142_),
    .A2(_13144_),
    .B1(_13145_),
    .Y(_13146_));
 sky130_fd_sc_hd__nand2_4 _43691_ (.A(_13139_),
    .B(_13140_),
    .Y(_13147_));
 sky130_vsdinv _43692_ (.A(_13141_),
    .Y(_13148_));
 sky130_fd_sc_hd__nand2_4 _43693_ (.A(_13147_),
    .B(_13148_),
    .Y(_13149_));
 sky130_vsdinv _43694_ (.A(_13145_),
    .Y(_13150_));
 sky130_fd_sc_hd__nand3_4 _43695_ (.A(_13149_),
    .B(_13150_),
    .C(_13143_),
    .Y(_13151_));
 sky130_fd_sc_hd__nand2_4 _43696_ (.A(_13146_),
    .B(_13151_),
    .Y(_13152_));
 sky130_fd_sc_hd__nand2_4 _43697_ (.A(_13082_),
    .B(_13152_),
    .Y(_13153_));
 sky130_fd_sc_hd__a21oi_4 _43698_ (.A1(_13149_),
    .A2(_13143_),
    .B1(_13150_),
    .Y(_13154_));
 sky130_vsdinv _43699_ (.A(_13151_),
    .Y(_13155_));
 sky130_fd_sc_hd__nor2_4 _43700_ (.A(_13154_),
    .B(_13155_),
    .Y(_13156_));
 sky130_fd_sc_hd__nand3_4 _43701_ (.A(_13156_),
    .B(_13081_),
    .C(_13079_),
    .Y(_13157_));
 sky130_fd_sc_hd__nand2_4 _43702_ (.A(_13153_),
    .B(_13157_),
    .Y(_13158_));
 sky130_vsdinv _43703_ (.A(_12790_),
    .Y(_13159_));
 sky130_fd_sc_hd__a21oi_4 _43704_ (.A1(_12860_),
    .A2(_12787_),
    .B1(_13159_),
    .Y(_13160_));
 sky130_fd_sc_hd__nand2_4 _43705_ (.A(_13158_),
    .B(_13160_),
    .Y(_13161_));
 sky130_fd_sc_hd__a21o_4 _43706_ (.A1(_12860_),
    .A2(_12787_),
    .B1(_13159_),
    .X(_13162_));
 sky130_fd_sc_hd__nand3_4 _43707_ (.A(_13162_),
    .B(_13157_),
    .C(_13153_),
    .Y(_13163_));
 sky130_fd_sc_hd__nand2_4 _43708_ (.A(_13161_),
    .B(_13163_),
    .Y(_13164_));
 sky130_fd_sc_hd__maj3_4 _43709_ (.A(_12831_),
    .B(_12833_),
    .C(_12829_),
    .X(_13165_));
 sky130_fd_sc_hd__nand2_4 _43710_ (.A(_11334_),
    .B(_07470_),
    .Y(_13166_));
 sky130_fd_sc_hd__nand2_4 _43711_ (.A(_11684_),
    .B(_06600_),
    .Y(_13167_));
 sky130_fd_sc_hd__nand2_4 _43712_ (.A(_13166_),
    .B(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__buf_1 _43713_ (.A(_10845_),
    .X(_13169_));
 sky130_fd_sc_hd__nand4_4 _43714_ (.A(_13169_),
    .B(_11690_),
    .C(_06478_),
    .D(_03492_),
    .Y(_13170_));
 sky130_fd_sc_hd__nand2_4 _43715_ (.A(\pcpi_mul.rs1[32] ),
    .B(\pcpi_mul.rs2[6] ),
    .Y(_13171_));
 sky130_vsdinv _43716_ (.A(_13171_),
    .Y(_13172_));
 sky130_fd_sc_hd__buf_1 _43717_ (.A(_13172_),
    .X(_13173_));
 sky130_fd_sc_hd__a21o_4 _43718_ (.A1(_13168_),
    .A2(_13170_),
    .B1(_13173_),
    .X(_13174_));
 sky130_fd_sc_hd__buf_1 _43719_ (.A(_13173_),
    .X(_13175_));
 sky130_fd_sc_hd__nand3_4 _43720_ (.A(_13168_),
    .B(_13170_),
    .C(_13175_),
    .Y(_13176_));
 sky130_fd_sc_hd__nand2_4 _43721_ (.A(_13174_),
    .B(_13176_),
    .Y(_13177_));
 sky130_fd_sc_hd__nor2_4 _43722_ (.A(_13165_),
    .B(_13177_),
    .Y(_13178_));
 sky130_vsdinv _43723_ (.A(_13178_),
    .Y(_13179_));
 sky130_fd_sc_hd__nand2_4 _43724_ (.A(_13177_),
    .B(_13165_),
    .Y(_13180_));
 sky130_fd_sc_hd__a21boi_4 _43725_ (.A1(_12877_),
    .A2(_12881_),
    .B1_N(_12879_),
    .Y(_13181_));
 sky130_vsdinv _43726_ (.A(_13181_),
    .Y(_13182_));
 sky130_fd_sc_hd__a21o_4 _43727_ (.A1(_13179_),
    .A2(_13180_),
    .B1(_13182_),
    .X(_13183_));
 sky130_fd_sc_hd__nand3_4 _43728_ (.A(_13179_),
    .B(_13182_),
    .C(_13180_),
    .Y(_13184_));
 sky130_fd_sc_hd__nand2_4 _43729_ (.A(_13183_),
    .B(_13184_),
    .Y(_13185_));
 sky130_vsdinv _43730_ (.A(_12827_),
    .Y(_13186_));
 sky130_fd_sc_hd__o21a_4 _43731_ (.A1(_12828_),
    .A2(_12838_),
    .B1(_13186_),
    .X(_13187_));
 sky130_fd_sc_hd__nand2_4 _43732_ (.A(_13185_),
    .B(_13187_),
    .Y(_13188_));
 sky130_vsdinv _43733_ (.A(_13187_),
    .Y(_13189_));
 sky130_fd_sc_hd__nand3_4 _43734_ (.A(_13189_),
    .B(_13183_),
    .C(_13184_),
    .Y(_13190_));
 sky130_fd_sc_hd__a21oi_4 _43735_ (.A1(_12887_),
    .A2(_12891_),
    .B1(_12885_),
    .Y(_13191_));
 sky130_vsdinv _43736_ (.A(_13191_),
    .Y(_13192_));
 sky130_fd_sc_hd__a21o_4 _43737_ (.A1(_13188_),
    .A2(_13190_),
    .B1(_13192_),
    .X(_13193_));
 sky130_fd_sc_hd__nand3_4 _43738_ (.A(_13188_),
    .B(_13190_),
    .C(_13192_),
    .Y(_13194_));
 sky130_fd_sc_hd__nand2_4 _43739_ (.A(_13193_),
    .B(_13194_),
    .Y(_13195_));
 sky130_fd_sc_hd__a21boi_4 _43740_ (.A1(_12894_),
    .A2(_12899_),
    .B1_N(_12895_),
    .Y(_13196_));
 sky130_fd_sc_hd__nand2_4 _43741_ (.A(_13195_),
    .B(_13196_),
    .Y(_13197_));
 sky130_vsdinv _43742_ (.A(_13196_),
    .Y(_13198_));
 sky130_fd_sc_hd__nand3_4 _43743_ (.A(_13198_),
    .B(_13193_),
    .C(_13194_),
    .Y(_13199_));
 sky130_fd_sc_hd__nand2_4 _43744_ (.A(_13197_),
    .B(_13199_),
    .Y(_13200_));
 sky130_fd_sc_hd__nand4_4 _43745_ (.A(_03408_),
    .B(_03455_),
    .C(_03466_),
    .D(_03473_),
    .Y(_13201_));
 sky130_fd_sc_hd__buf_1 _43746_ (.A(_13201_),
    .X(_13202_));
 sky130_fd_sc_hd__o21a_4 _43747_ (.A1(_12612_),
    .A2(_12908_),
    .B1(_13201_),
    .X(_13203_));
 sky130_fd_sc_hd__xor2_4 _43748_ (.A(_13203_),
    .B(_12005_),
    .X(_13204_));
 sky130_vsdinv _43749_ (.A(_13204_),
    .Y(_13205_));
 sky130_fd_sc_hd__a21o_4 _43750_ (.A1(_12919_),
    .A2(_13202_),
    .B1(_13205_),
    .X(_13206_));
 sky130_fd_sc_hd__nand3_4 _43751_ (.A(_13205_),
    .B(_12919_),
    .C(_13202_),
    .Y(_13207_));
 sky130_fd_sc_hd__a21oi_4 _43752_ (.A1(_13206_),
    .A2(_13207_),
    .B1(_12335_),
    .Y(_13208_));
 sky130_fd_sc_hd__nand3_4 _43753_ (.A(_13206_),
    .B(_12337_),
    .C(_13207_),
    .Y(_13209_));
 sky130_vsdinv _43754_ (.A(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__nor2_4 _43755_ (.A(_13208_),
    .B(_13210_),
    .Y(_13211_));
 sky130_vsdinv _43756_ (.A(_13211_),
    .Y(_13212_));
 sky130_fd_sc_hd__nand2_4 _43757_ (.A(_13200_),
    .B(_13212_),
    .Y(_13213_));
 sky130_fd_sc_hd__nand3_4 _43758_ (.A(_13197_),
    .B(_13211_),
    .C(_13199_),
    .Y(_13214_));
 sky130_fd_sc_hd__nand2_4 _43759_ (.A(_12856_),
    .B(_12851_),
    .Y(_13215_));
 sky130_fd_sc_hd__a21oi_4 _43760_ (.A1(_13213_),
    .A2(_13214_),
    .B1(_13215_),
    .Y(_13216_));
 sky130_fd_sc_hd__nand3_4 _43761_ (.A(_13213_),
    .B(_13215_),
    .C(_13214_),
    .Y(_13217_));
 sky130_vsdinv _43762_ (.A(_13217_),
    .Y(_13218_));
 sky130_fd_sc_hd__a21boi_4 _43763_ (.A1(_12928_),
    .A2(_12903_),
    .B1_N(_12905_),
    .Y(_13219_));
 sky130_fd_sc_hd__o21ai_4 _43764_ (.A1(_13216_),
    .A2(_13218_),
    .B1(_13219_),
    .Y(_13220_));
 sky130_fd_sc_hd__nand2_4 _43765_ (.A(_13213_),
    .B(_13214_),
    .Y(_13221_));
 sky130_vsdinv _43766_ (.A(_13215_),
    .Y(_13222_));
 sky130_fd_sc_hd__nand2_4 _43767_ (.A(_13221_),
    .B(_13222_),
    .Y(_13223_));
 sky130_vsdinv _43768_ (.A(_13219_),
    .Y(_13224_));
 sky130_fd_sc_hd__nand3_4 _43769_ (.A(_13223_),
    .B(_13224_),
    .C(_13217_),
    .Y(_13225_));
 sky130_fd_sc_hd__nand2_4 _43770_ (.A(_13220_),
    .B(_13225_),
    .Y(_13226_));
 sky130_fd_sc_hd__nand2_4 _43771_ (.A(_13164_),
    .B(_13226_),
    .Y(_13227_));
 sky130_fd_sc_hd__a21oi_4 _43772_ (.A1(_13223_),
    .A2(_13217_),
    .B1(_13224_),
    .Y(_13228_));
 sky130_vsdinv _43773_ (.A(_13225_),
    .Y(_13229_));
 sky130_fd_sc_hd__nor2_4 _43774_ (.A(_13228_),
    .B(_13229_),
    .Y(_13230_));
 sky130_fd_sc_hd__nand3_4 _43775_ (.A(_13230_),
    .B(_13163_),
    .C(_13161_),
    .Y(_13231_));
 sky130_fd_sc_hd__nand2_4 _43776_ (.A(_13227_),
    .B(_13231_),
    .Y(_13232_));
 sky130_vsdinv _43777_ (.A(_12867_),
    .Y(_13233_));
 sky130_fd_sc_hd__a21oi_4 _43778_ (.A1(_12943_),
    .A2(_12864_),
    .B1(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__nand2_4 _43779_ (.A(_13232_),
    .B(_13234_),
    .Y(_13235_));
 sky130_fd_sc_hd__a21o_4 _43780_ (.A1(_12943_),
    .A2(_12864_),
    .B1(_13233_),
    .X(_13236_));
 sky130_fd_sc_hd__nand3_4 _43781_ (.A(_13236_),
    .B(_13231_),
    .C(_13227_),
    .Y(_13237_));
 sky130_fd_sc_hd__nand2_4 _43782_ (.A(_13235_),
    .B(_13237_),
    .Y(_13238_));
 sky130_fd_sc_hd__a21boi_4 _43783_ (.A1(_12924_),
    .A2(_12658_),
    .B1_N(_12925_),
    .Y(_13239_));
 sky130_vsdinv _43784_ (.A(_13239_),
    .Y(_13240_));
 sky130_fd_sc_hd__a21boi_4 _43785_ (.A1(_12933_),
    .A2(_12936_),
    .B1_N(_12934_),
    .Y(_13241_));
 sky130_fd_sc_hd__xor2_4 _43786_ (.A(_13240_),
    .B(_13241_),
    .X(_13242_));
 sky130_fd_sc_hd__nand2_4 _43787_ (.A(_13238_),
    .B(_13242_),
    .Y(_13243_));
 sky130_vsdinv _43788_ (.A(_13242_),
    .Y(_13244_));
 sky130_fd_sc_hd__nand3_4 _43789_ (.A(_13235_),
    .B(_13244_),
    .C(_13237_),
    .Y(_13245_));
 sky130_fd_sc_hd__nand2_4 _43790_ (.A(_13243_),
    .B(_13245_),
    .Y(_13246_));
 sky130_fd_sc_hd__a21boi_4 _43791_ (.A1(_12947_),
    .A2(_12956_),
    .B1_N(_12950_),
    .Y(_13247_));
 sky130_fd_sc_hd__nand2_4 _43792_ (.A(_13246_),
    .B(_13247_),
    .Y(_13248_));
 sky130_vsdinv _43793_ (.A(_13247_),
    .Y(_13249_));
 sky130_fd_sc_hd__nand3_4 _43794_ (.A(_13249_),
    .B(_13243_),
    .C(_13245_),
    .Y(_13250_));
 sky130_fd_sc_hd__nand2_4 _43795_ (.A(_13248_),
    .B(_13250_),
    .Y(_13251_));
 sky130_fd_sc_hd__a21oi_4 _43796_ (.A1(_12645_),
    .A2(_12641_),
    .B1(_12952_),
    .Y(_13252_));
 sky130_vsdinv _43797_ (.A(_13252_),
    .Y(_13253_));
 sky130_fd_sc_hd__nand2_4 _43798_ (.A(_13251_),
    .B(_13253_),
    .Y(_13254_));
 sky130_fd_sc_hd__nand3_4 _43799_ (.A(_13248_),
    .B(_13250_),
    .C(_13252_),
    .Y(_13255_));
 sky130_fd_sc_hd__nand2_4 _43800_ (.A(_13254_),
    .B(_13255_),
    .Y(_13256_));
 sky130_fd_sc_hd__nand2_4 _43801_ (.A(_12968_),
    .B(_12963_),
    .Y(_13257_));
 sky130_vsdinv _43802_ (.A(_13257_),
    .Y(_13258_));
 sky130_fd_sc_hd__nand2_4 _43803_ (.A(_13256_),
    .B(_13258_),
    .Y(_13259_));
 sky130_fd_sc_hd__nand3_4 _43804_ (.A(_13254_),
    .B(_13257_),
    .C(_13255_),
    .Y(_13260_));
 sky130_fd_sc_hd__nand2_4 _43805_ (.A(_13259_),
    .B(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__nand4_4 _43806_ (.A(_12679_),
    .B(_12677_),
    .C(_12971_),
    .D(_12973_),
    .Y(_13262_));
 sky130_fd_sc_hd__nand2_4 _43807_ (.A(_12973_),
    .B(_12679_),
    .Y(_13263_));
 sky130_fd_sc_hd__nand2_4 _43808_ (.A(_13263_),
    .B(_12971_),
    .Y(_13264_));
 sky130_fd_sc_hd__o21ai_4 _43809_ (.A1(_13262_),
    .A2(_12686_),
    .B1(_13264_),
    .Y(_13265_));
 sky130_fd_sc_hd__xnor2_4 _43810_ (.A(_13261_),
    .B(_13265_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_4 _43811_ (.A(_03276_),
    .B(_12393_),
    .Y(_13266_));
 sky130_fd_sc_hd__o21ai_4 _43812_ (.A1(_03281_),
    .A2(_03629_),
    .B1(_13266_),
    .Y(_13267_));
 sky130_fd_sc_hd__nand4_4 _43813_ (.A(_03276_),
    .B(_07758_),
    .C(_11105_),
    .D(_12076_),
    .Y(_13268_));
 sky130_fd_sc_hd__nand2_4 _43814_ (.A(_13267_),
    .B(_13268_),
    .Y(_13269_));
 sky130_fd_sc_hd__nand2_4 _43815_ (.A(_07465_),
    .B(_10955_),
    .Y(_13270_));
 sky130_fd_sc_hd__nand2_4 _43816_ (.A(_13269_),
    .B(_13270_),
    .Y(_13271_));
 sky130_vsdinv _43817_ (.A(_13270_),
    .Y(_13272_));
 sky130_fd_sc_hd__nand3_4 _43818_ (.A(_13267_),
    .B(_13272_),
    .C(_13268_),
    .Y(_13273_));
 sky130_fd_sc_hd__nand2_4 _43819_ (.A(_13271_),
    .B(_13273_),
    .Y(_13274_));
 sky130_fd_sc_hd__a21boi_4 _43820_ (.A1(_12979_),
    .A2(_12981_),
    .B1_N(_12982_),
    .Y(_13275_));
 sky130_fd_sc_hd__nand2_4 _43821_ (.A(_13274_),
    .B(_13275_),
    .Y(_13276_));
 sky130_vsdinv _43822_ (.A(_13275_),
    .Y(_13277_));
 sky130_fd_sc_hd__nand3_4 _43823_ (.A(_13277_),
    .B(_13273_),
    .C(_13271_),
    .Y(_13278_));
 sky130_fd_sc_hd__nand2_4 _43824_ (.A(_13276_),
    .B(_13278_),
    .Y(_13279_));
 sky130_fd_sc_hd__nand2_4 _43825_ (.A(_07952_),
    .B(_11447_),
    .Y(_13280_));
 sky130_fd_sc_hd__nand2_4 _43826_ (.A(_08607_),
    .B(_11449_),
    .Y(_13281_));
 sky130_fd_sc_hd__nand2_4 _43827_ (.A(_13280_),
    .B(_13281_),
    .Y(_13282_));
 sky130_fd_sc_hd__nand4_4 _43828_ (.A(_08394_),
    .B(_07822_),
    .C(_03606_),
    .D(_11777_),
    .Y(_13283_));
 sky130_fd_sc_hd__nand2_4 _43829_ (.A(_11826_),
    .B(_12095_),
    .Y(_13284_));
 sky130_vsdinv _43830_ (.A(_13284_),
    .Y(_13285_));
 sky130_fd_sc_hd__a21o_4 _43831_ (.A1(_13282_),
    .A2(_13283_),
    .B1(_13285_),
    .X(_13286_));
 sky130_fd_sc_hd__nand3_4 _43832_ (.A(_13282_),
    .B(_13283_),
    .C(_13285_),
    .Y(_13287_));
 sky130_fd_sc_hd__and2_4 _43833_ (.A(_13286_),
    .B(_13287_),
    .X(_13288_));
 sky130_vsdinv _43834_ (.A(_13288_),
    .Y(_13289_));
 sky130_fd_sc_hd__nand2_4 _43835_ (.A(_13279_),
    .B(_13289_),
    .Y(_13290_));
 sky130_fd_sc_hd__nand3_4 _43836_ (.A(_13276_),
    .B(_13278_),
    .C(_13288_),
    .Y(_13291_));
 sky130_fd_sc_hd__nand2_4 _43837_ (.A(_13290_),
    .B(_13291_),
    .Y(_13292_));
 sky130_fd_sc_hd__nand2_4 _43838_ (.A(_13002_),
    .B(_12986_),
    .Y(_13293_));
 sky130_vsdinv _43839_ (.A(_13293_),
    .Y(_13294_));
 sky130_fd_sc_hd__nand2_4 _43840_ (.A(_13292_),
    .B(_13294_),
    .Y(_13295_));
 sky130_fd_sc_hd__nand3_4 _43841_ (.A(_13293_),
    .B(_13290_),
    .C(_13291_),
    .Y(_13296_));
 sky130_fd_sc_hd__nand2_4 _43842_ (.A(_13295_),
    .B(_13296_),
    .Y(_13297_));
 sky130_fd_sc_hd__buf_1 _43843_ (.A(_03595_),
    .X(_13298_));
 sky130_fd_sc_hd__nand2_4 _43844_ (.A(_07005_),
    .B(_13298_),
    .Y(_13299_));
 sky130_fd_sc_hd__nand2_4 _43845_ (.A(_10989_),
    .B(_12427_),
    .Y(_13300_));
 sky130_fd_sc_hd__nand2_4 _43846_ (.A(_13299_),
    .B(_13300_),
    .Y(_13301_));
 sky130_fd_sc_hd__nand4_4 _43847_ (.A(_07147_),
    .B(_07299_),
    .C(_12430_),
    .D(_12431_),
    .Y(_13302_));
 sky130_fd_sc_hd__buf_1 _43848_ (.A(_09346_),
    .X(_13303_));
 sky130_fd_sc_hd__nand2_4 _43849_ (.A(_07302_),
    .B(_13303_),
    .Y(_13304_));
 sky130_vsdinv _43850_ (.A(_13304_),
    .Y(_13305_));
 sky130_fd_sc_hd__a21o_4 _43851_ (.A1(_13301_),
    .A2(_13302_),
    .B1(_13305_),
    .X(_13306_));
 sky130_fd_sc_hd__nand3_4 _43852_ (.A(_13301_),
    .B(_13302_),
    .C(_13305_),
    .Y(_13307_));
 sky130_fd_sc_hd__nand2_4 _43853_ (.A(_13306_),
    .B(_13307_),
    .Y(_13308_));
 sky130_fd_sc_hd__a21o_4 _43854_ (.A1(_12993_),
    .A2(_12997_),
    .B1(_13308_),
    .X(_13309_));
 sky130_fd_sc_hd__a21boi_4 _43855_ (.A1(_12992_),
    .A2(_12995_),
    .B1_N(_12993_),
    .Y(_13310_));
 sky130_fd_sc_hd__nand2_4 _43856_ (.A(_13308_),
    .B(_13310_),
    .Y(_13311_));
 sky130_fd_sc_hd__a21boi_4 _43857_ (.A1(_13010_),
    .A2(_13014_),
    .B1_N(_13012_),
    .Y(_13312_));
 sky130_vsdinv _43858_ (.A(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__a21oi_4 _43859_ (.A1(_13309_),
    .A2(_13311_),
    .B1(_13313_),
    .Y(_13314_));
 sky130_fd_sc_hd__nand3_4 _43860_ (.A(_13309_),
    .B(_13313_),
    .C(_13311_),
    .Y(_13315_));
 sky130_vsdinv _43861_ (.A(_13315_),
    .Y(_13316_));
 sky130_fd_sc_hd__nor2_4 _43862_ (.A(_13314_),
    .B(_13316_),
    .Y(_13317_));
 sky130_vsdinv _43863_ (.A(_13317_),
    .Y(_13318_));
 sky130_fd_sc_hd__nand2_4 _43864_ (.A(_13297_),
    .B(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__nand3_4 _43865_ (.A(_13295_),
    .B(_13317_),
    .C(_13296_),
    .Y(_13320_));
 sky130_fd_sc_hd__nand2_4 _43866_ (.A(_13319_),
    .B(_13320_),
    .Y(_13321_));
 sky130_fd_sc_hd__a21boi_4 _43867_ (.A1(_13029_),
    .A2(_13004_),
    .B1_N(_13006_),
    .Y(_13322_));
 sky130_fd_sc_hd__nand2_4 _43868_ (.A(_13321_),
    .B(_13322_),
    .Y(_13323_));
 sky130_fd_sc_hd__a21oi_4 _43869_ (.A1(_13002_),
    .A2(_13001_),
    .B1(_13005_),
    .Y(_13324_));
 sky130_fd_sc_hd__o21ai_4 _43870_ (.A1(_13027_),
    .A2(_13324_),
    .B1(_13006_),
    .Y(_13325_));
 sky130_fd_sc_hd__nand3_4 _43871_ (.A(_13325_),
    .B(_13320_),
    .C(_13319_),
    .Y(_13326_));
 sky130_fd_sc_hd__nand2_4 _43872_ (.A(_13323_),
    .B(_13326_),
    .Y(_13327_));
 sky130_fd_sc_hd__nand2_4 _43873_ (.A(_10605_),
    .B(_10537_),
    .Y(_13328_));
 sky130_fd_sc_hd__nand2_4 _43874_ (.A(_08032_),
    .B(_08631_),
    .Y(_13329_));
 sky130_fd_sc_hd__nand2_4 _43875_ (.A(_13328_),
    .B(_13329_),
    .Y(_13330_));
 sky130_fd_sc_hd__buf_1 _43876_ (.A(_08289_),
    .X(_13331_));
 sky130_fd_sc_hd__nand4_4 _43877_ (.A(_13331_),
    .B(_07875_),
    .C(_12156_),
    .D(_12157_),
    .Y(_13332_));
 sky130_fd_sc_hd__nand2_4 _43878_ (.A(_11015_),
    .B(_11175_),
    .Y(_13333_));
 sky130_fd_sc_hd__a21bo_4 _43879_ (.A1(_13330_),
    .A2(_13332_),
    .B1_N(_13333_),
    .X(_13334_));
 sky130_fd_sc_hd__nand4_4 _43880_ (.A(_13054_),
    .B(_13330_),
    .C(_13332_),
    .D(_12754_),
    .Y(_13335_));
 sky130_fd_sc_hd__nand2_4 _43881_ (.A(_13334_),
    .B(_13335_),
    .Y(_13336_));
 sky130_fd_sc_hd__a21o_4 _43882_ (.A1(_13041_),
    .A2(_13045_),
    .B1(_13336_),
    .X(_13337_));
 sky130_fd_sc_hd__nand3_4 _43883_ (.A(_13336_),
    .B(_13041_),
    .C(_13045_),
    .Y(_13338_));
 sky130_fd_sc_hd__a2bb2o_4 _43884_ (.A1_N(_03348_),
    .A2_N(_03553_),
    .B1(_10624_),
    .B2(_12142_),
    .X(_13339_));
 sky130_fd_sc_hd__buf_1 _43885_ (.A(_08733_),
    .X(_13340_));
 sky130_fd_sc_hd__nand4_4 _43886_ (.A(_13340_),
    .B(_08523_),
    .C(_11842_),
    .D(_11522_),
    .Y(_13341_));
 sky130_fd_sc_hd__buf_1 _43887_ (.A(_08752_),
    .X(_13342_));
 sky130_fd_sc_hd__nand2_4 _43888_ (.A(_13342_),
    .B(_12144_),
    .Y(_13343_));
 sky130_vsdinv _43889_ (.A(_13343_),
    .Y(_13344_));
 sky130_fd_sc_hd__a21oi_4 _43890_ (.A1(_13339_),
    .A2(_13341_),
    .B1(_13344_),
    .Y(_13345_));
 sky130_fd_sc_hd__nand3_4 _43891_ (.A(_13339_),
    .B(_13344_),
    .C(_13341_),
    .Y(_13346_));
 sky130_vsdinv _43892_ (.A(_13346_),
    .Y(_13347_));
 sky130_fd_sc_hd__nor2_4 _43893_ (.A(_13345_),
    .B(_13347_),
    .Y(_13348_));
 sky130_fd_sc_hd__a21o_4 _43894_ (.A1(_13337_),
    .A2(_13338_),
    .B1(_13348_),
    .X(_13349_));
 sky130_fd_sc_hd__nand3_4 _43895_ (.A(_13337_),
    .B(_13348_),
    .C(_13338_),
    .Y(_13350_));
 sky130_fd_sc_hd__nand2_4 _43896_ (.A(_13349_),
    .B(_13350_),
    .Y(_13351_));
 sky130_fd_sc_hd__o21a_4 _43897_ (.A1(_13022_),
    .A2(_13018_),
    .B1(_13021_),
    .X(_13352_));
 sky130_fd_sc_hd__nand2_4 _43898_ (.A(_13351_),
    .B(_13352_),
    .Y(_13353_));
 sky130_vsdinv _43899_ (.A(_13352_),
    .Y(_13354_));
 sky130_fd_sc_hd__nand3_4 _43900_ (.A(_13349_),
    .B(_13354_),
    .C(_13350_),
    .Y(_13355_));
 sky130_fd_sc_hd__a21oi_4 _43901_ (.A1(_13058_),
    .A2(_13049_),
    .B1(_13047_),
    .Y(_13356_));
 sky130_vsdinv _43902_ (.A(_13356_),
    .Y(_13357_));
 sky130_fd_sc_hd__a21o_4 _43903_ (.A1(_13353_),
    .A2(_13355_),
    .B1(_13357_),
    .X(_13358_));
 sky130_fd_sc_hd__nand3_4 _43904_ (.A(_13353_),
    .B(_13357_),
    .C(_13355_),
    .Y(_13359_));
 sky130_fd_sc_hd__nand2_4 _43905_ (.A(_13358_),
    .B(_13359_),
    .Y(_13360_));
 sky130_fd_sc_hd__nand2_4 _43906_ (.A(_13327_),
    .B(_13360_),
    .Y(_13361_));
 sky130_fd_sc_hd__a21oi_4 _43907_ (.A1(_13353_),
    .A2(_13355_),
    .B1(_13357_),
    .Y(_13362_));
 sky130_vsdinv _43908_ (.A(_13359_),
    .Y(_13363_));
 sky130_fd_sc_hd__nor2_4 _43909_ (.A(_13362_),
    .B(_13363_),
    .Y(_13364_));
 sky130_fd_sc_hd__nand3_4 _43910_ (.A(_13364_),
    .B(_13326_),
    .C(_13323_),
    .Y(_13365_));
 sky130_fd_sc_hd__nand2_4 _43911_ (.A(_13361_),
    .B(_13365_),
    .Y(_13366_));
 sky130_fd_sc_hd__a21oi_4 _43912_ (.A1(_13028_),
    .A2(_13030_),
    .B1(_13034_),
    .Y(_13367_));
 sky130_fd_sc_hd__o21a_4 _43913_ (.A1(_13071_),
    .A2(_13367_),
    .B1(_13035_),
    .X(_13368_));
 sky130_fd_sc_hd__nand2_4 _43914_ (.A(_13366_),
    .B(_13368_),
    .Y(_13369_));
 sky130_fd_sc_hd__o21ai_4 _43915_ (.A1(_13071_),
    .A2(_13367_),
    .B1(_13035_),
    .Y(_13370_));
 sky130_fd_sc_hd__nand3_4 _43916_ (.A(_13370_),
    .B(_13365_),
    .C(_13361_),
    .Y(_13371_));
 sky130_fd_sc_hd__nand2_4 _43917_ (.A(_13369_),
    .B(_13371_),
    .Y(_13372_));
 sky130_vsdinv _43918_ (.A(_13050_),
    .Y(_13373_));
 sky130_fd_sc_hd__nand3_4 _43919_ (.A(_13053_),
    .B(_13056_),
    .C(_13373_),
    .Y(_13374_));
 sky130_fd_sc_hd__nand2_4 _43920_ (.A(_08531_),
    .B(_07915_),
    .Y(_13375_));
 sky130_fd_sc_hd__buf_1 _43921_ (.A(_03361_),
    .X(_13376_));
 sky130_fd_sc_hd__nand2_4 _43922_ (.A(_13376_),
    .B(_07917_),
    .Y(_13377_));
 sky130_fd_sc_hd__nand2_4 _43923_ (.A(_13375_),
    .B(_13377_),
    .Y(_13378_));
 sky130_fd_sc_hd__nand4_4 _43924_ (.A(_13084_),
    .B(_11595_),
    .C(_07920_),
    .D(_11873_),
    .Y(_13379_));
 sky130_fd_sc_hd__nand2_4 _43925_ (.A(_10785_),
    .B(_07563_),
    .Y(_13380_));
 sky130_vsdinv _43926_ (.A(_13380_),
    .Y(_13381_));
 sky130_fd_sc_hd__a21o_4 _43927_ (.A1(_13378_),
    .A2(_13379_),
    .B1(_13381_),
    .X(_13382_));
 sky130_fd_sc_hd__nand3_4 _43928_ (.A(_13378_),
    .B(_13379_),
    .C(_13381_),
    .Y(_13383_));
 sky130_fd_sc_hd__nand2_4 _43929_ (.A(_13382_),
    .B(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__a21o_4 _43930_ (.A1(_13056_),
    .A2(_13374_),
    .B1(_13384_),
    .X(_13385_));
 sky130_fd_sc_hd__a21boi_4 _43931_ (.A1(_13053_),
    .A2(_13373_),
    .B1_N(_13056_),
    .Y(_13386_));
 sky130_fd_sc_hd__nand2_4 _43932_ (.A(_13384_),
    .B(_13386_),
    .Y(_13387_));
 sky130_fd_sc_hd__a21boi_4 _43933_ (.A1(_13086_),
    .A2(_13092_),
    .B1_N(_13090_),
    .Y(_13388_));
 sky130_vsdinv _43934_ (.A(_13388_),
    .Y(_13389_));
 sky130_fd_sc_hd__a21o_4 _43935_ (.A1(_13385_),
    .A2(_13387_),
    .B1(_13389_),
    .X(_13390_));
 sky130_fd_sc_hd__nand3_4 _43936_ (.A(_13385_),
    .B(_13389_),
    .C(_13387_),
    .Y(_13391_));
 sky130_fd_sc_hd__maj3_4 _43937_ (.A(_13097_),
    .B(_13095_),
    .C(_13099_),
    .X(_13392_));
 sky130_vsdinv _43938_ (.A(_13392_),
    .Y(_13393_));
 sky130_fd_sc_hd__a21o_4 _43939_ (.A1(_13390_),
    .A2(_13391_),
    .B1(_13393_),
    .X(_13394_));
 sky130_fd_sc_hd__nand3_4 _43940_ (.A(_13393_),
    .B(_13390_),
    .C(_13391_),
    .Y(_13395_));
 sky130_fd_sc_hd__nand2_4 _43941_ (.A(_13394_),
    .B(_13395_),
    .Y(_13396_));
 sky130_fd_sc_hd__nand2_4 _43942_ (.A(_09578_),
    .B(_12528_),
    .Y(_13397_));
 sky130_fd_sc_hd__nand2_4 _43943_ (.A(_10080_),
    .B(_07522_),
    .Y(_13398_));
 sky130_fd_sc_hd__nand2_4 _43944_ (.A(_13397_),
    .B(_13398_),
    .Y(_13399_));
 sky130_fd_sc_hd__nand4_4 _43945_ (.A(_10791_),
    .B(_12830_),
    .C(_11907_),
    .D(_11905_),
    .Y(_13400_));
 sky130_fd_sc_hd__nand4_4 _43946_ (.A(_12277_),
    .B(_13399_),
    .C(_13400_),
    .D(_11023_),
    .Y(_13401_));
 sky130_fd_sc_hd__nand2_4 _43947_ (.A(_11951_),
    .B(_08598_),
    .Y(_13402_));
 sky130_fd_sc_hd__a21bo_4 _43948_ (.A1(_13399_),
    .A2(_13400_),
    .B1_N(_13402_),
    .X(_13403_));
 sky130_fd_sc_hd__maj3_4 _43949_ (.A(_13115_),
    .B(_13109_),
    .C(_13110_),
    .X(_13404_));
 sky130_fd_sc_hd__a21boi_4 _43950_ (.A1(_13401_),
    .A2(_13403_),
    .B1_N(_13404_),
    .Y(_13405_));
 sky130_vsdinv _43951_ (.A(_13405_),
    .Y(_13406_));
 sky130_fd_sc_hd__nand2_4 _43952_ (.A(_13403_),
    .B(_13401_),
    .Y(_13407_));
 sky130_fd_sc_hd__nor2_4 _43953_ (.A(_13404_),
    .B(_13407_),
    .Y(_13408_));
 sky130_vsdinv _43954_ (.A(_13408_),
    .Y(_13409_));
 sky130_fd_sc_hd__buf_1 _43955_ (.A(_12308_),
    .X(_13410_));
 sky130_fd_sc_hd__nand2_4 _43956_ (.A(_13410_),
    .B(_03497_),
    .Y(_13411_));
 sky130_fd_sc_hd__buf_1 _43957_ (.A(_10827_),
    .X(_13412_));
 sky130_fd_sc_hd__a2bb2o_4 _43958_ (.A1_N(_03394_),
    .A2_N(_03502_),
    .B1(_13412_),
    .B2(_07038_),
    .X(_13413_));
 sky130_fd_sc_hd__nand4_4 _43959_ (.A(_13412_),
    .B(_10844_),
    .C(_06507_),
    .D(_07038_),
    .Y(_13414_));
 sky130_fd_sc_hd__nand2_4 _43960_ (.A(_13413_),
    .B(_13414_),
    .Y(_13415_));
 sky130_fd_sc_hd__xor2_4 _43961_ (.A(_13411_),
    .B(_13415_),
    .X(_13416_));
 sky130_fd_sc_hd__a21oi_4 _43962_ (.A1(_13406_),
    .A2(_13409_),
    .B1(_13416_),
    .Y(_13417_));
 sky130_fd_sc_hd__nand3_4 _43963_ (.A(_13416_),
    .B(_13406_),
    .C(_13409_),
    .Y(_13418_));
 sky130_vsdinv _43964_ (.A(_13418_),
    .Y(_13419_));
 sky130_fd_sc_hd__nor2_4 _43965_ (.A(_13417_),
    .B(_13419_),
    .Y(_13420_));
 sky130_vsdinv _43966_ (.A(_13420_),
    .Y(_13421_));
 sky130_fd_sc_hd__nand2_4 _43967_ (.A(_13396_),
    .B(_13421_),
    .Y(_13422_));
 sky130_fd_sc_hd__nand3_4 _43968_ (.A(_13394_),
    .B(_13420_),
    .C(_13395_),
    .Y(_13423_));
 sky130_fd_sc_hd__nand2_4 _43969_ (.A(_13422_),
    .B(_13423_),
    .Y(_13424_));
 sky130_fd_sc_hd__o21ai_4 _43970_ (.A1(_13066_),
    .A2(_13063_),
    .B1(_13064_),
    .Y(_13425_));
 sky130_vsdinv _43971_ (.A(_13425_),
    .Y(_13426_));
 sky130_fd_sc_hd__nand2_4 _43972_ (.A(_13424_),
    .B(_13426_),
    .Y(_13427_));
 sky130_fd_sc_hd__nand3_4 _43973_ (.A(_13422_),
    .B(_13425_),
    .C(_13423_),
    .Y(_13428_));
 sky130_fd_sc_hd__nand2_4 _43974_ (.A(_13427_),
    .B(_13428_),
    .Y(_13429_));
 sky130_fd_sc_hd__a21boi_4 _43975_ (.A1(_13105_),
    .A2(_13137_),
    .B1_N(_13106_),
    .Y(_13430_));
 sky130_fd_sc_hd__nand2_4 _43976_ (.A(_13429_),
    .B(_13430_),
    .Y(_13431_));
 sky130_vsdinv _43977_ (.A(_13430_),
    .Y(_13432_));
 sky130_fd_sc_hd__nand3_4 _43978_ (.A(_13427_),
    .B(_13432_),
    .C(_13428_),
    .Y(_13433_));
 sky130_fd_sc_hd__nand2_4 _43979_ (.A(_13431_),
    .B(_13433_),
    .Y(_13434_));
 sky130_fd_sc_hd__nand2_4 _43980_ (.A(_13372_),
    .B(_13434_),
    .Y(_13435_));
 sky130_fd_sc_hd__nand4_4 _43981_ (.A(_13433_),
    .B(_13369_),
    .C(_13431_),
    .D(_13371_),
    .Y(_13436_));
 sky130_fd_sc_hd__nand2_4 _43982_ (.A(_13435_),
    .B(_13436_),
    .Y(_13437_));
 sky130_fd_sc_hd__a21boi_4 _43983_ (.A1(_13156_),
    .A2(_13079_),
    .B1_N(_13081_),
    .Y(_13438_));
 sky130_fd_sc_hd__nand2_4 _43984_ (.A(_13437_),
    .B(_13438_),
    .Y(_13439_));
 sky130_fd_sc_hd__a21oi_4 _43985_ (.A1(_13072_),
    .A2(_13073_),
    .B1(_13080_),
    .Y(_13440_));
 sky130_fd_sc_hd__o21ai_4 _43986_ (.A1(_13152_),
    .A2(_13440_),
    .B1(_13081_),
    .Y(_13441_));
 sky130_fd_sc_hd__nand3_4 _43987_ (.A(_13441_),
    .B(_13436_),
    .C(_13435_),
    .Y(_13442_));
 sky130_fd_sc_hd__nand2_4 _43988_ (.A(_13439_),
    .B(_13442_),
    .Y(_13443_));
 sky130_fd_sc_hd__a21boi_4 _43989_ (.A1(_13188_),
    .A2(_13192_),
    .B1_N(_13190_),
    .Y(_13444_));
 sky130_vsdinv _43990_ (.A(_13444_),
    .Y(_13445_));
 sky130_fd_sc_hd__maj3_4 _43991_ (.A(_13123_),
    .B(_13125_),
    .C(_13122_),
    .X(_13446_));
 sky130_fd_sc_hd__nand2_4 _43992_ (.A(_11684_),
    .B(_06594_),
    .Y(_13447_));
 sky130_fd_sc_hd__nand2_4 _43993_ (.A(_11339_),
    .B(_07095_),
    .Y(_13448_));
 sky130_fd_sc_hd__nand2_4 _43994_ (.A(_13447_),
    .B(_13448_),
    .Y(_13449_));
 sky130_fd_sc_hd__nand4_4 _43995_ (.A(_11690_),
    .B(_12909_),
    .C(_06478_),
    .D(_06789_),
    .Y(_13450_));
 sky130_fd_sc_hd__a21o_4 _43996_ (.A1(_13449_),
    .A2(_13450_),
    .B1(_13173_),
    .X(_13451_));
 sky130_fd_sc_hd__nand3_4 _43997_ (.A(_13449_),
    .B(_13450_),
    .C(_13175_),
    .Y(_13452_));
 sky130_fd_sc_hd__nand2_4 _43998_ (.A(_13451_),
    .B(_13452_),
    .Y(_13453_));
 sky130_fd_sc_hd__nor2_4 _43999_ (.A(_13446_),
    .B(_13453_),
    .Y(_13454_));
 sky130_vsdinv _44000_ (.A(_13454_),
    .Y(_13455_));
 sky130_fd_sc_hd__nand2_4 _44001_ (.A(_13453_),
    .B(_13446_),
    .Y(_13456_));
 sky130_fd_sc_hd__a21boi_4 _44002_ (.A1(_13168_),
    .A2(_13175_),
    .B1_N(_13170_),
    .Y(_13457_));
 sky130_vsdinv _44003_ (.A(_13457_),
    .Y(_13458_));
 sky130_fd_sc_hd__a21o_4 _44004_ (.A1(_13455_),
    .A2(_13456_),
    .B1(_13458_),
    .X(_13459_));
 sky130_fd_sc_hd__nand3_4 _44005_ (.A(_13455_),
    .B(_13458_),
    .C(_13456_),
    .Y(_13460_));
 sky130_fd_sc_hd__nand2_4 _44006_ (.A(_13459_),
    .B(_13460_),
    .Y(_13461_));
 sky130_vsdinv _44007_ (.A(_13120_),
    .Y(_13462_));
 sky130_fd_sc_hd__o21a_4 _44008_ (.A1(_13121_),
    .A2(_13132_),
    .B1(_13462_),
    .X(_13463_));
 sky130_fd_sc_hd__nand2_4 _44009_ (.A(_13461_),
    .B(_13463_),
    .Y(_13464_));
 sky130_vsdinv _44010_ (.A(_13463_),
    .Y(_13465_));
 sky130_fd_sc_hd__nand3_4 _44011_ (.A(_13465_),
    .B(_13459_),
    .C(_13460_),
    .Y(_13466_));
 sky130_fd_sc_hd__a21oi_4 _44012_ (.A1(_13180_),
    .A2(_13182_),
    .B1(_13178_),
    .Y(_13467_));
 sky130_vsdinv _44013_ (.A(_13467_),
    .Y(_13468_));
 sky130_fd_sc_hd__nand3_4 _44014_ (.A(_13464_),
    .B(_13466_),
    .C(_13468_),
    .Y(_13469_));
 sky130_fd_sc_hd__nand2_4 _44015_ (.A(_13464_),
    .B(_13466_),
    .Y(_13470_));
 sky130_fd_sc_hd__nand2_4 _44016_ (.A(_13470_),
    .B(_13467_),
    .Y(_13471_));
 sky130_fd_sc_hd__nand3_4 _44017_ (.A(_13445_),
    .B(_13469_),
    .C(_13471_),
    .Y(_13472_));
 sky130_fd_sc_hd__nand2_4 _44018_ (.A(_13471_),
    .B(_13469_),
    .Y(_13473_));
 sky130_fd_sc_hd__nand2_4 _44019_ (.A(_13473_),
    .B(_13444_),
    .Y(_13474_));
 sky130_fd_sc_hd__nand2_4 _44020_ (.A(_13472_),
    .B(_13474_),
    .Y(_13475_));
 sky130_fd_sc_hd__a211o_4 _44021_ (.A1(_12002_),
    .A2(_12003_),
    .B1(_12612_),
    .C1(_12908_),
    .X(_13476_));
 sky130_fd_sc_hd__o21a_4 _44022_ (.A1(_12920_),
    .A2(_13201_),
    .B1(_13476_),
    .X(_13477_));
 sky130_fd_sc_hd__xor2_4 _44023_ (.A(_12334_),
    .B(_13477_),
    .X(_13478_));
 sky130_vsdinv _44024_ (.A(_13478_),
    .Y(_13479_));
 sky130_fd_sc_hd__buf_1 _44025_ (.A(_13479_),
    .X(_13480_));
 sky130_fd_sc_hd__nand2_4 _44026_ (.A(_13475_),
    .B(_13480_),
    .Y(_13481_));
 sky130_fd_sc_hd__buf_1 _44027_ (.A(_13478_),
    .X(_13482_));
 sky130_fd_sc_hd__buf_1 _44028_ (.A(_13482_),
    .X(_13483_));
 sky130_fd_sc_hd__nand3_4 _44029_ (.A(_13472_),
    .B(_13474_),
    .C(_13483_),
    .Y(_13484_));
 sky130_fd_sc_hd__nand2_4 _44030_ (.A(_13481_),
    .B(_13484_),
    .Y(_13485_));
 sky130_fd_sc_hd__o21ai_4 _44031_ (.A1(_13145_),
    .A2(_13142_),
    .B1(_13143_),
    .Y(_13486_));
 sky130_vsdinv _44032_ (.A(_13486_),
    .Y(_13487_));
 sky130_fd_sc_hd__nand2_4 _44033_ (.A(_13485_),
    .B(_13487_),
    .Y(_13488_));
 sky130_fd_sc_hd__nand3_4 _44034_ (.A(_13486_),
    .B(_13481_),
    .C(_13484_),
    .Y(_13489_));
 sky130_fd_sc_hd__buf_1 _44035_ (.A(_13489_),
    .X(_13490_));
 sky130_fd_sc_hd__a21boi_4 _44036_ (.A1(_13197_),
    .A2(_13211_),
    .B1_N(_13199_),
    .Y(_13491_));
 sky130_vsdinv _44037_ (.A(_13491_),
    .Y(_13492_));
 sky130_fd_sc_hd__a21o_4 _44038_ (.A1(_13488_),
    .A2(_13490_),
    .B1(_13492_),
    .X(_13493_));
 sky130_fd_sc_hd__nand3_4 _44039_ (.A(_13488_),
    .B(_13492_),
    .C(_13489_),
    .Y(_13494_));
 sky130_fd_sc_hd__nand2_4 _44040_ (.A(_13493_),
    .B(_13494_),
    .Y(_13495_));
 sky130_fd_sc_hd__nand2_4 _44041_ (.A(_13443_),
    .B(_13495_),
    .Y(_13496_));
 sky130_fd_sc_hd__a21oi_4 _44042_ (.A1(_13488_),
    .A2(_13490_),
    .B1(_13492_),
    .Y(_13497_));
 sky130_vsdinv _44043_ (.A(_13494_),
    .Y(_13498_));
 sky130_fd_sc_hd__nor2_4 _44044_ (.A(_13497_),
    .B(_13498_),
    .Y(_13499_));
 sky130_fd_sc_hd__nand3_4 _44045_ (.A(_13499_),
    .B(_13442_),
    .C(_13439_),
    .Y(_13500_));
 sky130_fd_sc_hd__nand2_4 _44046_ (.A(_13496_),
    .B(_13500_),
    .Y(_13501_));
 sky130_fd_sc_hd__a21boi_4 _44047_ (.A1(_13230_),
    .A2(_13161_),
    .B1_N(_13163_),
    .Y(_13502_));
 sky130_fd_sc_hd__nand2_4 _44048_ (.A(_13501_),
    .B(_13502_),
    .Y(_13503_));
 sky130_fd_sc_hd__a21oi_4 _44049_ (.A1(_13153_),
    .A2(_13157_),
    .B1(_13162_),
    .Y(_13504_));
 sky130_fd_sc_hd__o21ai_4 _44050_ (.A1(_13226_),
    .A2(_13504_),
    .B1(_13163_),
    .Y(_13505_));
 sky130_fd_sc_hd__nand3_4 _44051_ (.A(_13505_),
    .B(_13500_),
    .C(_13496_),
    .Y(_13506_));
 sky130_fd_sc_hd__nand2_4 _44052_ (.A(_13503_),
    .B(_13506_),
    .Y(_13507_));
 sky130_fd_sc_hd__o21ai_4 _44053_ (.A1(_12920_),
    .A2(_13202_),
    .B1(_13209_),
    .Y(_13508_));
 sky130_fd_sc_hd__a21oi_4 _44054_ (.A1(_13223_),
    .A2(_13224_),
    .B1(_13218_),
    .Y(_13509_));
 sky130_fd_sc_hd__xor2_4 _44055_ (.A(_13508_),
    .B(_13509_),
    .X(_13510_));
 sky130_fd_sc_hd__nand2_4 _44056_ (.A(_13507_),
    .B(_13510_),
    .Y(_13511_));
 sky130_vsdinv _44057_ (.A(_13510_),
    .Y(_13512_));
 sky130_fd_sc_hd__nand3_4 _44058_ (.A(_13503_),
    .B(_13506_),
    .C(_13512_),
    .Y(_13513_));
 sky130_fd_sc_hd__nand2_4 _44059_ (.A(_13511_),
    .B(_13513_),
    .Y(_13514_));
 sky130_fd_sc_hd__a21boi_4 _44060_ (.A1(_13235_),
    .A2(_13244_),
    .B1_N(_13237_),
    .Y(_13515_));
 sky130_fd_sc_hd__nand2_4 _44061_ (.A(_13514_),
    .B(_13515_),
    .Y(_13516_));
 sky130_fd_sc_hd__nand2_4 _44062_ (.A(_13245_),
    .B(_13237_),
    .Y(_13517_));
 sky130_fd_sc_hd__nand3_4 _44063_ (.A(_13517_),
    .B(_13513_),
    .C(_13511_),
    .Y(_13518_));
 sky130_fd_sc_hd__nand2_4 _44064_ (.A(_13516_),
    .B(_13518_),
    .Y(_13519_));
 sky130_fd_sc_hd__a21oi_4 _44065_ (.A1(_12939_),
    .A2(_12934_),
    .B1(_13239_),
    .Y(_13520_));
 sky130_vsdinv _44066_ (.A(_13520_),
    .Y(_13521_));
 sky130_fd_sc_hd__nand2_4 _44067_ (.A(_13519_),
    .B(_13521_),
    .Y(_13522_));
 sky130_fd_sc_hd__nand3_4 _44068_ (.A(_13516_),
    .B(_13518_),
    .C(_13520_),
    .Y(_13523_));
 sky130_fd_sc_hd__nand2_4 _44069_ (.A(_13522_),
    .B(_13523_),
    .Y(_13524_));
 sky130_fd_sc_hd__a21boi_4 _44070_ (.A1(_13248_),
    .A2(_13252_),
    .B1_N(_13250_),
    .Y(_13525_));
 sky130_fd_sc_hd__nand2_4 _44071_ (.A(_13524_),
    .B(_13525_),
    .Y(_13526_));
 sky130_fd_sc_hd__nand2_4 _44072_ (.A(_13255_),
    .B(_13250_),
    .Y(_13527_));
 sky130_fd_sc_hd__nand3_4 _44073_ (.A(_13527_),
    .B(_13523_),
    .C(_13522_),
    .Y(_13528_));
 sky130_fd_sc_hd__nand2_4 _44074_ (.A(_13526_),
    .B(_13528_),
    .Y(_13529_));
 sky130_vsdinv _44075_ (.A(_13260_),
    .Y(_13530_));
 sky130_fd_sc_hd__a21oi_4 _44076_ (.A1(_13265_),
    .A2(_13259_),
    .B1(_13530_),
    .Y(_13531_));
 sky130_fd_sc_hd__xor2_4 _44077_ (.A(_13529_),
    .B(_13531_),
    .X(_01444_));
 sky130_fd_sc_hd__a21oi_4 _44078_ (.A1(_13496_),
    .A2(_13500_),
    .B1(_13505_),
    .Y(_13532_));
 sky130_fd_sc_hd__o21ai_4 _44079_ (.A1(_13510_),
    .A2(_13532_),
    .B1(_13506_),
    .Y(_13533_));
 sky130_vsdinv _44080_ (.A(_13533_),
    .Y(_13534_));
 sky130_fd_sc_hd__nand2_4 _44081_ (.A(_07753_),
    .B(_11102_),
    .Y(_13535_));
 sky130_fd_sc_hd__o21ai_4 _44082_ (.A1(_07762_),
    .A2(_03633_),
    .B1(_13535_),
    .Y(_13536_));
 sky130_fd_sc_hd__nand4_4 _44083_ (.A(_03281_),
    .B(_06451_),
    .C(_12075_),
    .D(_12393_),
    .Y(_13537_));
 sky130_fd_sc_hd__nand2_4 _44084_ (.A(_13536_),
    .B(_13537_),
    .Y(_13538_));
 sky130_fd_sc_hd__nand2_4 _44085_ (.A(_03294_),
    .B(_03619_),
    .Y(_13539_));
 sky130_fd_sc_hd__nand2_4 _44086_ (.A(_13538_),
    .B(_13539_),
    .Y(_13540_));
 sky130_vsdinv _44087_ (.A(_13539_),
    .Y(_13541_));
 sky130_fd_sc_hd__nand3_4 _44088_ (.A(_13536_),
    .B(_13541_),
    .C(_13537_),
    .Y(_13542_));
 sky130_fd_sc_hd__nand2_4 _44089_ (.A(_13540_),
    .B(_13542_),
    .Y(_13543_));
 sky130_fd_sc_hd__nand3_4 _44090_ (.A(_13543_),
    .B(_13268_),
    .C(_13273_),
    .Y(_13544_));
 sky130_fd_sc_hd__nand2_4 _44091_ (.A(_13273_),
    .B(_13268_),
    .Y(_13545_));
 sky130_fd_sc_hd__nand3_4 _44092_ (.A(_13545_),
    .B(_13542_),
    .C(_13540_),
    .Y(_13546_));
 sky130_fd_sc_hd__nand2_4 _44093_ (.A(_13544_),
    .B(_13546_),
    .Y(_13547_));
 sky130_fd_sc_hd__nand2_4 _44094_ (.A(_06847_),
    .B(_10499_),
    .Y(_13548_));
 sky130_fd_sc_hd__nand2_4 _44095_ (.A(_06849_),
    .B(_10502_),
    .Y(_13549_));
 sky130_fd_sc_hd__nand2_4 _44096_ (.A(_13548_),
    .B(_13549_),
    .Y(_13550_));
 sky130_fd_sc_hd__nand4_4 _44097_ (.A(_07284_),
    .B(_08835_),
    .C(_12092_),
    .D(_12093_),
    .Y(_13551_));
 sky130_fd_sc_hd__nand2_4 _44098_ (.A(_07147_),
    .B(_10509_),
    .Y(_13552_));
 sky130_fd_sc_hd__a21bo_4 _44099_ (.A1(_13550_),
    .A2(_13551_),
    .B1_N(_13552_),
    .X(_13553_));
 sky130_fd_sc_hd__nand4_4 _44100_ (.A(_07006_),
    .B(_13550_),
    .C(_13551_),
    .D(_10513_),
    .Y(_13554_));
 sky130_fd_sc_hd__nand2_4 _44101_ (.A(_13553_),
    .B(_13554_),
    .Y(_13555_));
 sky130_fd_sc_hd__nand2_4 _44102_ (.A(_13547_),
    .B(_13555_),
    .Y(_13556_));
 sky130_vsdinv _44103_ (.A(_13555_),
    .Y(_13557_));
 sky130_fd_sc_hd__nand3_4 _44104_ (.A(_13544_),
    .B(_13557_),
    .C(_13546_),
    .Y(_13558_));
 sky130_fd_sc_hd__nand2_4 _44105_ (.A(_13556_),
    .B(_13558_),
    .Y(_13559_));
 sky130_fd_sc_hd__a21boi_4 _44106_ (.A1(_13276_),
    .A2(_13288_),
    .B1_N(_13278_),
    .Y(_13560_));
 sky130_fd_sc_hd__nand2_4 _44107_ (.A(_13559_),
    .B(_13560_),
    .Y(_13561_));
 sky130_fd_sc_hd__nand2_4 _44108_ (.A(_13291_),
    .B(_13278_),
    .Y(_13562_));
 sky130_fd_sc_hd__nand3_4 _44109_ (.A(_13562_),
    .B(_13558_),
    .C(_13556_),
    .Y(_13563_));
 sky130_fd_sc_hd__nand2_4 _44110_ (.A(_13561_),
    .B(_13563_),
    .Y(_13564_));
 sky130_fd_sc_hd__nand2_4 _44111_ (.A(_08470_),
    .B(_11793_),
    .Y(_13565_));
 sky130_fd_sc_hd__nand2_4 _44112_ (.A(_10198_),
    .B(_10922_),
    .Y(_13566_));
 sky130_fd_sc_hd__nand2_4 _44113_ (.A(_13565_),
    .B(_13566_),
    .Y(_13567_));
 sky130_fd_sc_hd__nand4_4 _44114_ (.A(_07422_),
    .B(_07439_),
    .C(_11797_),
    .D(_11142_),
    .Y(_13568_));
 sky130_fd_sc_hd__nand2_4 _44115_ (.A(_03325_),
    .B(_10927_),
    .Y(_13569_));
 sky130_vsdinv _44116_ (.A(_13569_),
    .Y(_13570_));
 sky130_fd_sc_hd__a21o_4 _44117_ (.A1(_13567_),
    .A2(_13568_),
    .B1(_13570_),
    .X(_13571_));
 sky130_fd_sc_hd__nand3_4 _44118_ (.A(_13567_),
    .B(_13568_),
    .C(_13570_),
    .Y(_13572_));
 sky130_fd_sc_hd__nand2_4 _44119_ (.A(_13571_),
    .B(_13572_),
    .Y(_13573_));
 sky130_fd_sc_hd__a21boi_4 _44120_ (.A1(_13282_),
    .A2(_13285_),
    .B1_N(_13283_),
    .Y(_13574_));
 sky130_fd_sc_hd__nand2_4 _44121_ (.A(_13573_),
    .B(_13574_),
    .Y(_13575_));
 sky130_vsdinv _44122_ (.A(_13574_),
    .Y(_13576_));
 sky130_fd_sc_hd__nand3_4 _44123_ (.A(_13576_),
    .B(_13571_),
    .C(_13572_),
    .Y(_13577_));
 sky130_fd_sc_hd__a21boi_4 _44124_ (.A1(_13301_),
    .A2(_13305_),
    .B1_N(_13302_),
    .Y(_13578_));
 sky130_vsdinv _44125_ (.A(_13578_),
    .Y(_13579_));
 sky130_fd_sc_hd__a21o_4 _44126_ (.A1(_13575_),
    .A2(_13577_),
    .B1(_13579_),
    .X(_13580_));
 sky130_fd_sc_hd__nand3_4 _44127_ (.A(_13575_),
    .B(_13577_),
    .C(_13579_),
    .Y(_13581_));
 sky130_fd_sc_hd__nand2_4 _44128_ (.A(_13580_),
    .B(_13581_),
    .Y(_13582_));
 sky130_fd_sc_hd__nand2_4 _44129_ (.A(_13564_),
    .B(_13582_),
    .Y(_13583_));
 sky130_vsdinv _44130_ (.A(_13582_),
    .Y(_13584_));
 sky130_fd_sc_hd__nand3_4 _44131_ (.A(_13561_),
    .B(_13584_),
    .C(_13563_),
    .Y(_13585_));
 sky130_fd_sc_hd__nand2_4 _44132_ (.A(_13583_),
    .B(_13585_),
    .Y(_13586_));
 sky130_vsdinv _44133_ (.A(_13296_),
    .Y(_13587_));
 sky130_fd_sc_hd__a21oi_4 _44134_ (.A1(_13295_),
    .A2(_13317_),
    .B1(_13587_),
    .Y(_13588_));
 sky130_fd_sc_hd__nand2_4 _44135_ (.A(_13586_),
    .B(_13588_),
    .Y(_13589_));
 sky130_fd_sc_hd__a21o_4 _44136_ (.A1(_13295_),
    .A2(_13317_),
    .B1(_13587_),
    .X(_13590_));
 sky130_fd_sc_hd__nand3_4 _44137_ (.A(_13590_),
    .B(_13583_),
    .C(_13585_),
    .Y(_13591_));
 sky130_fd_sc_hd__nand2_4 _44138_ (.A(_13589_),
    .B(_13591_),
    .Y(_13592_));
 sky130_fd_sc_hd__maj3_4 _44139_ (.A(_13328_),
    .B(_13333_),
    .C(_13329_),
    .X(_13593_));
 sky130_fd_sc_hd__nand2_4 _44140_ (.A(_07626_),
    .B(_03576_),
    .Y(_13594_));
 sky130_fd_sc_hd__nand2_4 _44141_ (.A(_07871_),
    .B(_10536_),
    .Y(_13595_));
 sky130_fd_sc_hd__nand2_4 _44142_ (.A(_13594_),
    .B(_13595_),
    .Y(_13596_));
 sky130_fd_sc_hd__nand4_4 _44143_ (.A(_07875_),
    .B(_08051_),
    .C(_11829_),
    .D(_11824_),
    .Y(_13597_));
 sky130_fd_sc_hd__nand2_4 _44144_ (.A(_08052_),
    .B(_10887_),
    .Y(_13598_));
 sky130_vsdinv _44145_ (.A(_13598_),
    .Y(_13599_));
 sky130_fd_sc_hd__a21o_4 _44146_ (.A1(_13596_),
    .A2(_13597_),
    .B1(_13599_),
    .X(_13600_));
 sky130_fd_sc_hd__nand3_4 _44147_ (.A(_13596_),
    .B(_13597_),
    .C(_13599_),
    .Y(_13601_));
 sky130_fd_sc_hd__nand2_4 _44148_ (.A(_13600_),
    .B(_13601_),
    .Y(_13602_));
 sky130_fd_sc_hd__nor2_4 _44149_ (.A(_13593_),
    .B(_13602_),
    .Y(_13603_));
 sky130_vsdinv _44150_ (.A(_13603_),
    .Y(_13604_));
 sky130_fd_sc_hd__nand2_4 _44151_ (.A(_13602_),
    .B(_13593_),
    .Y(_13605_));
 sky130_fd_sc_hd__nand2_4 _44152_ (.A(_13088_),
    .B(_11514_),
    .Y(_13606_));
 sky130_fd_sc_hd__nand2_4 _44153_ (.A(_11243_),
    .B(_11516_),
    .Y(_13607_));
 sky130_fd_sc_hd__nand2_4 _44154_ (.A(_13087_),
    .B(_11518_),
    .Y(_13608_));
 sky130_fd_sc_hd__nand2_4 _44155_ (.A(_13607_),
    .B(_13608_),
    .Y(_13609_));
 sky130_fd_sc_hd__buf_1 _44156_ (.A(_11034_),
    .X(_13610_));
 sky130_fd_sc_hd__buf_1 _44157_ (.A(_11842_),
    .X(_13611_));
 sky130_fd_sc_hd__nand4_4 _44158_ (.A(_11910_),
    .B(_13610_),
    .C(_13611_),
    .D(_11523_),
    .Y(_13612_));
 sky130_fd_sc_hd__nand2_4 _44159_ (.A(_13609_),
    .B(_13612_),
    .Y(_13613_));
 sky130_fd_sc_hd__xor2_4 _44160_ (.A(_13606_),
    .B(_13613_),
    .X(_13614_));
 sky130_fd_sc_hd__a21oi_4 _44161_ (.A1(_13604_),
    .A2(_13605_),
    .B1(_13614_),
    .Y(_13615_));
 sky130_fd_sc_hd__nand3_4 _44162_ (.A(_13604_),
    .B(_13614_),
    .C(_13605_),
    .Y(_13616_));
 sky130_vsdinv _44163_ (.A(_13616_),
    .Y(_13617_));
 sky130_fd_sc_hd__maj3_4 _44164_ (.A(_13312_),
    .B(_13308_),
    .C(_13310_),
    .X(_13618_));
 sky130_fd_sc_hd__o21ai_4 _44165_ (.A1(_13615_),
    .A2(_13617_),
    .B1(_13618_),
    .Y(_13619_));
 sky130_vsdinv _44166_ (.A(_13615_),
    .Y(_13620_));
 sky130_vsdinv _44167_ (.A(_13618_),
    .Y(_13621_));
 sky130_fd_sc_hd__nand3_4 _44168_ (.A(_13620_),
    .B(_13621_),
    .C(_13616_),
    .Y(_13622_));
 sky130_fd_sc_hd__a21boi_4 _44169_ (.A1(_13348_),
    .A2(_13338_),
    .B1_N(_13337_),
    .Y(_13623_));
 sky130_vsdinv _44170_ (.A(_13623_),
    .Y(_13624_));
 sky130_fd_sc_hd__a21oi_4 _44171_ (.A1(_13619_),
    .A2(_13622_),
    .B1(_13624_),
    .Y(_13625_));
 sky130_vsdinv _44172_ (.A(_13625_),
    .Y(_13626_));
 sky130_fd_sc_hd__nand3_4 _44173_ (.A(_13619_),
    .B(_13622_),
    .C(_13624_),
    .Y(_13627_));
 sky130_fd_sc_hd__nand2_4 _44174_ (.A(_13626_),
    .B(_13627_),
    .Y(_13628_));
 sky130_fd_sc_hd__nand2_4 _44175_ (.A(_13592_),
    .B(_13628_),
    .Y(_13629_));
 sky130_vsdinv _44176_ (.A(_13627_),
    .Y(_13630_));
 sky130_fd_sc_hd__nor2_4 _44177_ (.A(_13625_),
    .B(_13630_),
    .Y(_13631_));
 sky130_fd_sc_hd__nand3_4 _44178_ (.A(_13631_),
    .B(_13591_),
    .C(_13589_),
    .Y(_13632_));
 sky130_fd_sc_hd__nand2_4 _44179_ (.A(_13629_),
    .B(_13632_),
    .Y(_13633_));
 sky130_fd_sc_hd__a21boi_4 _44180_ (.A1(_13364_),
    .A2(_13323_),
    .B1_N(_13326_),
    .Y(_13634_));
 sky130_fd_sc_hd__nand2_4 _44181_ (.A(_13633_),
    .B(_13634_),
    .Y(_13635_));
 sky130_fd_sc_hd__a21oi_4 _44182_ (.A1(_13319_),
    .A2(_13320_),
    .B1(_13325_),
    .Y(_13636_));
 sky130_fd_sc_hd__o21ai_4 _44183_ (.A1(_13636_),
    .A2(_13360_),
    .B1(_13326_),
    .Y(_13637_));
 sky130_fd_sc_hd__nand3_4 _44184_ (.A(_13637_),
    .B(_13632_),
    .C(_13629_),
    .Y(_13638_));
 sky130_fd_sc_hd__nand2_4 _44185_ (.A(_13635_),
    .B(_13638_),
    .Y(_13639_));
 sky130_fd_sc_hd__nand2_4 _44186_ (.A(_13376_),
    .B(_08358_),
    .Y(_13640_));
 sky130_fd_sc_hd__nand2_4 _44187_ (.A(_09574_),
    .B(_08357_),
    .Y(_13641_));
 sky130_fd_sc_hd__nand2_4 _44188_ (.A(_13640_),
    .B(_13641_),
    .Y(_13642_));
 sky130_fd_sc_hd__buf_1 _44189_ (.A(_08568_),
    .X(_13643_));
 sky130_fd_sc_hd__buf_1 _44190_ (.A(_08566_),
    .X(_13644_));
 sky130_fd_sc_hd__nand4_4 _44191_ (.A(_10783_),
    .B(_11287_),
    .C(_13643_),
    .D(_13644_),
    .Y(_13645_));
 sky130_fd_sc_hd__nand2_4 _44192_ (.A(_09578_),
    .B(_07720_),
    .Y(_13646_));
 sky130_vsdinv _44193_ (.A(_13646_),
    .Y(_13647_));
 sky130_fd_sc_hd__a21o_4 _44194_ (.A1(_13642_),
    .A2(_13645_),
    .B1(_13647_),
    .X(_13648_));
 sky130_fd_sc_hd__nand3_4 _44195_ (.A(_13642_),
    .B(_13645_),
    .C(_13647_),
    .Y(_13649_));
 sky130_fd_sc_hd__nand2_4 _44196_ (.A(_13648_),
    .B(_13649_),
    .Y(_13650_));
 sky130_fd_sc_hd__a21o_4 _44197_ (.A1(_13346_),
    .A2(_13341_),
    .B1(_13650_),
    .X(_13651_));
 sky130_fd_sc_hd__nand3_4 _44198_ (.A(_13650_),
    .B(_13346_),
    .C(_13341_),
    .Y(_13652_));
 sky130_fd_sc_hd__a21boi_4 _44199_ (.A1(_13378_),
    .A2(_13381_),
    .B1_N(_13379_),
    .Y(_13653_));
 sky130_vsdinv _44200_ (.A(_13653_),
    .Y(_13654_));
 sky130_fd_sc_hd__a21o_4 _44201_ (.A1(_13651_),
    .A2(_13652_),
    .B1(_13654_),
    .X(_13655_));
 sky130_fd_sc_hd__nand3_4 _44202_ (.A(_13651_),
    .B(_13654_),
    .C(_13652_),
    .Y(_13656_));
 sky130_fd_sc_hd__nand2_4 _44203_ (.A(_13655_),
    .B(_13656_),
    .Y(_13657_));
 sky130_fd_sc_hd__maj3_4 _44204_ (.A(_13388_),
    .B(_13384_),
    .C(_13386_),
    .X(_13658_));
 sky130_fd_sc_hd__nand2_4 _44205_ (.A(_13657_),
    .B(_13658_),
    .Y(_13659_));
 sky130_vsdinv _44206_ (.A(_13658_),
    .Y(_13660_));
 sky130_fd_sc_hd__nand3_4 _44207_ (.A(_13655_),
    .B(_13660_),
    .C(_13656_),
    .Y(_13661_));
 sky130_fd_sc_hd__nand2_4 _44208_ (.A(_13659_),
    .B(_13661_),
    .Y(_13662_));
 sky130_fd_sc_hd__maj3_4 _44209_ (.A(_13402_),
    .B(_13397_),
    .C(_13398_),
    .X(_13663_));
 sky130_fd_sc_hd__nand2_4 _44210_ (.A(_09580_),
    .B(_12523_),
    .Y(_13664_));
 sky130_fd_sc_hd__nand2_4 _44211_ (.A(_03383_),
    .B(_07051_),
    .Y(_13665_));
 sky130_fd_sc_hd__nand2_4 _44212_ (.A(_13664_),
    .B(_13665_),
    .Y(_13666_));
 sky130_fd_sc_hd__nand4_4 _44213_ (.A(_11639_),
    .B(_12832_),
    .C(_11016_),
    .D(_11017_),
    .Y(_13667_));
 sky130_fd_sc_hd__nand2_4 _44214_ (.A(_13124_),
    .B(_07744_),
    .Y(_13668_));
 sky130_vsdinv _44215_ (.A(_13668_),
    .Y(_13669_));
 sky130_fd_sc_hd__a21o_4 _44216_ (.A1(_13666_),
    .A2(_13667_),
    .B1(_13669_),
    .X(_13670_));
 sky130_fd_sc_hd__nand3_4 _44217_ (.A(_13666_),
    .B(_13667_),
    .C(_13669_),
    .Y(_13671_));
 sky130_fd_sc_hd__nand2_4 _44218_ (.A(_13670_),
    .B(_13671_),
    .Y(_13672_));
 sky130_fd_sc_hd__nor2_4 _44219_ (.A(_13663_),
    .B(_13672_),
    .Y(_13673_));
 sky130_fd_sc_hd__a21boi_4 _44220_ (.A1(_13670_),
    .A2(_13671_),
    .B1_N(_13663_),
    .Y(_13674_));
 sky130_fd_sc_hd__nand2_4 _44221_ (.A(_11337_),
    .B(_11590_),
    .Y(_13675_));
 sky130_fd_sc_hd__nand2_4 _44222_ (.A(_11988_),
    .B(_07215_),
    .Y(_13676_));
 sky130_fd_sc_hd__nand2_4 _44223_ (.A(_10846_),
    .B(_07213_),
    .Y(_13677_));
 sky130_fd_sc_hd__nand2_4 _44224_ (.A(_13676_),
    .B(_13677_),
    .Y(_13678_));
 sky130_fd_sc_hd__nand4_4 _44225_ (.A(_10840_),
    .B(_13169_),
    .C(_06888_),
    .D(_06894_),
    .Y(_13679_));
 sky130_fd_sc_hd__nand2_4 _44226_ (.A(_13678_),
    .B(_13679_),
    .Y(_13680_));
 sky130_fd_sc_hd__xor2_4 _44227_ (.A(_13675_),
    .B(_13680_),
    .X(_13681_));
 sky130_vsdinv _44228_ (.A(_13681_),
    .Y(_13682_));
 sky130_fd_sc_hd__o21a_4 _44229_ (.A1(_13673_),
    .A2(_13674_),
    .B1(_13682_),
    .X(_13683_));
 sky130_fd_sc_hd__nor2_4 _44230_ (.A(_13673_),
    .B(_13674_),
    .Y(_13684_));
 sky130_fd_sc_hd__nand2_4 _44231_ (.A(_13684_),
    .B(_13681_),
    .Y(_13685_));
 sky130_vsdinv _44232_ (.A(_13685_),
    .Y(_13686_));
 sky130_fd_sc_hd__nor2_4 _44233_ (.A(_13683_),
    .B(_13686_),
    .Y(_13687_));
 sky130_vsdinv _44234_ (.A(_13687_),
    .Y(_13688_));
 sky130_fd_sc_hd__nand2_4 _44235_ (.A(_13662_),
    .B(_13688_),
    .Y(_13689_));
 sky130_fd_sc_hd__nand3_4 _44236_ (.A(_13659_),
    .B(_13687_),
    .C(_13661_),
    .Y(_13690_));
 sky130_fd_sc_hd__nand2_4 _44237_ (.A(_13689_),
    .B(_13690_),
    .Y(_13691_));
 sky130_vsdinv _44238_ (.A(_13355_),
    .Y(_13692_));
 sky130_fd_sc_hd__a21oi_4 _44239_ (.A1(_13353_),
    .A2(_13357_),
    .B1(_13692_),
    .Y(_13693_));
 sky130_fd_sc_hd__nand2_4 _44240_ (.A(_13691_),
    .B(_13693_),
    .Y(_13694_));
 sky130_vsdinv _44241_ (.A(_13693_),
    .Y(_13695_));
 sky130_fd_sc_hd__nand3_4 _44242_ (.A(_13695_),
    .B(_13689_),
    .C(_13690_),
    .Y(_13696_));
 sky130_fd_sc_hd__a21boi_4 _44243_ (.A1(_13394_),
    .A2(_13420_),
    .B1_N(_13395_),
    .Y(_13697_));
 sky130_vsdinv _44244_ (.A(_13697_),
    .Y(_13698_));
 sky130_fd_sc_hd__a21o_4 _44245_ (.A1(_13694_),
    .A2(_13696_),
    .B1(_13698_),
    .X(_13699_));
 sky130_fd_sc_hd__nand3_4 _44246_ (.A(_13694_),
    .B(_13696_),
    .C(_13698_),
    .Y(_13700_));
 sky130_fd_sc_hd__nand2_4 _44247_ (.A(_13699_),
    .B(_13700_),
    .Y(_13701_));
 sky130_fd_sc_hd__nand2_4 _44248_ (.A(_13639_),
    .B(_13701_),
    .Y(_13702_));
 sky130_fd_sc_hd__nand4_4 _44249_ (.A(_13700_),
    .B(_13635_),
    .C(_13699_),
    .D(_13638_),
    .Y(_13703_));
 sky130_fd_sc_hd__nand2_4 _44250_ (.A(_13702_),
    .B(_13703_),
    .Y(_13704_));
 sky130_fd_sc_hd__a21oi_4 _44251_ (.A1(_13361_),
    .A2(_13365_),
    .B1(_13370_),
    .Y(_13705_));
 sky130_fd_sc_hd__o21a_4 _44252_ (.A1(_13434_),
    .A2(_13705_),
    .B1(_13371_),
    .X(_13706_));
 sky130_fd_sc_hd__nand2_4 _44253_ (.A(_13704_),
    .B(_13706_),
    .Y(_13707_));
 sky130_fd_sc_hd__o21ai_4 _44254_ (.A1(_13434_),
    .A2(_13705_),
    .B1(_13371_),
    .Y(_13708_));
 sky130_fd_sc_hd__nand3_4 _44255_ (.A(_13708_),
    .B(_13703_),
    .C(_13702_),
    .Y(_13709_));
 sky130_fd_sc_hd__nand2_4 _44256_ (.A(_13707_),
    .B(_13709_),
    .Y(_13710_));
 sky130_vsdinv _44257_ (.A(_13411_),
    .Y(_13711_));
 sky130_fd_sc_hd__a21bo_4 _44258_ (.A1(_13413_),
    .A2(_13711_),
    .B1_N(_13414_),
    .X(_13712_));
 sky130_fd_sc_hd__nand2_4 _44259_ (.A(_12315_),
    .B(_08081_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand2_4 _44260_ (.A(_13448_),
    .B(_13713_),
    .Y(_13714_));
 sky130_fd_sc_hd__nand3_4 _44261_ (.A(_11686_),
    .B(_08259_),
    .C(_08257_),
    .Y(_13715_));
 sky130_fd_sc_hd__a21o_4 _44262_ (.A1(_13714_),
    .A2(_13715_),
    .B1(_13172_),
    .X(_13716_));
 sky130_fd_sc_hd__nand3_4 _44263_ (.A(_13714_),
    .B(_13172_),
    .C(_13715_),
    .Y(_13717_));
 sky130_fd_sc_hd__nand2_4 _44264_ (.A(_13716_),
    .B(_13717_),
    .Y(_13718_));
 sky130_vsdinv _44265_ (.A(_13718_),
    .Y(_13719_));
 sky130_fd_sc_hd__nand2_4 _44266_ (.A(_13712_),
    .B(_13719_),
    .Y(_13720_));
 sky130_fd_sc_hd__a21boi_4 _44267_ (.A1(_13413_),
    .A2(_13711_),
    .B1_N(_13414_),
    .Y(_13721_));
 sky130_fd_sc_hd__buf_1 _44268_ (.A(_13718_),
    .X(_13722_));
 sky130_fd_sc_hd__nand2_4 _44269_ (.A(_13721_),
    .B(_13722_),
    .Y(_13723_));
 sky130_fd_sc_hd__a21boi_4 _44270_ (.A1(_13449_),
    .A2(_13175_),
    .B1_N(_13450_),
    .Y(_13724_));
 sky130_vsdinv _44271_ (.A(_13724_),
    .Y(_13725_));
 sky130_fd_sc_hd__a21o_4 _44272_ (.A1(_13720_),
    .A2(_13723_),
    .B1(_13725_),
    .X(_13726_));
 sky130_fd_sc_hd__nand3_4 _44273_ (.A(_13720_),
    .B(_13725_),
    .C(_13723_),
    .Y(_13727_));
 sky130_fd_sc_hd__nand2_4 _44274_ (.A(_13726_),
    .B(_13727_),
    .Y(_13728_));
 sky130_fd_sc_hd__a21oi_4 _44275_ (.A1(_13416_),
    .A2(_13406_),
    .B1(_13408_),
    .Y(_13729_));
 sky130_fd_sc_hd__nand2_4 _44276_ (.A(_13728_),
    .B(_13729_),
    .Y(_13730_));
 sky130_fd_sc_hd__xor2_4 _44277_ (.A(_13711_),
    .B(_13415_),
    .X(_13731_));
 sky130_fd_sc_hd__o21ai_4 _44278_ (.A1(_13405_),
    .A2(_13731_),
    .B1(_13409_),
    .Y(_13732_));
 sky130_fd_sc_hd__nand3_4 _44279_ (.A(_13732_),
    .B(_13727_),
    .C(_13726_),
    .Y(_13733_));
 sky130_fd_sc_hd__nand2_4 _44280_ (.A(_13730_),
    .B(_13733_),
    .Y(_13734_));
 sky130_fd_sc_hd__a21oi_4 _44281_ (.A1(_13456_),
    .A2(_13458_),
    .B1(_13454_),
    .Y(_13735_));
 sky130_fd_sc_hd__nand2_4 _44282_ (.A(_13734_),
    .B(_13735_),
    .Y(_13736_));
 sky130_vsdinv _44283_ (.A(_13735_),
    .Y(_13737_));
 sky130_fd_sc_hd__nand3_4 _44284_ (.A(_13730_),
    .B(_13733_),
    .C(_13737_),
    .Y(_13738_));
 sky130_fd_sc_hd__nand2_4 _44285_ (.A(_13736_),
    .B(_13738_),
    .Y(_13739_));
 sky130_fd_sc_hd__a21boi_4 _44286_ (.A1(_13464_),
    .A2(_13468_),
    .B1_N(_13466_),
    .Y(_13740_));
 sky130_fd_sc_hd__nand2_4 _44287_ (.A(_13739_),
    .B(_13740_),
    .Y(_13741_));
 sky130_fd_sc_hd__nand2_4 _44288_ (.A(_13469_),
    .B(_13466_),
    .Y(_13742_));
 sky130_fd_sc_hd__nand3_4 _44289_ (.A(_13742_),
    .B(_13736_),
    .C(_13738_),
    .Y(_13743_));
 sky130_fd_sc_hd__nand2_4 _44290_ (.A(_13741_),
    .B(_13743_),
    .Y(_13744_));
 sky130_fd_sc_hd__buf_1 _44291_ (.A(_13479_),
    .X(_13745_));
 sky130_fd_sc_hd__nand2_4 _44292_ (.A(_13744_),
    .B(_13745_),
    .Y(_13746_));
 sky130_fd_sc_hd__buf_1 _44293_ (.A(_13482_),
    .X(_13747_));
 sky130_fd_sc_hd__nand3_4 _44294_ (.A(_13741_),
    .B(_13747_),
    .C(_13743_),
    .Y(_13748_));
 sky130_fd_sc_hd__nand2_4 _44295_ (.A(_13746_),
    .B(_13748_),
    .Y(_13749_));
 sky130_vsdinv _44296_ (.A(_13428_),
    .Y(_13750_));
 sky130_fd_sc_hd__a21oi_4 _44297_ (.A1(_13427_),
    .A2(_13432_),
    .B1(_13750_),
    .Y(_13751_));
 sky130_fd_sc_hd__nand2_4 _44298_ (.A(_13749_),
    .B(_13751_),
    .Y(_13752_));
 sky130_fd_sc_hd__a21o_4 _44299_ (.A1(_13427_),
    .A2(_13432_),
    .B1(_13750_),
    .X(_13753_));
 sky130_fd_sc_hd__nand3_4 _44300_ (.A(_13753_),
    .B(_13746_),
    .C(_13748_),
    .Y(_13754_));
 sky130_fd_sc_hd__buf_1 _44301_ (.A(_13754_),
    .X(_13755_));
 sky130_fd_sc_hd__buf_1 _44302_ (.A(_13482_),
    .X(_13756_));
 sky130_fd_sc_hd__a21boi_4 _44303_ (.A1(_13756_),
    .A2(_13474_),
    .B1_N(_13472_),
    .Y(_13757_));
 sky130_vsdinv _44304_ (.A(_13757_),
    .Y(_13758_));
 sky130_fd_sc_hd__a21o_4 _44305_ (.A1(_13752_),
    .A2(_13755_),
    .B1(_13758_),
    .X(_13759_));
 sky130_fd_sc_hd__nand3_4 _44306_ (.A(_13752_),
    .B(_13754_),
    .C(_13758_),
    .Y(_13760_));
 sky130_fd_sc_hd__nand2_4 _44307_ (.A(_13759_),
    .B(_13760_),
    .Y(_13761_));
 sky130_fd_sc_hd__nand2_4 _44308_ (.A(_13710_),
    .B(_13761_),
    .Y(_13762_));
 sky130_fd_sc_hd__a21oi_4 _44309_ (.A1(_13752_),
    .A2(_13755_),
    .B1(_13758_),
    .Y(_13763_));
 sky130_vsdinv _44310_ (.A(_13760_),
    .Y(_13764_));
 sky130_fd_sc_hd__nor2_4 _44311_ (.A(_13763_),
    .B(_13764_),
    .Y(_13765_));
 sky130_fd_sc_hd__nand3_4 _44312_ (.A(_13765_),
    .B(_13709_),
    .C(_13707_),
    .Y(_13766_));
 sky130_fd_sc_hd__nand2_4 _44313_ (.A(_13762_),
    .B(_13766_),
    .Y(_13767_));
 sky130_fd_sc_hd__a21boi_4 _44314_ (.A1(_13499_),
    .A2(_13439_),
    .B1_N(_13442_),
    .Y(_13768_));
 sky130_fd_sc_hd__nand2_4 _44315_ (.A(_13767_),
    .B(_13768_),
    .Y(_13769_));
 sky130_fd_sc_hd__a21oi_4 _44316_ (.A1(_13435_),
    .A2(_13436_),
    .B1(_13441_),
    .Y(_13770_));
 sky130_fd_sc_hd__o21ai_4 _44317_ (.A1(_13770_),
    .A2(_13495_),
    .B1(_13442_),
    .Y(_13771_));
 sky130_fd_sc_hd__nand3_4 _44318_ (.A(_13771_),
    .B(_13766_),
    .C(_13762_),
    .Y(_13772_));
 sky130_fd_sc_hd__nand2_4 _44319_ (.A(_13769_),
    .B(_13772_),
    .Y(_13773_));
 sky130_fd_sc_hd__a2bb2oi_4 _44320_ (.A1_N(_12920_),
    .A2_N(_13202_),
    .B1(_12658_),
    .B2(_13476_),
    .Y(_13774_));
 sky130_vsdinv _44321_ (.A(_13774_),
    .Y(_13775_));
 sky130_fd_sc_hd__buf_8 _44322_ (.A(_13775_),
    .X(_13776_));
 sky130_fd_sc_hd__a21boi_4 _44323_ (.A1(_13488_),
    .A2(_13492_),
    .B1_N(_13490_),
    .Y(_13777_));
 sky130_fd_sc_hd__xor2_4 _44324_ (.A(_13776_),
    .B(_13777_),
    .X(_13778_));
 sky130_fd_sc_hd__nand2_4 _44325_ (.A(_13773_),
    .B(_13778_),
    .Y(_13779_));
 sky130_vsdinv _44326_ (.A(_13778_),
    .Y(_13780_));
 sky130_fd_sc_hd__nand3_4 _44327_ (.A(_13769_),
    .B(_13772_),
    .C(_13780_),
    .Y(_13781_));
 sky130_fd_sc_hd__nand2_4 _44328_ (.A(_13779_),
    .B(_13781_),
    .Y(_13782_));
 sky130_fd_sc_hd__nand2_4 _44329_ (.A(_13534_),
    .B(_13782_),
    .Y(_13783_));
 sky130_fd_sc_hd__nand3_4 _44330_ (.A(_13533_),
    .B(_13779_),
    .C(_13781_),
    .Y(_13784_));
 sky130_fd_sc_hd__nand2_4 _44331_ (.A(_13783_),
    .B(_13784_),
    .Y(_13785_));
 sky130_fd_sc_hd__a21boi_4 _44332_ (.A1(_13225_),
    .A2(_13217_),
    .B1_N(_13508_),
    .Y(_13786_));
 sky130_vsdinv _44333_ (.A(_13786_),
    .Y(_13787_));
 sky130_fd_sc_hd__nand2_4 _44334_ (.A(_13785_),
    .B(_13787_),
    .Y(_13788_));
 sky130_fd_sc_hd__nand3_4 _44335_ (.A(_13783_),
    .B(_13786_),
    .C(_13784_),
    .Y(_13789_));
 sky130_fd_sc_hd__nand2_4 _44336_ (.A(_13788_),
    .B(_13789_),
    .Y(_13790_));
 sky130_fd_sc_hd__a21oi_4 _44337_ (.A1(_13511_),
    .A2(_13513_),
    .B1(_13517_),
    .Y(_13791_));
 sky130_fd_sc_hd__o21ai_4 _44338_ (.A1(_13521_),
    .A2(_13791_),
    .B1(_13518_),
    .Y(_13792_));
 sky130_vsdinv _44339_ (.A(_13792_),
    .Y(_13793_));
 sky130_fd_sc_hd__nand2_4 _44340_ (.A(_13790_),
    .B(_13793_),
    .Y(_13794_));
 sky130_fd_sc_hd__nand3_4 _44341_ (.A(_13792_),
    .B(_13788_),
    .C(_13789_),
    .Y(_13795_));
 sky130_fd_sc_hd__nand2_4 _44342_ (.A(_13794_),
    .B(_13795_),
    .Y(_13796_));
 sky130_fd_sc_hd__nand4_4 _44343_ (.A(_13260_),
    .B(_13259_),
    .C(_13526_),
    .D(_13528_),
    .Y(_13797_));
 sky130_fd_sc_hd__nor2_4 _44344_ (.A(_13262_),
    .B(_13797_),
    .Y(_13798_));
 sky130_fd_sc_hd__nand2_4 _44345_ (.A(_12685_),
    .B(_13798_),
    .Y(_13799_));
 sky130_fd_sc_hd__a21boi_4 _44346_ (.A1(_13530_),
    .A2(_13526_),
    .B1_N(_13528_),
    .Y(_13800_));
 sky130_fd_sc_hd__o21a_4 _44347_ (.A1(_13264_),
    .A2(_13797_),
    .B1(_13800_),
    .X(_13801_));
 sky130_fd_sc_hd__nand2_4 _44348_ (.A(_13799_),
    .B(_13801_),
    .Y(_13802_));
 sky130_fd_sc_hd__nand2_4 _44349_ (.A(_12682_),
    .B(_13798_),
    .Y(_13803_));
 sky130_fd_sc_hd__a21oi_4 _44350_ (.A1(_11424_),
    .A2(_11425_),
    .B1(_13803_),
    .Y(_13804_));
 sky130_fd_sc_hd__nor2_4 _44351_ (.A(_13802_),
    .B(_13804_),
    .Y(_13805_));
 sky130_fd_sc_hd__xor2_4 _44352_ (.A(_13796_),
    .B(_13805_),
    .X(_01445_));
 sky130_fd_sc_hd__a21boi_4 _44353_ (.A1(_13544_),
    .A2(_13557_),
    .B1_N(_13546_),
    .Y(_13806_));
 sky130_vsdinv _44354_ (.A(_13806_),
    .Y(_13807_));
 sky130_fd_sc_hd__buf_1 _44355_ (.A(_03632_),
    .X(_13808_));
 sky130_fd_sc_hd__nand2_4 _44356_ (.A(_06567_),
    .B(_12075_),
    .Y(_13809_));
 sky130_fd_sc_hd__o21ai_4 _44357_ (.A1(_08168_),
    .A2(_13808_),
    .B1(_13809_),
    .Y(_13810_));
 sky130_fd_sc_hd__nand4_4 _44358_ (.A(_03291_),
    .B(_07654_),
    .C(_11438_),
    .D(_11107_),
    .Y(_13811_));
 sky130_fd_sc_hd__nand2_4 _44359_ (.A(_06847_),
    .B(_10955_),
    .Y(_13812_));
 sky130_vsdinv _44360_ (.A(_13812_),
    .Y(_13813_));
 sky130_fd_sc_hd__a21o_4 _44361_ (.A1(_13810_),
    .A2(_13811_),
    .B1(_13813_),
    .X(_13814_));
 sky130_fd_sc_hd__nand3_4 _44362_ (.A(_13810_),
    .B(_13813_),
    .C(_13811_),
    .Y(_13815_));
 sky130_fd_sc_hd__nand2_4 _44363_ (.A(_13814_),
    .B(_13815_),
    .Y(_13816_));
 sky130_fd_sc_hd__a21boi_4 _44364_ (.A1(_13536_),
    .A2(_13541_),
    .B1_N(_13537_),
    .Y(_13817_));
 sky130_fd_sc_hd__nand2_4 _44365_ (.A(_13816_),
    .B(_13817_),
    .Y(_13818_));
 sky130_vsdinv _44366_ (.A(_13817_),
    .Y(_13819_));
 sky130_fd_sc_hd__nand3_4 _44367_ (.A(_13819_),
    .B(_13815_),
    .C(_13814_),
    .Y(_13820_));
 sky130_fd_sc_hd__nand2_4 _44368_ (.A(_06849_),
    .B(_11447_),
    .Y(_13821_));
 sky130_fd_sc_hd__nand2_4 _44369_ (.A(_07150_),
    .B(_11449_),
    .Y(_13822_));
 sky130_fd_sc_hd__nand2_4 _44370_ (.A(_13821_),
    .B(_13822_),
    .Y(_13823_));
 sky130_fd_sc_hd__nand4_4 _44371_ (.A(_07660_),
    .B(_07150_),
    .C(_10502_),
    .D(_10499_),
    .Y(_13824_));
 sky130_fd_sc_hd__buf_1 _44372_ (.A(_03313_),
    .X(_13825_));
 sky130_fd_sc_hd__nand2_4 _44373_ (.A(_13825_),
    .B(_03600_),
    .Y(_13826_));
 sky130_vsdinv _44374_ (.A(_13826_),
    .Y(_13827_));
 sky130_fd_sc_hd__a21o_4 _44375_ (.A1(_13823_),
    .A2(_13824_),
    .B1(_13827_),
    .X(_13828_));
 sky130_fd_sc_hd__nand3_4 _44376_ (.A(_13823_),
    .B(_13824_),
    .C(_13827_),
    .Y(_13829_));
 sky130_fd_sc_hd__and2_4 _44377_ (.A(_13828_),
    .B(_13829_),
    .X(_13830_));
 sky130_fd_sc_hd__nand3_4 _44378_ (.A(_13818_),
    .B(_13820_),
    .C(_13830_),
    .Y(_13831_));
 sky130_fd_sc_hd__nand2_4 _44379_ (.A(_13818_),
    .B(_13820_),
    .Y(_13832_));
 sky130_vsdinv _44380_ (.A(_13830_),
    .Y(_13833_));
 sky130_fd_sc_hd__nand2_4 _44381_ (.A(_13832_),
    .B(_13833_),
    .Y(_13834_));
 sky130_fd_sc_hd__nand3_4 _44382_ (.A(_13807_),
    .B(_13831_),
    .C(_13834_),
    .Y(_13835_));
 sky130_fd_sc_hd__nand2_4 _44383_ (.A(_13834_),
    .B(_13831_),
    .Y(_13836_));
 sky130_fd_sc_hd__nand2_4 _44384_ (.A(_13836_),
    .B(_13806_),
    .Y(_13837_));
 sky130_fd_sc_hd__nand2_4 _44385_ (.A(_13835_),
    .B(_13837_),
    .Y(_13838_));
 sky130_fd_sc_hd__nand2_4 _44386_ (.A(_11513_),
    .B(_12719_),
    .Y(_13839_));
 sky130_fd_sc_hd__nand2_4 _44387_ (.A(_12458_),
    .B(_12721_),
    .Y(_13840_));
 sky130_fd_sc_hd__nand2_4 _44388_ (.A(_13839_),
    .B(_13840_),
    .Y(_13841_));
 sky130_fd_sc_hd__buf_1 _44389_ (.A(_12427_),
    .X(_13842_));
 sky130_fd_sc_hd__nand4_4 _44390_ (.A(_11513_),
    .B(_07625_),
    .C(_13842_),
    .D(_03597_),
    .Y(_13843_));
 sky130_fd_sc_hd__nand2_4 _44391_ (.A(_07627_),
    .B(_03582_),
    .Y(_13844_));
 sky130_vsdinv _44392_ (.A(_13844_),
    .Y(_13845_));
 sky130_fd_sc_hd__a21o_4 _44393_ (.A1(_13841_),
    .A2(_13843_),
    .B1(_13845_),
    .X(_13846_));
 sky130_fd_sc_hd__nand3_4 _44394_ (.A(_13841_),
    .B(_13843_),
    .C(_13845_),
    .Y(_13847_));
 sky130_fd_sc_hd__maj3_4 _44395_ (.A(_13548_),
    .B(_13552_),
    .C(_13549_),
    .X(_13848_));
 sky130_fd_sc_hd__a21boi_4 _44396_ (.A1(_13846_),
    .A2(_13847_),
    .B1_N(_13848_),
    .Y(_13849_));
 sky130_vsdinv _44397_ (.A(_13849_),
    .Y(_13850_));
 sky130_vsdinv _44398_ (.A(_13848_),
    .Y(_13851_));
 sky130_fd_sc_hd__nand3_4 _44399_ (.A(_13851_),
    .B(_13846_),
    .C(_13847_),
    .Y(_13852_));
 sky130_fd_sc_hd__a21boi_4 _44400_ (.A1(_13567_),
    .A2(_13570_),
    .B1_N(_13568_),
    .Y(_13853_));
 sky130_vsdinv _44401_ (.A(_13853_),
    .Y(_13854_));
 sky130_fd_sc_hd__a21o_4 _44402_ (.A1(_13850_),
    .A2(_13852_),
    .B1(_13854_),
    .X(_13855_));
 sky130_fd_sc_hd__nand3_4 _44403_ (.A(_13850_),
    .B(_13854_),
    .C(_13852_),
    .Y(_13856_));
 sky130_fd_sc_hd__nand2_4 _44404_ (.A(_13855_),
    .B(_13856_),
    .Y(_13857_));
 sky130_fd_sc_hd__nand2_4 _44405_ (.A(_13838_),
    .B(_13857_),
    .Y(_13858_));
 sky130_fd_sc_hd__a21oi_4 _44406_ (.A1(_13850_),
    .A2(_13852_),
    .B1(_13854_),
    .Y(_13859_));
 sky130_vsdinv _44407_ (.A(_13856_),
    .Y(_13860_));
 sky130_fd_sc_hd__nor2_4 _44408_ (.A(_13859_),
    .B(_13860_),
    .Y(_13861_));
 sky130_fd_sc_hd__nand3_4 _44409_ (.A(_13861_),
    .B(_13835_),
    .C(_13837_),
    .Y(_13862_));
 sky130_fd_sc_hd__nand2_4 _44410_ (.A(_13858_),
    .B(_13862_),
    .Y(_13863_));
 sky130_fd_sc_hd__a21boi_4 _44411_ (.A1(_13561_),
    .A2(_13584_),
    .B1_N(_13563_),
    .Y(_13864_));
 sky130_fd_sc_hd__nand2_4 _44412_ (.A(_13863_),
    .B(_13864_),
    .Y(_13865_));
 sky130_vsdinv _44413_ (.A(_13864_),
    .Y(_13866_));
 sky130_fd_sc_hd__nand3_4 _44414_ (.A(_13866_),
    .B(_13862_),
    .C(_13858_),
    .Y(_13867_));
 sky130_fd_sc_hd__nand2_4 _44415_ (.A(_13865_),
    .B(_13867_),
    .Y(_13868_));
 sky130_fd_sc_hd__nand2_4 _44416_ (.A(_12192_),
    .B(_12466_),
    .Y(_13869_));
 sky130_fd_sc_hd__o21ai_4 _44417_ (.A1(_03338_),
    .A2(_03577_),
    .B1(_13869_),
    .Y(_13870_));
 sky130_fd_sc_hd__nand4_4 _44418_ (.A(_11871_),
    .B(_08307_),
    .C(_11172_),
    .D(_11173_),
    .Y(_13871_));
 sky130_fd_sc_hd__buf_1 _44419_ (.A(_10887_),
    .X(_13872_));
 sky130_fd_sc_hd__nand2_4 _44420_ (.A(_08526_),
    .B(_13872_),
    .Y(_13873_));
 sky130_vsdinv _44421_ (.A(_13873_),
    .Y(_13874_));
 sky130_fd_sc_hd__a21o_4 _44422_ (.A1(_13870_),
    .A2(_13871_),
    .B1(_13874_),
    .X(_13875_));
 sky130_fd_sc_hd__nand3_4 _44423_ (.A(_13870_),
    .B(_13874_),
    .C(_13871_),
    .Y(_13876_));
 sky130_fd_sc_hd__a21boi_4 _44424_ (.A1(_13596_),
    .A2(_13599_),
    .B1_N(_13597_),
    .Y(_13877_));
 sky130_vsdinv _44425_ (.A(_13877_),
    .Y(_13878_));
 sky130_fd_sc_hd__a21o_4 _44426_ (.A1(_13875_),
    .A2(_13876_),
    .B1(_13878_),
    .X(_13879_));
 sky130_fd_sc_hd__nand3_4 _44427_ (.A(_13875_),
    .B(_13878_),
    .C(_13876_),
    .Y(_13880_));
 sky130_fd_sc_hd__nand2_4 _44428_ (.A(_08760_),
    .B(_07980_),
    .Y(_13881_));
 sky130_fd_sc_hd__nand2_4 _44429_ (.A(_13088_),
    .B(_11186_),
    .Y(_13882_));
 sky130_fd_sc_hd__o21ai_4 _44430_ (.A1(_03355_),
    .A2(_03559_),
    .B1(_13882_),
    .Y(_13883_));
 sky130_fd_sc_hd__buf_1 _44431_ (.A(_07977_),
    .X(_13884_));
 sky130_fd_sc_hd__buf_1 _44432_ (.A(_11187_),
    .X(_13885_));
 sky130_fd_sc_hd__nand4_4 _44433_ (.A(_13610_),
    .B(_11915_),
    .C(_13884_),
    .D(_13885_),
    .Y(_13886_));
 sky130_fd_sc_hd__nand2_4 _44434_ (.A(_13883_),
    .B(_13886_),
    .Y(_13887_));
 sky130_fd_sc_hd__xor2_4 _44435_ (.A(_13881_),
    .B(_13887_),
    .X(_13888_));
 sky130_fd_sc_hd__a21o_4 _44436_ (.A1(_13879_),
    .A2(_13880_),
    .B1(_13888_),
    .X(_13889_));
 sky130_fd_sc_hd__nand3_4 _44437_ (.A(_13879_),
    .B(_13888_),
    .C(_13880_),
    .Y(_13890_));
 sky130_fd_sc_hd__a21boi_4 _44438_ (.A1(_13575_),
    .A2(_13579_),
    .B1_N(_13577_),
    .Y(_13891_));
 sky130_vsdinv _44439_ (.A(_13891_),
    .Y(_13892_));
 sky130_fd_sc_hd__a21oi_4 _44440_ (.A1(_13889_),
    .A2(_13890_),
    .B1(_13892_),
    .Y(_13893_));
 sky130_fd_sc_hd__nand3_4 _44441_ (.A(_13889_),
    .B(_13892_),
    .C(_13890_),
    .Y(_13894_));
 sky130_vsdinv _44442_ (.A(_13894_),
    .Y(_13895_));
 sky130_fd_sc_hd__a21oi_4 _44443_ (.A1(_13605_),
    .A2(_13614_),
    .B1(_13603_),
    .Y(_13896_));
 sky130_fd_sc_hd__o21ai_4 _44444_ (.A1(_13893_),
    .A2(_13895_),
    .B1(_13896_),
    .Y(_13897_));
 sky130_fd_sc_hd__a21o_4 _44445_ (.A1(_13889_),
    .A2(_13890_),
    .B1(_13892_),
    .X(_13898_));
 sky130_vsdinv _44446_ (.A(_13896_),
    .Y(_13899_));
 sky130_fd_sc_hd__nand3_4 _44447_ (.A(_13898_),
    .B(_13899_),
    .C(_13894_),
    .Y(_13900_));
 sky130_fd_sc_hd__nand2_4 _44448_ (.A(_13897_),
    .B(_13900_),
    .Y(_13901_));
 sky130_fd_sc_hd__nand2_4 _44449_ (.A(_13868_),
    .B(_13901_),
    .Y(_13902_));
 sky130_fd_sc_hd__a21oi_4 _44450_ (.A1(_13898_),
    .A2(_13894_),
    .B1(_13899_),
    .Y(_13903_));
 sky130_vsdinv _44451_ (.A(_13900_),
    .Y(_13904_));
 sky130_fd_sc_hd__nor2_4 _44452_ (.A(_13903_),
    .B(_13904_),
    .Y(_13905_));
 sky130_fd_sc_hd__nand3_4 _44453_ (.A(_13905_),
    .B(_13867_),
    .C(_13865_),
    .Y(_13906_));
 sky130_fd_sc_hd__nand2_4 _44454_ (.A(_13902_),
    .B(_13906_),
    .Y(_13907_));
 sky130_vsdinv _44455_ (.A(_13591_),
    .Y(_13908_));
 sky130_fd_sc_hd__a21oi_4 _44456_ (.A1(_13631_),
    .A2(_13589_),
    .B1(_13908_),
    .Y(_13909_));
 sky130_fd_sc_hd__nand2_4 _44457_ (.A(_13907_),
    .B(_13909_),
    .Y(_13910_));
 sky130_fd_sc_hd__a21o_4 _44458_ (.A1(_13631_),
    .A2(_13589_),
    .B1(_13908_),
    .X(_13911_));
 sky130_fd_sc_hd__nand3_4 _44459_ (.A(_13911_),
    .B(_13906_),
    .C(_13902_),
    .Y(_13912_));
 sky130_fd_sc_hd__nand2_4 _44460_ (.A(_13910_),
    .B(_13912_),
    .Y(_13913_));
 sky130_fd_sc_hd__a21boi_4 _44461_ (.A1(_13666_),
    .A2(_13669_),
    .B1_N(_13667_),
    .Y(_13914_));
 sky130_fd_sc_hd__nand2_4 _44462_ (.A(_10085_),
    .B(_11017_),
    .Y(_13915_));
 sky130_fd_sc_hd__nand2_4 _44463_ (.A(_13128_),
    .B(_11016_),
    .Y(_13916_));
 sky130_fd_sc_hd__nand2_4 _44464_ (.A(_13915_),
    .B(_13916_),
    .Y(_13917_));
 sky130_fd_sc_hd__nand4_4 _44465_ (.A(_11951_),
    .B(_13128_),
    .C(_03518_),
    .D(_12221_),
    .Y(_13918_));
 sky130_fd_sc_hd__nand2_4 _44466_ (.A(_11988_),
    .B(_08598_),
    .Y(_13919_));
 sky130_vsdinv _44467_ (.A(_13919_),
    .Y(_13920_));
 sky130_fd_sc_hd__a21o_4 _44468_ (.A1(_13917_),
    .A2(_13918_),
    .B1(_13920_),
    .X(_13921_));
 sky130_fd_sc_hd__nand3_4 _44469_ (.A(_13917_),
    .B(_13918_),
    .C(_13920_),
    .Y(_13922_));
 sky130_fd_sc_hd__nand2_4 _44470_ (.A(_13921_),
    .B(_13922_),
    .Y(_13923_));
 sky130_fd_sc_hd__nor2_4 _44471_ (.A(_13914_),
    .B(_13923_),
    .Y(_13924_));
 sky130_vsdinv _44472_ (.A(_13924_),
    .Y(_13925_));
 sky130_fd_sc_hd__nand2_4 _44473_ (.A(_12315_),
    .B(_07204_),
    .Y(_13926_));
 sky130_fd_sc_hd__nand2_4 _44474_ (.A(_10846_),
    .B(_07537_),
    .Y(_13927_));
 sky130_fd_sc_hd__nand2_4 _44475_ (.A(_12313_),
    .B(_06632_),
    .Y(_13928_));
 sky130_fd_sc_hd__nand2_4 _44476_ (.A(_13927_),
    .B(_13928_),
    .Y(_13929_));
 sky130_fd_sc_hd__nand4_4 _44477_ (.A(_11989_),
    .B(_11991_),
    .C(_07213_),
    .D(_07215_),
    .Y(_13930_));
 sky130_fd_sc_hd__nand2_4 _44478_ (.A(_13929_),
    .B(_13930_),
    .Y(_13931_));
 sky130_fd_sc_hd__xor2_4 _44479_ (.A(_13926_),
    .B(_13931_),
    .X(_13932_));
 sky130_fd_sc_hd__a21boi_4 _44480_ (.A1(_13921_),
    .A2(_13922_),
    .B1_N(_13914_),
    .Y(_13933_));
 sky130_vsdinv _44481_ (.A(_13933_),
    .Y(_13934_));
 sky130_fd_sc_hd__nand3_4 _44482_ (.A(_13925_),
    .B(_13932_),
    .C(_13934_),
    .Y(_13935_));
 sky130_vsdinv _44483_ (.A(_13935_),
    .Y(_13936_));
 sky130_fd_sc_hd__a21oi_4 _44484_ (.A1(_13925_),
    .A2(_13934_),
    .B1(_13932_),
    .Y(_13937_));
 sky130_fd_sc_hd__a21boi_4 _44485_ (.A1(_13654_),
    .A2(_13652_),
    .B1_N(_13651_),
    .Y(_13938_));
 sky130_vsdinv _44486_ (.A(_13938_),
    .Y(_13939_));
 sky130_fd_sc_hd__nand2_4 _44487_ (.A(_09577_),
    .B(_13644_),
    .Y(_13940_));
 sky130_fd_sc_hd__nand2_4 _44488_ (.A(_13112_),
    .B(_13643_),
    .Y(_13941_));
 sky130_fd_sc_hd__nand2_4 _44489_ (.A(_13940_),
    .B(_13941_),
    .Y(_13942_));
 sky130_fd_sc_hd__buf_1 _44490_ (.A(_10666_),
    .X(_13943_));
 sky130_fd_sc_hd__nand4_4 _44491_ (.A(_13943_),
    .B(_11893_),
    .C(_13089_),
    .D(_12190_),
    .Y(_13944_));
 sky130_fd_sc_hd__nand2_4 _44492_ (.A(_10084_),
    .B(_03531_),
    .Y(_13945_));
 sky130_vsdinv _44493_ (.A(_13945_),
    .Y(_13946_));
 sky130_fd_sc_hd__a21o_4 _44494_ (.A1(_13942_),
    .A2(_13944_),
    .B1(_13946_),
    .X(_13947_));
 sky130_fd_sc_hd__nand3_4 _44495_ (.A(_13942_),
    .B(_13944_),
    .C(_13946_),
    .Y(_13948_));
 sky130_vsdinv _44496_ (.A(_13606_),
    .Y(_13949_));
 sky130_fd_sc_hd__a21boi_4 _44497_ (.A1(_13609_),
    .A2(_13949_),
    .B1_N(_13612_),
    .Y(_13950_));
 sky130_fd_sc_hd__a21boi_4 _44498_ (.A1(_13947_),
    .A2(_13948_),
    .B1_N(_13950_),
    .Y(_13951_));
 sky130_fd_sc_hd__nand2_4 _44499_ (.A(_13947_),
    .B(_13948_),
    .Y(_13952_));
 sky130_fd_sc_hd__nor2_4 _44500_ (.A(_13950_),
    .B(_13952_),
    .Y(_13953_));
 sky130_fd_sc_hd__a21boi_4 _44501_ (.A1(_13642_),
    .A2(_13647_),
    .B1_N(_13645_),
    .Y(_13954_));
 sky130_fd_sc_hd__o21ai_4 _44502_ (.A1(_13951_),
    .A2(_13953_),
    .B1(_13954_),
    .Y(_13955_));
 sky130_fd_sc_hd__a211o_4 _44503_ (.A1(_13645_),
    .A2(_13649_),
    .B1(_13951_),
    .C1(_13953_),
    .X(_13956_));
 sky130_fd_sc_hd__nand3_4 _44504_ (.A(_13939_),
    .B(_13955_),
    .C(_13956_),
    .Y(_13957_));
 sky130_fd_sc_hd__nand2_4 _44505_ (.A(_13956_),
    .B(_13955_),
    .Y(_13958_));
 sky130_fd_sc_hd__nand2_4 _44506_ (.A(_13958_),
    .B(_13938_),
    .Y(_13959_));
 sky130_fd_sc_hd__nand2_4 _44507_ (.A(_13957_),
    .B(_13959_),
    .Y(_13960_));
 sky130_fd_sc_hd__o21ai_4 _44508_ (.A1(_13936_),
    .A2(_13937_),
    .B1(_13960_),
    .Y(_13961_));
 sky130_fd_sc_hd__nor2_4 _44509_ (.A(_13937_),
    .B(_13936_),
    .Y(_13962_));
 sky130_fd_sc_hd__nand3_4 _44510_ (.A(_13957_),
    .B(_13962_),
    .C(_13959_),
    .Y(_13963_));
 sky130_fd_sc_hd__a21boi_4 _44511_ (.A1(_13619_),
    .A2(_13624_),
    .B1_N(_13622_),
    .Y(_13964_));
 sky130_vsdinv _44512_ (.A(_13964_),
    .Y(_13965_));
 sky130_fd_sc_hd__a21oi_4 _44513_ (.A1(_13961_),
    .A2(_13963_),
    .B1(_13965_),
    .Y(_13966_));
 sky130_fd_sc_hd__nand3_4 _44514_ (.A(_13965_),
    .B(_13961_),
    .C(_13963_),
    .Y(_13967_));
 sky130_vsdinv _44515_ (.A(_13967_),
    .Y(_13968_));
 sky130_fd_sc_hd__a21boi_4 _44516_ (.A1(_13659_),
    .A2(_13687_),
    .B1_N(_13661_),
    .Y(_13969_));
 sky130_fd_sc_hd__o21ai_4 _44517_ (.A1(_13966_),
    .A2(_13968_),
    .B1(_13969_),
    .Y(_13970_));
 sky130_fd_sc_hd__a21o_4 _44518_ (.A1(_13961_),
    .A2(_13963_),
    .B1(_13965_),
    .X(_13971_));
 sky130_vsdinv _44519_ (.A(_13969_),
    .Y(_13972_));
 sky130_fd_sc_hd__nand3_4 _44520_ (.A(_13971_),
    .B(_13972_),
    .C(_13967_),
    .Y(_13973_));
 sky130_fd_sc_hd__nand2_4 _44521_ (.A(_13970_),
    .B(_13973_),
    .Y(_13974_));
 sky130_fd_sc_hd__nand2_4 _44522_ (.A(_13913_),
    .B(_13974_),
    .Y(_13975_));
 sky130_fd_sc_hd__nand4_4 _44523_ (.A(_13973_),
    .B(_13910_),
    .C(_13970_),
    .D(_13912_),
    .Y(_13976_));
 sky130_fd_sc_hd__nand2_4 _44524_ (.A(_13975_),
    .B(_13976_),
    .Y(_13977_));
 sky130_vsdinv _44525_ (.A(_13635_),
    .Y(_13978_));
 sky130_fd_sc_hd__o21a_4 _44526_ (.A1(_13701_),
    .A2(_13978_),
    .B1(_13638_),
    .X(_13979_));
 sky130_fd_sc_hd__nand2_4 _44527_ (.A(_13977_),
    .B(_13979_),
    .Y(_13980_));
 sky130_fd_sc_hd__o21ai_4 _44528_ (.A1(_13701_),
    .A2(_13978_),
    .B1(_13638_),
    .Y(_13981_));
 sky130_fd_sc_hd__nand3_4 _44529_ (.A(_13981_),
    .B(_13976_),
    .C(_13975_),
    .Y(_13982_));
 sky130_fd_sc_hd__nand2_4 _44530_ (.A(_13980_),
    .B(_13982_),
    .Y(_13983_));
 sky130_fd_sc_hd__nand2_4 _44531_ (.A(_13700_),
    .B(_13696_),
    .Y(_13984_));
 sky130_vsdinv _44532_ (.A(_13984_),
    .Y(_13985_));
 sky130_vsdinv _44533_ (.A(_13673_),
    .Y(_13986_));
 sky130_fd_sc_hd__o21a_4 _44534_ (.A1(_13674_),
    .A2(_13682_),
    .B1(_13986_),
    .X(_13987_));
 sky130_vsdinv _44535_ (.A(_13987_),
    .Y(_13988_));
 sky130_fd_sc_hd__maj3_4 _44536_ (.A(_13676_),
    .B(_13677_),
    .C(_13675_),
    .X(_13989_));
 sky130_vsdinv _44537_ (.A(_13989_),
    .Y(_13990_));
 sky130_fd_sc_hd__buf_1 _44538_ (.A(_13717_),
    .X(_13991_));
 sky130_fd_sc_hd__buf_1 _44539_ (.A(_13716_),
    .X(_13992_));
 sky130_fd_sc_hd__nand3_4 _44540_ (.A(_13990_),
    .B(_13991_),
    .C(_13992_),
    .Y(_13993_));
 sky130_fd_sc_hd__buf_1 _44541_ (.A(_13722_),
    .X(_13994_));
 sky130_fd_sc_hd__nand2_4 _44542_ (.A(_13994_),
    .B(_13989_),
    .Y(_13995_));
 sky130_fd_sc_hd__a21boi_4 _44543_ (.A1(_13714_),
    .A2(_13173_),
    .B1_N(_13715_),
    .Y(_13996_));
 sky130_vsdinv _44544_ (.A(_13996_),
    .Y(_13997_));
 sky130_fd_sc_hd__buf_1 _44545_ (.A(_13997_),
    .X(_13998_));
 sky130_fd_sc_hd__a21o_4 _44546_ (.A1(_13993_),
    .A2(_13995_),
    .B1(_13998_),
    .X(_13999_));
 sky130_fd_sc_hd__nand3_4 _44547_ (.A(_13993_),
    .B(_13998_),
    .C(_13995_),
    .Y(_14000_));
 sky130_fd_sc_hd__nand3_4 _44548_ (.A(_13988_),
    .B(_13999_),
    .C(_14000_),
    .Y(_14001_));
 sky130_fd_sc_hd__nand2_4 _44549_ (.A(_13999_),
    .B(_14000_),
    .Y(_14002_));
 sky130_fd_sc_hd__nand2_4 _44550_ (.A(_14002_),
    .B(_13987_),
    .Y(_14003_));
 sky130_fd_sc_hd__maj3_4 _44551_ (.A(_13724_),
    .B(_13721_),
    .C(_13994_),
    .X(_14004_));
 sky130_vsdinv _44552_ (.A(_14004_),
    .Y(_14005_));
 sky130_fd_sc_hd__a21o_4 _44553_ (.A1(_14001_),
    .A2(_14003_),
    .B1(_14005_),
    .X(_14006_));
 sky130_fd_sc_hd__nand3_4 _44554_ (.A(_14001_),
    .B(_14005_),
    .C(_14003_),
    .Y(_14007_));
 sky130_fd_sc_hd__nand2_4 _44555_ (.A(_14006_),
    .B(_14007_),
    .Y(_14008_));
 sky130_fd_sc_hd__a21boi_4 _44556_ (.A1(_13730_),
    .A2(_13737_),
    .B1_N(_13733_),
    .Y(_14009_));
 sky130_fd_sc_hd__nand2_4 _44557_ (.A(_14008_),
    .B(_14009_),
    .Y(_14010_));
 sky130_vsdinv _44558_ (.A(_14009_),
    .Y(_14011_));
 sky130_fd_sc_hd__nand3_4 _44559_ (.A(_14011_),
    .B(_14007_),
    .C(_14006_),
    .Y(_14012_));
 sky130_fd_sc_hd__nand2_4 _44560_ (.A(_14010_),
    .B(_14012_),
    .Y(_14013_));
 sky130_fd_sc_hd__nand2_4 _44561_ (.A(_14013_),
    .B(_13745_),
    .Y(_14014_));
 sky130_fd_sc_hd__buf_1 _44562_ (.A(_13478_),
    .X(_14015_));
 sky130_fd_sc_hd__nand3_4 _44563_ (.A(_14010_),
    .B(_14012_),
    .C(_14015_),
    .Y(_14016_));
 sky130_fd_sc_hd__nand2_4 _44564_ (.A(_14014_),
    .B(_14016_),
    .Y(_14017_));
 sky130_fd_sc_hd__nand2_4 _44565_ (.A(_13985_),
    .B(_14017_),
    .Y(_14018_));
 sky130_fd_sc_hd__nand3_4 _44566_ (.A(_13984_),
    .B(_14014_),
    .C(_14016_),
    .Y(_14019_));
 sky130_fd_sc_hd__buf_1 _44567_ (.A(_14019_),
    .X(_14020_));
 sky130_fd_sc_hd__nand2_4 _44568_ (.A(_14018_),
    .B(_14020_),
    .Y(_14021_));
 sky130_fd_sc_hd__a21boi_4 _44569_ (.A1(_13741_),
    .A2(_13756_),
    .B1_N(_13743_),
    .Y(_14022_));
 sky130_fd_sc_hd__nand2_4 _44570_ (.A(_14021_),
    .B(_14022_),
    .Y(_14023_));
 sky130_vsdinv _44571_ (.A(_14022_),
    .Y(_14024_));
 sky130_fd_sc_hd__nand3_4 _44572_ (.A(_14018_),
    .B(_14024_),
    .C(_14019_),
    .Y(_14025_));
 sky130_fd_sc_hd__nand2_4 _44573_ (.A(_14023_),
    .B(_14025_),
    .Y(_14026_));
 sky130_fd_sc_hd__nand2_4 _44574_ (.A(_13983_),
    .B(_14026_),
    .Y(_14027_));
 sky130_fd_sc_hd__a21oi_4 _44575_ (.A1(_14018_),
    .A2(_14020_),
    .B1(_14024_),
    .Y(_14028_));
 sky130_vsdinv _44576_ (.A(_14025_),
    .Y(_14029_));
 sky130_fd_sc_hd__nor2_4 _44577_ (.A(_14028_),
    .B(_14029_),
    .Y(_14030_));
 sky130_fd_sc_hd__nand3_4 _44578_ (.A(_14030_),
    .B(_13982_),
    .C(_13980_),
    .Y(_14031_));
 sky130_fd_sc_hd__nand2_4 _44579_ (.A(_14027_),
    .B(_14031_),
    .Y(_14032_));
 sky130_fd_sc_hd__a21boi_4 _44580_ (.A1(_13765_),
    .A2(_13707_),
    .B1_N(_13709_),
    .Y(_14033_));
 sky130_fd_sc_hd__nand2_4 _44581_ (.A(_14032_),
    .B(_14033_),
    .Y(_14034_));
 sky130_vsdinv _44582_ (.A(_13707_),
    .Y(_14035_));
 sky130_fd_sc_hd__o21ai_4 _44583_ (.A1(_13761_),
    .A2(_14035_),
    .B1(_13709_),
    .Y(_14036_));
 sky130_fd_sc_hd__nand3_4 _44584_ (.A(_14036_),
    .B(_14031_),
    .C(_14027_),
    .Y(_14037_));
 sky130_fd_sc_hd__nand2_4 _44585_ (.A(_14034_),
    .B(_14037_),
    .Y(_14038_));
 sky130_fd_sc_hd__a21boi_4 _44586_ (.A1(_13752_),
    .A2(_13758_),
    .B1_N(_13755_),
    .Y(_14039_));
 sky130_fd_sc_hd__xor2_4 _44587_ (.A(_13776_),
    .B(_14039_),
    .X(_14040_));
 sky130_fd_sc_hd__nand2_4 _44588_ (.A(_14038_),
    .B(_14040_),
    .Y(_14041_));
 sky130_vsdinv _44589_ (.A(_14040_),
    .Y(_14042_));
 sky130_fd_sc_hd__nand3_4 _44590_ (.A(_14034_),
    .B(_14037_),
    .C(_14042_),
    .Y(_14043_));
 sky130_fd_sc_hd__nand2_4 _44591_ (.A(_14041_),
    .B(_14043_),
    .Y(_14044_));
 sky130_fd_sc_hd__a21boi_4 _44592_ (.A1(_13769_),
    .A2(_13780_),
    .B1_N(_13772_),
    .Y(_14045_));
 sky130_fd_sc_hd__nand2_4 _44593_ (.A(_14044_),
    .B(_14045_),
    .Y(_14046_));
 sky130_fd_sc_hd__nand2_4 _44594_ (.A(_13781_),
    .B(_13772_),
    .Y(_14047_));
 sky130_fd_sc_hd__nand3_4 _44595_ (.A(_14047_),
    .B(_14041_),
    .C(_14043_),
    .Y(_14048_));
 sky130_fd_sc_hd__nand2_4 _44596_ (.A(_14046_),
    .B(_14048_),
    .Y(_14049_));
 sky130_fd_sc_hd__buf_1 _44597_ (.A(_13774_),
    .X(_14050_));
 sky130_fd_sc_hd__a21oi_4 _44598_ (.A1(_13494_),
    .A2(_13490_),
    .B1(_14050_),
    .Y(_14051_));
 sky130_vsdinv _44599_ (.A(_14051_),
    .Y(_14052_));
 sky130_fd_sc_hd__nand2_4 _44600_ (.A(_14049_),
    .B(_14052_),
    .Y(_14053_));
 sky130_fd_sc_hd__nand3_4 _44601_ (.A(_14046_),
    .B(_14051_),
    .C(_14048_),
    .Y(_14054_));
 sky130_fd_sc_hd__a21oi_4 _44602_ (.A1(_13779_),
    .A2(_13781_),
    .B1(_13533_),
    .Y(_14055_));
 sky130_fd_sc_hd__o21ai_4 _44603_ (.A1(_13787_),
    .A2(_14055_),
    .B1(_13784_),
    .Y(_14056_));
 sky130_fd_sc_hd__a21o_4 _44604_ (.A1(_14053_),
    .A2(_14054_),
    .B1(_14056_),
    .X(_14057_));
 sky130_fd_sc_hd__nand3_4 _44605_ (.A(_14053_),
    .B(_14056_),
    .C(_14054_),
    .Y(_14058_));
 sky130_fd_sc_hd__nand2_4 _44606_ (.A(_14057_),
    .B(_14058_),
    .Y(_14059_));
 sky130_fd_sc_hd__o21ai_4 _44607_ (.A1(_13796_),
    .A2(_13805_),
    .B1(_13795_),
    .Y(_14060_));
 sky130_fd_sc_hd__xnor2_4 _44608_ (.A(_14059_),
    .B(_14060_),
    .Y(_01446_));
 sky130_fd_sc_hd__a21boi_4 _44609_ (.A1(_13810_),
    .A2(_13813_),
    .B1_N(_13811_),
    .Y(_14061_));
 sky130_vsdinv _44610_ (.A(_14061_),
    .Y(_14062_));
 sky130_fd_sc_hd__nand2_4 _44611_ (.A(_08607_),
    .B(_11102_),
    .Y(_14063_));
 sky130_fd_sc_hd__o21ai_4 _44612_ (.A1(_08394_),
    .A2(_03633_),
    .B1(_14063_),
    .Y(_14064_));
 sky130_fd_sc_hd__nand2_4 _44613_ (.A(_03303_),
    .B(_11762_),
    .Y(_14065_));
 sky130_vsdinv _44614_ (.A(_14065_),
    .Y(_14066_));
 sky130_fd_sc_hd__nand4_4 _44615_ (.A(_03295_),
    .B(_07822_),
    .C(_11105_),
    .D(_12076_),
    .Y(_14067_));
 sky130_fd_sc_hd__nand3_4 _44616_ (.A(_14064_),
    .B(_14066_),
    .C(_14067_),
    .Y(_14068_));
 sky130_fd_sc_hd__nand2_4 _44617_ (.A(_14064_),
    .B(_14067_),
    .Y(_14069_));
 sky130_fd_sc_hd__nand2_4 _44618_ (.A(_14069_),
    .B(_14065_),
    .Y(_14070_));
 sky130_fd_sc_hd__nand3_4 _44619_ (.A(_14062_),
    .B(_14068_),
    .C(_14070_),
    .Y(_14071_));
 sky130_fd_sc_hd__nand2_4 _44620_ (.A(_14070_),
    .B(_14068_),
    .Y(_14072_));
 sky130_fd_sc_hd__nand2_4 _44621_ (.A(_14072_),
    .B(_14061_),
    .Y(_14073_));
 sky130_fd_sc_hd__nand2_4 _44622_ (.A(_14071_),
    .B(_14073_),
    .Y(_14074_));
 sky130_fd_sc_hd__nand2_4 _44623_ (.A(_06999_),
    .B(_11119_),
    .Y(_14075_));
 sky130_fd_sc_hd__nand2_4 _44624_ (.A(_07152_),
    .B(_11121_),
    .Y(_14076_));
 sky130_fd_sc_hd__nand2_4 _44625_ (.A(_14075_),
    .B(_14076_),
    .Y(_14077_));
 sky130_fd_sc_hd__nand4_4 _44626_ (.A(_10584_),
    .B(_06992_),
    .C(_11776_),
    .D(_10499_),
    .Y(_14078_));
 sky130_fd_sc_hd__nand2_4 _44627_ (.A(_10198_),
    .B(_03600_),
    .Y(_14079_));
 sky130_vsdinv _44628_ (.A(_14079_),
    .Y(_14080_));
 sky130_fd_sc_hd__a21o_4 _44629_ (.A1(_14077_),
    .A2(_14078_),
    .B1(_14080_),
    .X(_14081_));
 sky130_fd_sc_hd__nand3_4 _44630_ (.A(_14077_),
    .B(_14078_),
    .C(_14080_),
    .Y(_14082_));
 sky130_fd_sc_hd__nand2_4 _44631_ (.A(_14081_),
    .B(_14082_),
    .Y(_14083_));
 sky130_fd_sc_hd__nand2_4 _44632_ (.A(_14074_),
    .B(_14083_),
    .Y(_14084_));
 sky130_vsdinv _44633_ (.A(_14083_),
    .Y(_14085_));
 sky130_fd_sc_hd__nand3_4 _44634_ (.A(_14071_),
    .B(_14073_),
    .C(_14085_),
    .Y(_14086_));
 sky130_fd_sc_hd__nand2_4 _44635_ (.A(_14084_),
    .B(_14086_),
    .Y(_14087_));
 sky130_fd_sc_hd__a21boi_4 _44636_ (.A1(_13818_),
    .A2(_13830_),
    .B1_N(_13820_),
    .Y(_14088_));
 sky130_fd_sc_hd__nand2_4 _44637_ (.A(_14087_),
    .B(_14088_),
    .Y(_14089_));
 sky130_fd_sc_hd__nand2_4 _44638_ (.A(_13831_),
    .B(_13820_),
    .Y(_14090_));
 sky130_fd_sc_hd__nand3_4 _44639_ (.A(_14090_),
    .B(_14086_),
    .C(_14084_),
    .Y(_14091_));
 sky130_fd_sc_hd__nand2_4 _44640_ (.A(_14089_),
    .B(_14091_),
    .Y(_14092_));
 sky130_fd_sc_hd__nand2_4 _44641_ (.A(_03325_),
    .B(_03596_),
    .Y(_14093_));
 sky130_fd_sc_hd__nand2_4 _44642_ (.A(_11010_),
    .B(_13011_),
    .Y(_14094_));
 sky130_fd_sc_hd__nand2_4 _44643_ (.A(_14093_),
    .B(_14094_),
    .Y(_14095_));
 sky130_fd_sc_hd__buf_1 _44644_ (.A(_09038_),
    .X(_14096_));
 sky130_fd_sc_hd__nand4_4 _44645_ (.A(_11556_),
    .B(_14096_),
    .C(_11797_),
    .D(_12431_),
    .Y(_14097_));
 sky130_fd_sc_hd__nand2_4 _44646_ (.A(_11559_),
    .B(_09347_),
    .Y(_14098_));
 sky130_vsdinv _44647_ (.A(_14098_),
    .Y(_14099_));
 sky130_fd_sc_hd__a21o_4 _44648_ (.A1(_14095_),
    .A2(_14097_),
    .B1(_14099_),
    .X(_14100_));
 sky130_fd_sc_hd__nand3_4 _44649_ (.A(_14095_),
    .B(_14097_),
    .C(_14099_),
    .Y(_14101_));
 sky130_fd_sc_hd__nand2_4 _44650_ (.A(_14100_),
    .B(_14101_),
    .Y(_14102_));
 sky130_fd_sc_hd__a21boi_4 _44651_ (.A1(_13823_),
    .A2(_13827_),
    .B1_N(_13824_),
    .Y(_14103_));
 sky130_fd_sc_hd__nand2_4 _44652_ (.A(_14102_),
    .B(_14103_),
    .Y(_14104_));
 sky130_vsdinv _44653_ (.A(_14103_),
    .Y(_14105_));
 sky130_fd_sc_hd__nand3_4 _44654_ (.A(_14105_),
    .B(_14100_),
    .C(_14101_),
    .Y(_14106_));
 sky130_fd_sc_hd__a21boi_4 _44655_ (.A1(_13841_),
    .A2(_13845_),
    .B1_N(_13843_),
    .Y(_14107_));
 sky130_vsdinv _44656_ (.A(_14107_),
    .Y(_14108_));
 sky130_fd_sc_hd__a21o_4 _44657_ (.A1(_14104_),
    .A2(_14106_),
    .B1(_14108_),
    .X(_14109_));
 sky130_fd_sc_hd__nand3_4 _44658_ (.A(_14104_),
    .B(_14106_),
    .C(_14108_),
    .Y(_14110_));
 sky130_fd_sc_hd__nand2_4 _44659_ (.A(_14109_),
    .B(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__nand2_4 _44660_ (.A(_14092_),
    .B(_14111_),
    .Y(_14112_));
 sky130_vsdinv _44661_ (.A(_14111_),
    .Y(_14113_));
 sky130_fd_sc_hd__nand3_4 _44662_ (.A(_14089_),
    .B(_14091_),
    .C(_14113_),
    .Y(_14114_));
 sky130_fd_sc_hd__nand2_4 _44663_ (.A(_14112_),
    .B(_14114_),
    .Y(_14115_));
 sky130_fd_sc_hd__a21boi_4 _44664_ (.A1(_13861_),
    .A2(_13837_),
    .B1_N(_13835_),
    .Y(_14116_));
 sky130_fd_sc_hd__nand2_4 _44665_ (.A(_14115_),
    .B(_14116_),
    .Y(_14117_));
 sky130_fd_sc_hd__a21boi_4 _44666_ (.A1(_13834_),
    .A2(_13831_),
    .B1_N(_13806_),
    .Y(_14118_));
 sky130_fd_sc_hd__o21ai_4 _44667_ (.A1(_13857_),
    .A2(_14118_),
    .B1(_13835_),
    .Y(_14119_));
 sky130_fd_sc_hd__nand3_4 _44668_ (.A(_14119_),
    .B(_14114_),
    .C(_14112_),
    .Y(_14120_));
 sky130_fd_sc_hd__nand2_4 _44669_ (.A(_14117_),
    .B(_14120_),
    .Y(_14121_));
 sky130_fd_sc_hd__nand2_4 _44670_ (.A(_13340_),
    .B(_11167_),
    .Y(_14122_));
 sky130_fd_sc_hd__nand2_4 _44671_ (.A(_08523_),
    .B(_11169_),
    .Y(_14123_));
 sky130_fd_sc_hd__nand2_4 _44672_ (.A(_14122_),
    .B(_14123_),
    .Y(_14124_));
 sky130_fd_sc_hd__nand4_4 _44673_ (.A(_13340_),
    .B(_10625_),
    .C(_12156_),
    .D(_11167_),
    .Y(_14125_));
 sky130_fd_sc_hd__nand2_4 _44674_ (.A(_08315_),
    .B(_10540_),
    .Y(_14126_));
 sky130_vsdinv _44675_ (.A(_14126_),
    .Y(_14127_));
 sky130_fd_sc_hd__a21o_4 _44676_ (.A1(_14124_),
    .A2(_14125_),
    .B1(_14127_),
    .X(_14128_));
 sky130_fd_sc_hd__nand3_4 _44677_ (.A(_14124_),
    .B(_14125_),
    .C(_14127_),
    .Y(_14129_));
 sky130_fd_sc_hd__a21boi_4 _44678_ (.A1(_13870_),
    .A2(_13874_),
    .B1_N(_13871_),
    .Y(_14130_));
 sky130_vsdinv _44679_ (.A(_14130_),
    .Y(_14131_));
 sky130_fd_sc_hd__a21o_4 _44680_ (.A1(_14128_),
    .A2(_14129_),
    .B1(_14131_),
    .X(_14132_));
 sky130_fd_sc_hd__nand3_4 _44681_ (.A(_14131_),
    .B(_14128_),
    .C(_14129_),
    .Y(_14133_));
 sky130_fd_sc_hd__nand2_4 _44682_ (.A(_14132_),
    .B(_14133_),
    .Y(_14134_));
 sky130_fd_sc_hd__nand2_4 _44683_ (.A(_10789_),
    .B(_07980_),
    .Y(_14135_));
 sky130_fd_sc_hd__nand2_4 _44684_ (.A(_11912_),
    .B(_11516_),
    .Y(_14136_));
 sky130_fd_sc_hd__buf_1 _44685_ (.A(_11249_),
    .X(_14137_));
 sky130_fd_sc_hd__nand2_4 _44686_ (.A(_14137_),
    .B(_11186_),
    .Y(_14138_));
 sky130_fd_sc_hd__nand2_4 _44687_ (.A(_14136_),
    .B(_14138_),
    .Y(_14139_));
 sky130_fd_sc_hd__buf_1 _44688_ (.A(_03358_),
    .X(_14140_));
 sky130_fd_sc_hd__nand4_4 _44689_ (.A(_14140_),
    .B(_12226_),
    .C(_13611_),
    .D(_11523_),
    .Y(_14141_));
 sky130_fd_sc_hd__nand2_4 _44690_ (.A(_14139_),
    .B(_14141_),
    .Y(_14142_));
 sky130_fd_sc_hd__xor2_4 _44691_ (.A(_14135_),
    .B(_14142_),
    .X(_14143_));
 sky130_vsdinv _44692_ (.A(_14143_),
    .Y(_14144_));
 sky130_fd_sc_hd__nand2_4 _44693_ (.A(_14134_),
    .B(_14144_),
    .Y(_14145_));
 sky130_fd_sc_hd__nand3_4 _44694_ (.A(_14132_),
    .B(_14143_),
    .C(_14133_),
    .Y(_14146_));
 sky130_fd_sc_hd__o21ai_4 _44695_ (.A1(_13853_),
    .A2(_13849_),
    .B1(_13852_),
    .Y(_14147_));
 sky130_fd_sc_hd__a21oi_4 _44696_ (.A1(_14145_),
    .A2(_14146_),
    .B1(_14147_),
    .Y(_14148_));
 sky130_fd_sc_hd__nand3_4 _44697_ (.A(_14145_),
    .B(_14147_),
    .C(_14146_),
    .Y(_14149_));
 sky130_vsdinv _44698_ (.A(_14149_),
    .Y(_14150_));
 sky130_vsdinv _44699_ (.A(_13880_),
    .Y(_14151_));
 sky130_fd_sc_hd__a21oi_4 _44700_ (.A1(_13879_),
    .A2(_13888_),
    .B1(_14151_),
    .Y(_14152_));
 sky130_fd_sc_hd__o21ai_4 _44701_ (.A1(_14148_),
    .A2(_14150_),
    .B1(_14152_),
    .Y(_14153_));
 sky130_vsdinv _44702_ (.A(_14148_),
    .Y(_14154_));
 sky130_vsdinv _44703_ (.A(_14152_),
    .Y(_14155_));
 sky130_fd_sc_hd__nand3_4 _44704_ (.A(_14154_),
    .B(_14155_),
    .C(_14149_),
    .Y(_14156_));
 sky130_fd_sc_hd__nand2_4 _44705_ (.A(_14153_),
    .B(_14156_),
    .Y(_14157_));
 sky130_fd_sc_hd__nand2_4 _44706_ (.A(_14121_),
    .B(_14157_),
    .Y(_14158_));
 sky130_fd_sc_hd__nand4_4 _44707_ (.A(_14156_),
    .B(_14117_),
    .C(_14120_),
    .D(_14153_),
    .Y(_14159_));
 sky130_fd_sc_hd__nand2_4 _44708_ (.A(_14158_),
    .B(_14159_),
    .Y(_14160_));
 sky130_fd_sc_hd__a21boi_4 _44709_ (.A1(_13858_),
    .A2(_13862_),
    .B1_N(_13864_),
    .Y(_14161_));
 sky130_fd_sc_hd__o21a_4 _44710_ (.A1(_13901_),
    .A2(_14161_),
    .B1(_13867_),
    .X(_14162_));
 sky130_fd_sc_hd__nand2_4 _44711_ (.A(_14160_),
    .B(_14162_),
    .Y(_14163_));
 sky130_fd_sc_hd__o21ai_4 _44712_ (.A1(_13901_),
    .A2(_14161_),
    .B1(_13867_),
    .Y(_14164_));
 sky130_fd_sc_hd__nand3_4 _44713_ (.A(_14164_),
    .B(_14159_),
    .C(_14158_),
    .Y(_14165_));
 sky130_fd_sc_hd__nand2_4 _44714_ (.A(_14163_),
    .B(_14165_),
    .Y(_14166_));
 sky130_fd_sc_hd__nand2_4 _44715_ (.A(_13087_),
    .B(_13055_),
    .Y(_14167_));
 sky130_fd_sc_hd__maj3_4 _44716_ (.A(_14167_),
    .B(_13882_),
    .C(_13881_),
    .X(_14168_));
 sky130_fd_sc_hd__nand2_4 _44717_ (.A(_11635_),
    .B(_07717_),
    .Y(_14169_));
 sky130_fd_sc_hd__nand2_4 _44718_ (.A(_09580_),
    .B(_03536_),
    .Y(_14170_));
 sky130_fd_sc_hd__nand2_4 _44719_ (.A(_14169_),
    .B(_14170_),
    .Y(_14171_));
 sky130_fd_sc_hd__nand4_4 _44720_ (.A(_13112_),
    .B(_11639_),
    .C(_13643_),
    .D(_13644_),
    .Y(_14172_));
 sky130_fd_sc_hd__nand2_4 _44721_ (.A(_10822_),
    .B(_07720_),
    .Y(_14173_));
 sky130_vsdinv _44722_ (.A(_14173_),
    .Y(_14174_));
 sky130_fd_sc_hd__a21o_4 _44723_ (.A1(_14171_),
    .A2(_14172_),
    .B1(_14174_),
    .X(_14175_));
 sky130_fd_sc_hd__nand3_4 _44724_ (.A(_14171_),
    .B(_14172_),
    .C(_14174_),
    .Y(_14176_));
 sky130_fd_sc_hd__nand2_4 _44725_ (.A(_14175_),
    .B(_14176_),
    .Y(_14177_));
 sky130_fd_sc_hd__or2_4 _44726_ (.A(_14168_),
    .B(_14177_),
    .X(_14178_));
 sky130_fd_sc_hd__nand2_4 _44727_ (.A(_14177_),
    .B(_14168_),
    .Y(_14179_));
 sky130_fd_sc_hd__a21boi_4 _44728_ (.A1(_13942_),
    .A2(_13946_),
    .B1_N(_13944_),
    .Y(_14180_));
 sky130_vsdinv _44729_ (.A(_14180_),
    .Y(_14181_));
 sky130_fd_sc_hd__a21o_4 _44730_ (.A1(_14178_),
    .A2(_14179_),
    .B1(_14181_),
    .X(_14182_));
 sky130_fd_sc_hd__nand3_4 _44731_ (.A(_14178_),
    .B(_14181_),
    .C(_14179_),
    .Y(_14183_));
 sky130_fd_sc_hd__nand2_4 _44732_ (.A(_14182_),
    .B(_14183_),
    .Y(_14184_));
 sky130_fd_sc_hd__maj3_4 _44733_ (.A(_13950_),
    .B(_13952_),
    .C(_13954_),
    .X(_14185_));
 sky130_fd_sc_hd__nand2_4 _44734_ (.A(_14184_),
    .B(_14185_),
    .Y(_14186_));
 sky130_vsdinv _44735_ (.A(_14185_),
    .Y(_14187_));
 sky130_fd_sc_hd__nand3_4 _44736_ (.A(_14182_),
    .B(_14187_),
    .C(_14183_),
    .Y(_14188_));
 sky130_fd_sc_hd__nand2_4 _44737_ (.A(_14186_),
    .B(_14188_),
    .Y(_14189_));
 sky130_fd_sc_hd__a21boi_4 _44738_ (.A1(_13917_),
    .A2(_13920_),
    .B1_N(_13918_),
    .Y(_14190_));
 sky130_fd_sc_hd__nand2_4 _44739_ (.A(_12278_),
    .B(_07187_),
    .Y(_14191_));
 sky130_fd_sc_hd__nand2_4 _44740_ (.A(_12878_),
    .B(_07189_),
    .Y(_14192_));
 sky130_fd_sc_hd__nand2_4 _44741_ (.A(_14191_),
    .B(_14192_),
    .Y(_14193_));
 sky130_fd_sc_hd__nand4_4 _44742_ (.A(_13124_),
    .B(_11323_),
    .C(_07522_),
    .D(_07194_),
    .Y(_14194_));
 sky130_fd_sc_hd__nand2_4 _44743_ (.A(_12308_),
    .B(_07197_),
    .Y(_14195_));
 sky130_vsdinv _44744_ (.A(_14195_),
    .Y(_14196_));
 sky130_fd_sc_hd__a21o_4 _44745_ (.A1(_14193_),
    .A2(_14194_),
    .B1(_14196_),
    .X(_14197_));
 sky130_fd_sc_hd__nand3_4 _44746_ (.A(_14193_),
    .B(_14194_),
    .C(_14196_),
    .Y(_14198_));
 sky130_fd_sc_hd__nand2_4 _44747_ (.A(_14197_),
    .B(_14198_),
    .Y(_14199_));
 sky130_fd_sc_hd__nor2_4 _44748_ (.A(_14190_),
    .B(_14199_),
    .Y(_14200_));
 sky130_vsdinv _44749_ (.A(_14200_),
    .Y(_14201_));
 sky130_fd_sc_hd__a21boi_4 _44750_ (.A1(_14197_),
    .A2(_14198_),
    .B1_N(_14190_),
    .Y(_14202_));
 sky130_vsdinv _44751_ (.A(_14202_),
    .Y(_14203_));
 sky130_fd_sc_hd__buf_1 _44752_ (.A(_12310_),
    .X(_14204_));
 sky130_fd_sc_hd__nand2_4 _44753_ (.A(_14204_),
    .B(_07669_),
    .Y(_14205_));
 sky130_fd_sc_hd__nand2_4 _44754_ (.A(_12907_),
    .B(_06892_),
    .Y(_14206_));
 sky130_fd_sc_hd__nand2_4 _44755_ (.A(_14205_),
    .B(_14206_),
    .Y(_14207_));
 sky130_fd_sc_hd__nand4_4 _44756_ (.A(_14204_),
    .B(_12907_),
    .C(_06892_),
    .D(_07669_),
    .Y(_14208_));
 sky130_fd_sc_hd__nand2_4 _44757_ (.A(_14207_),
    .B(_14208_),
    .Y(_14209_));
 sky130_fd_sc_hd__xor2_4 _44758_ (.A(_13926_),
    .B(_14209_),
    .X(_14210_));
 sky130_fd_sc_hd__a21oi_4 _44759_ (.A1(_14201_),
    .A2(_14203_),
    .B1(_14210_),
    .Y(_14211_));
 sky130_fd_sc_hd__nand3_4 _44760_ (.A(_14201_),
    .B(_14210_),
    .C(_14203_),
    .Y(_14212_));
 sky130_vsdinv _44761_ (.A(_14212_),
    .Y(_14213_));
 sky130_fd_sc_hd__nor2_4 _44762_ (.A(_14211_),
    .B(_14213_),
    .Y(_14214_));
 sky130_vsdinv _44763_ (.A(_14214_),
    .Y(_14215_));
 sky130_fd_sc_hd__nand2_4 _44764_ (.A(_14189_),
    .B(_14215_),
    .Y(_14216_));
 sky130_fd_sc_hd__nand3_4 _44765_ (.A(_14186_),
    .B(_14214_),
    .C(_14188_),
    .Y(_14217_));
 sky130_fd_sc_hd__nand2_4 _44766_ (.A(_14216_),
    .B(_14217_),
    .Y(_14218_));
 sky130_fd_sc_hd__o21ai_4 _44767_ (.A1(_13896_),
    .A2(_13893_),
    .B1(_13894_),
    .Y(_14219_));
 sky130_vsdinv _44768_ (.A(_14219_),
    .Y(_14220_));
 sky130_fd_sc_hd__nand2_4 _44769_ (.A(_14218_),
    .B(_14220_),
    .Y(_14221_));
 sky130_fd_sc_hd__nand3_4 _44770_ (.A(_14216_),
    .B(_14219_),
    .C(_14217_),
    .Y(_14222_));
 sky130_fd_sc_hd__buf_1 _44771_ (.A(_14222_),
    .X(_14223_));
 sky130_fd_sc_hd__a21boi_4 _44772_ (.A1(_13962_),
    .A2(_13959_),
    .B1_N(_13957_),
    .Y(_14224_));
 sky130_vsdinv _44773_ (.A(_14224_),
    .Y(_14225_));
 sky130_fd_sc_hd__a21o_4 _44774_ (.A1(_14221_),
    .A2(_14223_),
    .B1(_14225_),
    .X(_14226_));
 sky130_fd_sc_hd__nand3_4 _44775_ (.A(_14221_),
    .B(_14225_),
    .C(_14222_),
    .Y(_14227_));
 sky130_fd_sc_hd__nand2_4 _44776_ (.A(_14226_),
    .B(_14227_),
    .Y(_14228_));
 sky130_fd_sc_hd__nand2_4 _44777_ (.A(_14166_),
    .B(_14228_),
    .Y(_14229_));
 sky130_fd_sc_hd__a21oi_4 _44778_ (.A1(_14221_),
    .A2(_14223_),
    .B1(_14225_),
    .Y(_14230_));
 sky130_vsdinv _44779_ (.A(_14227_),
    .Y(_14231_));
 sky130_fd_sc_hd__nor2_4 _44780_ (.A(_14230_),
    .B(_14231_),
    .Y(_14232_));
 sky130_fd_sc_hd__nand3_4 _44781_ (.A(_14232_),
    .B(_14165_),
    .C(_14163_),
    .Y(_14233_));
 sky130_fd_sc_hd__nand2_4 _44782_ (.A(_14229_),
    .B(_14233_),
    .Y(_14234_));
 sky130_fd_sc_hd__a21oi_4 _44783_ (.A1(_13902_),
    .A2(_13906_),
    .B1(_13911_),
    .Y(_14235_));
 sky130_fd_sc_hd__o21a_4 _44784_ (.A1(_14235_),
    .A2(_13974_),
    .B1(_13912_),
    .X(_14236_));
 sky130_fd_sc_hd__nand2_4 _44785_ (.A(_14234_),
    .B(_14236_),
    .Y(_14237_));
 sky130_fd_sc_hd__o21ai_4 _44786_ (.A1(_14235_),
    .A2(_13974_),
    .B1(_13912_),
    .Y(_14238_));
 sky130_fd_sc_hd__nand3_4 _44787_ (.A(_14238_),
    .B(_14233_),
    .C(_14229_),
    .Y(_14239_));
 sky130_fd_sc_hd__nand2_4 _44788_ (.A(_14237_),
    .B(_14239_),
    .Y(_14240_));
 sky130_fd_sc_hd__maj3_4 _44789_ (.A(_14004_),
    .B(_14002_),
    .C(_13987_),
    .X(_14241_));
 sky130_vsdinv _44790_ (.A(_14241_),
    .Y(_14242_));
 sky130_vsdinv _44791_ (.A(_13926_),
    .Y(_14243_));
 sky130_fd_sc_hd__a21boi_4 _44792_ (.A1(_13929_),
    .A2(_14243_),
    .B1_N(_13930_),
    .Y(_14244_));
 sky130_fd_sc_hd__nand2_4 _44793_ (.A(_13722_),
    .B(_14244_),
    .Y(_14245_));
 sky130_vsdinv _44794_ (.A(_14244_),
    .Y(_14246_));
 sky130_fd_sc_hd__nand3_4 _44795_ (.A(_14246_),
    .B(_13991_),
    .C(_13992_),
    .Y(_14247_));
 sky130_fd_sc_hd__buf_1 _44796_ (.A(_13997_),
    .X(_14248_));
 sky130_fd_sc_hd__a21o_4 _44797_ (.A1(_14245_),
    .A2(_14247_),
    .B1(_14248_),
    .X(_14249_));
 sky130_fd_sc_hd__nand3_4 _44798_ (.A(_14245_),
    .B(_14247_),
    .C(_13998_),
    .Y(_14250_));
 sky130_fd_sc_hd__nand2_4 _44799_ (.A(_14249_),
    .B(_14250_),
    .Y(_14251_));
 sky130_fd_sc_hd__a21o_4 _44800_ (.A1(_13925_),
    .A2(_13935_),
    .B1(_14251_),
    .X(_14252_));
 sky130_fd_sc_hd__a21oi_4 _44801_ (.A1(_13934_),
    .A2(_13932_),
    .B1(_13924_),
    .Y(_14253_));
 sky130_fd_sc_hd__nand2_4 _44802_ (.A(_14251_),
    .B(_14253_),
    .Y(_14254_));
 sky130_fd_sc_hd__nand2_4 _44803_ (.A(_14252_),
    .B(_14254_),
    .Y(_14255_));
 sky130_fd_sc_hd__maj3_4 _44804_ (.A(_13996_),
    .B(_13994_),
    .C(_13989_),
    .X(_14256_));
 sky130_fd_sc_hd__nand2_4 _44805_ (.A(_14255_),
    .B(_14256_),
    .Y(_14257_));
 sky130_vsdinv _44806_ (.A(_14256_),
    .Y(_14258_));
 sky130_fd_sc_hd__nand3_4 _44807_ (.A(_14252_),
    .B(_14254_),
    .C(_14258_),
    .Y(_14259_));
 sky130_fd_sc_hd__nand3_4 _44808_ (.A(_14242_),
    .B(_14257_),
    .C(_14259_),
    .Y(_14260_));
 sky130_fd_sc_hd__nand2_4 _44809_ (.A(_14257_),
    .B(_14259_),
    .Y(_14261_));
 sky130_fd_sc_hd__nand2_4 _44810_ (.A(_14261_),
    .B(_14241_),
    .Y(_14262_));
 sky130_fd_sc_hd__nand2_4 _44811_ (.A(_14260_),
    .B(_14262_),
    .Y(_14263_));
 sky130_fd_sc_hd__nand2_4 _44812_ (.A(_14263_),
    .B(_13479_),
    .Y(_14264_));
 sky130_fd_sc_hd__nand3_4 _44813_ (.A(_14260_),
    .B(_14262_),
    .C(_14015_),
    .Y(_14265_));
 sky130_fd_sc_hd__nand2_4 _44814_ (.A(_14264_),
    .B(_14265_),
    .Y(_14266_));
 sky130_fd_sc_hd__o21ai_4 _44815_ (.A1(_13969_),
    .A2(_13966_),
    .B1(_13967_),
    .Y(_14267_));
 sky130_vsdinv _44816_ (.A(_14267_),
    .Y(_14268_));
 sky130_fd_sc_hd__nand2_4 _44817_ (.A(_14266_),
    .B(_14268_),
    .Y(_14269_));
 sky130_fd_sc_hd__nand3_4 _44818_ (.A(_14267_),
    .B(_14264_),
    .C(_14265_),
    .Y(_14270_));
 sky130_fd_sc_hd__buf_1 _44819_ (.A(_14270_),
    .X(_14271_));
 sky130_fd_sc_hd__nand2_4 _44820_ (.A(_14269_),
    .B(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__buf_1 _44821_ (.A(_13482_),
    .X(_14273_));
 sky130_fd_sc_hd__a21boi_4 _44822_ (.A1(_14010_),
    .A2(_14273_),
    .B1_N(_14012_),
    .Y(_14274_));
 sky130_fd_sc_hd__nand2_4 _44823_ (.A(_14272_),
    .B(_14274_),
    .Y(_14275_));
 sky130_vsdinv _44824_ (.A(_14274_),
    .Y(_14276_));
 sky130_fd_sc_hd__nand3_4 _44825_ (.A(_14269_),
    .B(_14276_),
    .C(_14270_),
    .Y(_14277_));
 sky130_fd_sc_hd__nand2_4 _44826_ (.A(_14275_),
    .B(_14277_),
    .Y(_14278_));
 sky130_fd_sc_hd__nand2_4 _44827_ (.A(_14240_),
    .B(_14278_),
    .Y(_14279_));
 sky130_fd_sc_hd__a21oi_4 _44828_ (.A1(_14269_),
    .A2(_14271_),
    .B1(_14276_),
    .Y(_14280_));
 sky130_vsdinv _44829_ (.A(_14277_),
    .Y(_14281_));
 sky130_fd_sc_hd__nor2_4 _44830_ (.A(_14280_),
    .B(_14281_),
    .Y(_14282_));
 sky130_fd_sc_hd__nand3_4 _44831_ (.A(_14282_),
    .B(_14239_),
    .C(_14237_),
    .Y(_14283_));
 sky130_fd_sc_hd__nand2_4 _44832_ (.A(_14279_),
    .B(_14283_),
    .Y(_14284_));
 sky130_fd_sc_hd__a21boi_4 _44833_ (.A1(_14030_),
    .A2(_13980_),
    .B1_N(_13982_),
    .Y(_14285_));
 sky130_fd_sc_hd__nand2_4 _44834_ (.A(_14284_),
    .B(_14285_),
    .Y(_14286_));
 sky130_fd_sc_hd__a21oi_4 _44835_ (.A1(_13975_),
    .A2(_13976_),
    .B1(_13981_),
    .Y(_14287_));
 sky130_fd_sc_hd__o21ai_4 _44836_ (.A1(_14026_),
    .A2(_14287_),
    .B1(_13982_),
    .Y(_14288_));
 sky130_fd_sc_hd__nand3_4 _44837_ (.A(_14288_),
    .B(_14283_),
    .C(_14279_),
    .Y(_14289_));
 sky130_fd_sc_hd__nand2_4 _44838_ (.A(_14286_),
    .B(_14289_),
    .Y(_14290_));
 sky130_fd_sc_hd__buf_1 _44839_ (.A(_13775_),
    .X(_14291_));
 sky130_fd_sc_hd__a21boi_4 _44840_ (.A1(_14018_),
    .A2(_14024_),
    .B1_N(_14020_),
    .Y(_14292_));
 sky130_fd_sc_hd__xor2_4 _44841_ (.A(_14291_),
    .B(_14292_),
    .X(_14293_));
 sky130_fd_sc_hd__nand2_4 _44842_ (.A(_14290_),
    .B(_14293_),
    .Y(_14294_));
 sky130_vsdinv _44843_ (.A(_14293_),
    .Y(_14295_));
 sky130_fd_sc_hd__nand3_4 _44844_ (.A(_14286_),
    .B(_14289_),
    .C(_14295_),
    .Y(_14296_));
 sky130_fd_sc_hd__nand2_4 _44845_ (.A(_14294_),
    .B(_14296_),
    .Y(_14297_));
 sky130_fd_sc_hd__a21boi_4 _44846_ (.A1(_14034_),
    .A2(_14042_),
    .B1_N(_14037_),
    .Y(_14298_));
 sky130_fd_sc_hd__nand2_4 _44847_ (.A(_14297_),
    .B(_14298_),
    .Y(_14299_));
 sky130_fd_sc_hd__nand2_4 _44848_ (.A(_14043_),
    .B(_14037_),
    .Y(_14300_));
 sky130_fd_sc_hd__nand3_4 _44849_ (.A(_14300_),
    .B(_14296_),
    .C(_14294_),
    .Y(_14301_));
 sky130_fd_sc_hd__nand2_4 _44850_ (.A(_14299_),
    .B(_14301_),
    .Y(_14302_));
 sky130_fd_sc_hd__buf_1 _44851_ (.A(_13774_),
    .X(_14303_));
 sky130_fd_sc_hd__a21oi_4 _44852_ (.A1(_13760_),
    .A2(_13755_),
    .B1(_14303_),
    .Y(_14304_));
 sky130_vsdinv _44853_ (.A(_14304_),
    .Y(_14305_));
 sky130_fd_sc_hd__nand2_4 _44854_ (.A(_14302_),
    .B(_14305_),
    .Y(_14306_));
 sky130_fd_sc_hd__nand3_4 _44855_ (.A(_14299_),
    .B(_14301_),
    .C(_14304_),
    .Y(_14307_));
 sky130_fd_sc_hd__nand2_4 _44856_ (.A(_14306_),
    .B(_14307_),
    .Y(_14308_));
 sky130_fd_sc_hd__a21boi_4 _44857_ (.A1(_14046_),
    .A2(_14051_),
    .B1_N(_14048_),
    .Y(_14309_));
 sky130_fd_sc_hd__nand2_4 _44858_ (.A(_14308_),
    .B(_14309_),
    .Y(_14310_));
 sky130_fd_sc_hd__nand2_4 _44859_ (.A(_14054_),
    .B(_14048_),
    .Y(_14311_));
 sky130_fd_sc_hd__nand3_4 _44860_ (.A(_14311_),
    .B(_14307_),
    .C(_14306_),
    .Y(_14312_));
 sky130_fd_sc_hd__nand2_4 _44861_ (.A(_14310_),
    .B(_14312_),
    .Y(_14313_));
 sky130_fd_sc_hd__nor2_4 _44862_ (.A(_13796_),
    .B(_14059_),
    .Y(_14314_));
 sky130_fd_sc_hd__o21ai_4 _44863_ (.A1(_13802_),
    .A2(_13804_),
    .B1(_14314_),
    .Y(_14315_));
 sky130_fd_sc_hd__nand2_4 _44864_ (.A(_13795_),
    .B(_14058_),
    .Y(_14316_));
 sky130_fd_sc_hd__nand2_4 _44865_ (.A(_14316_),
    .B(_14057_),
    .Y(_14317_));
 sky130_fd_sc_hd__nand2_4 _44866_ (.A(_14315_),
    .B(_14317_),
    .Y(_14318_));
 sky130_fd_sc_hd__xnor2_4 _44867_ (.A(_14313_),
    .B(_14318_),
    .Y(_01447_));
 sky130_fd_sc_hd__a21boi_4 _44868_ (.A1(_14064_),
    .A2(_14066_),
    .B1_N(_14067_),
    .Y(_14319_));
 sky130_vsdinv _44869_ (.A(_14319_),
    .Y(_14320_));
 sky130_fd_sc_hd__nand2_4 _44870_ (.A(_08392_),
    .B(_03628_),
    .Y(_14321_));
 sky130_fd_sc_hd__o21ai_4 _44871_ (.A1(_10900_),
    .A2(_11432_),
    .B1(_14321_),
    .Y(_14322_));
 sky130_fd_sc_hd__nand2_4 _44872_ (.A(_07824_),
    .B(_11762_),
    .Y(_14323_));
 sky130_vsdinv _44873_ (.A(_14323_),
    .Y(_14324_));
 sky130_fd_sc_hd__nand4_4 _44874_ (.A(_03299_),
    .B(_06995_),
    .C(_12075_),
    .D(_12076_),
    .Y(_14325_));
 sky130_fd_sc_hd__nand3_4 _44875_ (.A(_14322_),
    .B(_14324_),
    .C(_14325_),
    .Y(_14326_));
 sky130_fd_sc_hd__nand2_4 _44876_ (.A(_14322_),
    .B(_14325_),
    .Y(_14327_));
 sky130_fd_sc_hd__nand2_4 _44877_ (.A(_14327_),
    .B(_14323_),
    .Y(_14328_));
 sky130_fd_sc_hd__nand3_4 _44878_ (.A(_14320_),
    .B(_14326_),
    .C(_14328_),
    .Y(_14329_));
 sky130_fd_sc_hd__nand2_4 _44879_ (.A(_14328_),
    .B(_14326_),
    .Y(_14330_));
 sky130_fd_sc_hd__nand2_4 _44880_ (.A(_14330_),
    .B(_14319_),
    .Y(_14331_));
 sky130_fd_sc_hd__nand2_4 _44881_ (.A(_14329_),
    .B(_14331_),
    .Y(_14332_));
 sky130_fd_sc_hd__nand2_4 _44882_ (.A(_13825_),
    .B(_11119_),
    .Y(_14333_));
 sky130_fd_sc_hd__nand2_4 _44883_ (.A(_07305_),
    .B(_11121_),
    .Y(_14334_));
 sky130_fd_sc_hd__nand2_4 _44884_ (.A(_14333_),
    .B(_14334_),
    .Y(_14335_));
 sky130_fd_sc_hd__nand4_4 _44885_ (.A(_13825_),
    .B(_07305_),
    .C(_11121_),
    .D(_11119_),
    .Y(_14336_));
 sky130_fd_sc_hd__nand2_4 _44886_ (.A(_07435_),
    .B(_10508_),
    .Y(_14337_));
 sky130_vsdinv _44887_ (.A(_14337_),
    .Y(_14338_));
 sky130_fd_sc_hd__a21o_4 _44888_ (.A1(_14335_),
    .A2(_14336_),
    .B1(_14338_),
    .X(_14339_));
 sky130_fd_sc_hd__nand3_4 _44889_ (.A(_14335_),
    .B(_14336_),
    .C(_14338_),
    .Y(_14340_));
 sky130_fd_sc_hd__nand2_4 _44890_ (.A(_14339_),
    .B(_14340_),
    .Y(_14341_));
 sky130_fd_sc_hd__nand2_4 _44891_ (.A(_14332_),
    .B(_14341_),
    .Y(_14342_));
 sky130_fd_sc_hd__nand4_4 _44892_ (.A(_14339_),
    .B(_14329_),
    .C(_14331_),
    .D(_14340_),
    .Y(_14343_));
 sky130_fd_sc_hd__nand2_4 _44893_ (.A(_14342_),
    .B(_14343_),
    .Y(_14344_));
 sky130_fd_sc_hd__a21boi_4 _44894_ (.A1(_14085_),
    .A2(_14073_),
    .B1_N(_14071_),
    .Y(_14345_));
 sky130_fd_sc_hd__nand2_4 _44895_ (.A(_14344_),
    .B(_14345_),
    .Y(_14346_));
 sky130_fd_sc_hd__nand2_4 _44896_ (.A(_14086_),
    .B(_14071_),
    .Y(_14347_));
 sky130_fd_sc_hd__nand3_4 _44897_ (.A(_14347_),
    .B(_14343_),
    .C(_14342_),
    .Y(_14348_));
 sky130_fd_sc_hd__nand2_4 _44898_ (.A(_14346_),
    .B(_14348_),
    .Y(_14349_));
 sky130_fd_sc_hd__nand2_4 _44899_ (.A(_08032_),
    .B(_10920_),
    .Y(_14350_));
 sky130_fd_sc_hd__nand2_4 _44900_ (.A(_07871_),
    .B(_03587_),
    .Y(_14351_));
 sky130_fd_sc_hd__nand2_4 _44901_ (.A(_14350_),
    .B(_14351_),
    .Y(_14352_));
 sky130_fd_sc_hd__nand4_4 _44902_ (.A(_11557_),
    .B(_11559_),
    .C(_12111_),
    .D(_10925_),
    .Y(_14353_));
 sky130_fd_sc_hd__nand2_4 _44903_ (.A(_10619_),
    .B(_11473_),
    .Y(_14354_));
 sky130_vsdinv _44904_ (.A(_14354_),
    .Y(_14355_));
 sky130_fd_sc_hd__a21o_4 _44905_ (.A1(_14352_),
    .A2(_14353_),
    .B1(_14355_),
    .X(_14356_));
 sky130_fd_sc_hd__nand3_4 _44906_ (.A(_14352_),
    .B(_14353_),
    .C(_14355_),
    .Y(_14357_));
 sky130_fd_sc_hd__nand2_4 _44907_ (.A(_14356_),
    .B(_14357_),
    .Y(_14358_));
 sky130_fd_sc_hd__a21boi_4 _44908_ (.A1(_14077_),
    .A2(_14080_),
    .B1_N(_14078_),
    .Y(_14359_));
 sky130_fd_sc_hd__nand2_4 _44909_ (.A(_14358_),
    .B(_14359_),
    .Y(_14360_));
 sky130_vsdinv _44910_ (.A(_14359_),
    .Y(_14361_));
 sky130_fd_sc_hd__nand3_4 _44911_ (.A(_14361_),
    .B(_14356_),
    .C(_14357_),
    .Y(_14362_));
 sky130_fd_sc_hd__a21boi_4 _44912_ (.A1(_14095_),
    .A2(_14099_),
    .B1_N(_14097_),
    .Y(_14363_));
 sky130_vsdinv _44913_ (.A(_14363_),
    .Y(_14364_));
 sky130_fd_sc_hd__a21o_4 _44914_ (.A1(_14360_),
    .A2(_14362_),
    .B1(_14364_),
    .X(_14365_));
 sky130_fd_sc_hd__nand3_4 _44915_ (.A(_14360_),
    .B(_14362_),
    .C(_14364_),
    .Y(_14366_));
 sky130_fd_sc_hd__nand2_4 _44916_ (.A(_14365_),
    .B(_14366_),
    .Y(_14367_));
 sky130_fd_sc_hd__nand2_4 _44917_ (.A(_14349_),
    .B(_14367_),
    .Y(_14368_));
 sky130_vsdinv _44918_ (.A(_14367_),
    .Y(_14369_));
 sky130_fd_sc_hd__nand3_4 _44919_ (.A(_14346_),
    .B(_14369_),
    .C(_14348_),
    .Y(_14370_));
 sky130_fd_sc_hd__nand2_4 _44920_ (.A(_14368_),
    .B(_14370_),
    .Y(_14371_));
 sky130_fd_sc_hd__a21boi_4 _44921_ (.A1(_14089_),
    .A2(_14113_),
    .B1_N(_14091_),
    .Y(_14372_));
 sky130_fd_sc_hd__nand2_4 _44922_ (.A(_14371_),
    .B(_14372_),
    .Y(_14373_));
 sky130_fd_sc_hd__nand2_4 _44923_ (.A(_14114_),
    .B(_14091_),
    .Y(_14374_));
 sky130_fd_sc_hd__nand3_4 _44924_ (.A(_14374_),
    .B(_14370_),
    .C(_14368_),
    .Y(_14375_));
 sky130_fd_sc_hd__nand2_4 _44925_ (.A(_14373_),
    .B(_14375_),
    .Y(_14376_));
 sky130_fd_sc_hd__buf_1 _44926_ (.A(_10537_),
    .X(_14377_));
 sky130_fd_sc_hd__nand2_4 _44927_ (.A(_08526_),
    .B(_14377_),
    .Y(_14378_));
 sky130_fd_sc_hd__nand2_4 _44928_ (.A(_08749_),
    .B(_11172_),
    .Y(_14379_));
 sky130_fd_sc_hd__nand2_4 _44929_ (.A(_14378_),
    .B(_14379_),
    .Y(_14380_));
 sky130_fd_sc_hd__nand4_4 _44930_ (.A(_11904_),
    .B(_08749_),
    .C(_08632_),
    .D(_14377_),
    .Y(_14381_));
 sky130_fd_sc_hd__nand2_4 _44931_ (.A(_13084_),
    .B(_03564_),
    .Y(_14382_));
 sky130_vsdinv _44932_ (.A(_14382_),
    .Y(_14383_));
 sky130_fd_sc_hd__a21o_4 _44933_ (.A1(_14380_),
    .A2(_14381_),
    .B1(_14383_),
    .X(_14384_));
 sky130_fd_sc_hd__nand3_4 _44934_ (.A(_14380_),
    .B(_14381_),
    .C(_14383_),
    .Y(_14385_));
 sky130_fd_sc_hd__a21boi_4 _44935_ (.A1(_14124_),
    .A2(_14127_),
    .B1_N(_14125_),
    .Y(_14386_));
 sky130_vsdinv _44936_ (.A(_14386_),
    .Y(_14387_));
 sky130_fd_sc_hd__a21o_4 _44937_ (.A1(_14384_),
    .A2(_14385_),
    .B1(_14387_),
    .X(_14388_));
 sky130_fd_sc_hd__nand3_4 _44938_ (.A(_14387_),
    .B(_14384_),
    .C(_14385_),
    .Y(_14389_));
 sky130_fd_sc_hd__nand2_4 _44939_ (.A(_10703_),
    .B(_12144_),
    .Y(_14390_));
 sky130_fd_sc_hd__nand2_4 _44940_ (.A(_13376_),
    .B(_08198_),
    .Y(_14391_));
 sky130_fd_sc_hd__nand2_4 _44941_ (.A(_12817_),
    .B(_12762_),
    .Y(_14392_));
 sky130_fd_sc_hd__nand2_4 _44942_ (.A(_14391_),
    .B(_14392_),
    .Y(_14393_));
 sky130_fd_sc_hd__nand4_4 _44943_ (.A(_12225_),
    .B(_09574_),
    .C(_12762_),
    .D(_11522_),
    .Y(_14394_));
 sky130_fd_sc_hd__nand2_4 _44944_ (.A(_14393_),
    .B(_14394_),
    .Y(_14395_));
 sky130_fd_sc_hd__xor2_4 _44945_ (.A(_14390_),
    .B(_14395_),
    .X(_14396_));
 sky130_fd_sc_hd__a21o_4 _44946_ (.A1(_14388_),
    .A2(_14389_),
    .B1(_14396_),
    .X(_14397_));
 sky130_fd_sc_hd__nand3_4 _44947_ (.A(_14388_),
    .B(_14396_),
    .C(_14389_),
    .Y(_14398_));
 sky130_fd_sc_hd__a21boi_4 _44948_ (.A1(_14104_),
    .A2(_14108_),
    .B1_N(_14106_),
    .Y(_14399_));
 sky130_vsdinv _44949_ (.A(_14399_),
    .Y(_14400_));
 sky130_fd_sc_hd__a21o_4 _44950_ (.A1(_14397_),
    .A2(_14398_),
    .B1(_14400_),
    .X(_14401_));
 sky130_fd_sc_hd__nand3_4 _44951_ (.A(_14397_),
    .B(_14400_),
    .C(_14398_),
    .Y(_14402_));
 sky130_fd_sc_hd__a21boi_4 _44952_ (.A1(_14132_),
    .A2(_14143_),
    .B1_N(_14133_),
    .Y(_14403_));
 sky130_vsdinv _44953_ (.A(_14403_),
    .Y(_14404_));
 sky130_fd_sc_hd__a21oi_4 _44954_ (.A1(_14401_),
    .A2(_14402_),
    .B1(_14404_),
    .Y(_14405_));
 sky130_vsdinv _44955_ (.A(_14405_),
    .Y(_14406_));
 sky130_fd_sc_hd__nand3_4 _44956_ (.A(_14401_),
    .B(_14404_),
    .C(_14402_),
    .Y(_14407_));
 sky130_fd_sc_hd__nand2_4 _44957_ (.A(_14406_),
    .B(_14407_),
    .Y(_14408_));
 sky130_fd_sc_hd__nand2_4 _44958_ (.A(_14376_),
    .B(_14408_),
    .Y(_14409_));
 sky130_vsdinv _44959_ (.A(_14407_),
    .Y(_14410_));
 sky130_fd_sc_hd__nor2_4 _44960_ (.A(_14405_),
    .B(_14410_),
    .Y(_14411_));
 sky130_fd_sc_hd__nand3_4 _44961_ (.A(_14411_),
    .B(_14375_),
    .C(_14373_),
    .Y(_14412_));
 sky130_fd_sc_hd__nand2_4 _44962_ (.A(_14409_),
    .B(_14412_),
    .Y(_14413_));
 sky130_fd_sc_hd__a21oi_4 _44963_ (.A1(_14114_),
    .A2(_14112_),
    .B1(_14119_),
    .Y(_14414_));
 sky130_fd_sc_hd__o21a_4 _44964_ (.A1(_14157_),
    .A2(_14414_),
    .B1(_14120_),
    .X(_14415_));
 sky130_fd_sc_hd__nand2_4 _44965_ (.A(_14413_),
    .B(_14415_),
    .Y(_14416_));
 sky130_fd_sc_hd__o21ai_4 _44966_ (.A1(_14157_),
    .A2(_14414_),
    .B1(_14120_),
    .Y(_14417_));
 sky130_fd_sc_hd__nand3_4 _44967_ (.A(_14417_),
    .B(_14409_),
    .C(_14412_),
    .Y(_14418_));
 sky130_fd_sc_hd__nand2_4 _44968_ (.A(_14416_),
    .B(_14418_),
    .Y(_14419_));
 sky130_fd_sc_hd__maj3_4 _44969_ (.A(_14136_),
    .B(_14138_),
    .C(_14135_),
    .X(_14420_));
 sky130_vsdinv _44970_ (.A(_14420_),
    .Y(_14421_));
 sky130_fd_sc_hd__nand2_4 _44971_ (.A(_12830_),
    .B(_07923_),
    .Y(_14422_));
 sky130_fd_sc_hd__nand2_4 _44972_ (.A(_10085_),
    .B(_13643_),
    .Y(_14423_));
 sky130_fd_sc_hd__nand2_4 _44973_ (.A(_14422_),
    .B(_14423_),
    .Y(_14424_));
 sky130_fd_sc_hd__nand4_4 _44974_ (.A(_13114_),
    .B(_12273_),
    .C(_13089_),
    .D(_12190_),
    .Y(_14425_));
 sky130_fd_sc_hd__buf_1 _44975_ (.A(_10406_),
    .X(_14426_));
 sky130_fd_sc_hd__nand2_4 _44976_ (.A(_14426_),
    .B(_03531_),
    .Y(_14427_));
 sky130_vsdinv _44977_ (.A(_14427_),
    .Y(_14428_));
 sky130_fd_sc_hd__a21o_4 _44978_ (.A1(_14424_),
    .A2(_14425_),
    .B1(_14428_),
    .X(_14429_));
 sky130_fd_sc_hd__nand3_4 _44979_ (.A(_14424_),
    .B(_14425_),
    .C(_14428_),
    .Y(_14430_));
 sky130_fd_sc_hd__nand3_4 _44980_ (.A(_14421_),
    .B(_14429_),
    .C(_14430_),
    .Y(_14431_));
 sky130_fd_sc_hd__nand2_4 _44981_ (.A(_14429_),
    .B(_14430_),
    .Y(_14432_));
 sky130_fd_sc_hd__nand2_4 _44982_ (.A(_14432_),
    .B(_14420_),
    .Y(_14433_));
 sky130_fd_sc_hd__a21boi_4 _44983_ (.A1(_14171_),
    .A2(_14174_),
    .B1_N(_14172_),
    .Y(_14434_));
 sky130_vsdinv _44984_ (.A(_14434_),
    .Y(_14435_));
 sky130_fd_sc_hd__a21o_4 _44985_ (.A1(_14431_),
    .A2(_14433_),
    .B1(_14435_),
    .X(_14436_));
 sky130_fd_sc_hd__nand3_4 _44986_ (.A(_14431_),
    .B(_14435_),
    .C(_14433_),
    .Y(_14437_));
 sky130_fd_sc_hd__nand2_4 _44987_ (.A(_14436_),
    .B(_14437_),
    .Y(_14438_));
 sky130_fd_sc_hd__maj3_4 _44988_ (.A(_14180_),
    .B(_14177_),
    .C(_14168_),
    .X(_14439_));
 sky130_fd_sc_hd__nand2_4 _44989_ (.A(_14438_),
    .B(_14439_),
    .Y(_14440_));
 sky130_vsdinv _44990_ (.A(_14439_),
    .Y(_14441_));
 sky130_fd_sc_hd__nand3_4 _44991_ (.A(_14441_),
    .B(_14437_),
    .C(_14436_),
    .Y(_14442_));
 sky130_fd_sc_hd__a21boi_4 _44992_ (.A1(_14193_),
    .A2(_14196_),
    .B1_N(_14194_),
    .Y(_14443_));
 sky130_fd_sc_hd__nand2_4 _44993_ (.A(_12878_),
    .B(_07741_),
    .Y(_14444_));
 sky130_fd_sc_hd__nand2_4 _44994_ (.A(_03396_),
    .B(_07189_),
    .Y(_14445_));
 sky130_fd_sc_hd__nand2_4 _44995_ (.A(_14444_),
    .B(_14445_),
    .Y(_14446_));
 sky130_fd_sc_hd__nand4_4 _44996_ (.A(_11673_),
    .B(_11675_),
    .C(_07192_),
    .D(_07194_),
    .Y(_14447_));
 sky130_fd_sc_hd__nand2_4 _44997_ (.A(_12310_),
    .B(_07197_),
    .Y(_14448_));
 sky130_vsdinv _44998_ (.A(_14448_),
    .Y(_14449_));
 sky130_fd_sc_hd__a21o_4 _44999_ (.A1(_14446_),
    .A2(_14447_),
    .B1(_14449_),
    .X(_14450_));
 sky130_fd_sc_hd__nand3_4 _45000_ (.A(_14446_),
    .B(_14447_),
    .C(_14449_),
    .Y(_14451_));
 sky130_fd_sc_hd__nand2_4 _45001_ (.A(_14450_),
    .B(_14451_),
    .Y(_14452_));
 sky130_fd_sc_hd__nor2_4 _45002_ (.A(_14443_),
    .B(_14452_),
    .Y(_14453_));
 sky130_vsdinv _45003_ (.A(_14453_),
    .Y(_14454_));
 sky130_fd_sc_hd__nand2_4 _45004_ (.A(_14452_),
    .B(_14443_),
    .Y(_14455_));
 sky130_fd_sc_hd__o21ai_4 _45005_ (.A1(_06505_),
    .A2(_06636_),
    .B1(_03406_),
    .Y(_14456_));
 sky130_vsdinv _45006_ (.A(_14456_),
    .Y(_14457_));
 sky130_fd_sc_hd__nand3_4 _45007_ (.A(_03406_),
    .B(_07212_),
    .C(_07214_),
    .Y(_14458_));
 sky130_fd_sc_hd__a21o_4 _45008_ (.A1(_14457_),
    .A2(_14458_),
    .B1(_14243_),
    .X(_14459_));
 sky130_fd_sc_hd__nand3_4 _45009_ (.A(_14457_),
    .B(_14243_),
    .C(_14458_),
    .Y(_14460_));
 sky130_fd_sc_hd__nand2_4 _45010_ (.A(_14459_),
    .B(_14460_),
    .Y(_14461_));
 sky130_vsdinv _45011_ (.A(_14461_),
    .Y(_14462_));
 sky130_fd_sc_hd__buf_1 _45012_ (.A(_14462_),
    .X(_14463_));
 sky130_fd_sc_hd__buf_1 _45013_ (.A(_14463_),
    .X(_14464_));
 sky130_fd_sc_hd__a21oi_4 _45014_ (.A1(_14454_),
    .A2(_14455_),
    .B1(_14464_),
    .Y(_14465_));
 sky130_fd_sc_hd__nand3_4 _45015_ (.A(_14454_),
    .B(_14463_),
    .C(_14455_),
    .Y(_14466_));
 sky130_vsdinv _45016_ (.A(_14466_),
    .Y(_14467_));
 sky130_fd_sc_hd__nor2_4 _45017_ (.A(_14465_),
    .B(_14467_),
    .Y(_14468_));
 sky130_fd_sc_hd__a21o_4 _45018_ (.A1(_14440_),
    .A2(_14442_),
    .B1(_14468_),
    .X(_14469_));
 sky130_fd_sc_hd__nand3_4 _45019_ (.A(_14440_),
    .B(_14442_),
    .C(_14468_),
    .Y(_14470_));
 sky130_fd_sc_hd__nand2_4 _45020_ (.A(_14469_),
    .B(_14470_),
    .Y(_14471_));
 sky130_fd_sc_hd__o21ai_4 _45021_ (.A1(_14152_),
    .A2(_14148_),
    .B1(_14149_),
    .Y(_14472_));
 sky130_vsdinv _45022_ (.A(_14472_),
    .Y(_14473_));
 sky130_fd_sc_hd__nand2_4 _45023_ (.A(_14471_),
    .B(_14473_),
    .Y(_14474_));
 sky130_fd_sc_hd__nand3_4 _45024_ (.A(_14469_),
    .B(_14472_),
    .C(_14470_),
    .Y(_14475_));
 sky130_fd_sc_hd__a21boi_4 _45025_ (.A1(_14186_),
    .A2(_14214_),
    .B1_N(_14188_),
    .Y(_14476_));
 sky130_vsdinv _45026_ (.A(_14476_),
    .Y(_14477_));
 sky130_fd_sc_hd__a21oi_4 _45027_ (.A1(_14474_),
    .A2(_14475_),
    .B1(_14477_),
    .Y(_14478_));
 sky130_vsdinv _45028_ (.A(_14478_),
    .Y(_14479_));
 sky130_fd_sc_hd__nand3_4 _45029_ (.A(_14474_),
    .B(_14477_),
    .C(_14475_),
    .Y(_14480_));
 sky130_fd_sc_hd__nand2_4 _45030_ (.A(_14479_),
    .B(_14480_),
    .Y(_14481_));
 sky130_fd_sc_hd__nand2_4 _45031_ (.A(_14419_),
    .B(_14481_),
    .Y(_14482_));
 sky130_vsdinv _45032_ (.A(_14480_),
    .Y(_14483_));
 sky130_fd_sc_hd__nor2_4 _45033_ (.A(_14478_),
    .B(_14483_),
    .Y(_14484_));
 sky130_fd_sc_hd__nand3_4 _45034_ (.A(_14484_),
    .B(_14416_),
    .C(_14418_),
    .Y(_14485_));
 sky130_fd_sc_hd__nand2_4 _45035_ (.A(_14482_),
    .B(_14485_),
    .Y(_14486_));
 sky130_fd_sc_hd__a21boi_4 _45036_ (.A1(_14232_),
    .A2(_14163_),
    .B1_N(_14165_),
    .Y(_14487_));
 sky130_fd_sc_hd__nand2_4 _45037_ (.A(_14486_),
    .B(_14487_),
    .Y(_14488_));
 sky130_fd_sc_hd__a21oi_4 _45038_ (.A1(_14158_),
    .A2(_14159_),
    .B1(_14164_),
    .Y(_14489_));
 sky130_fd_sc_hd__o21ai_4 _45039_ (.A1(_14489_),
    .A2(_14228_),
    .B1(_14165_),
    .Y(_14490_));
 sky130_fd_sc_hd__nand3_4 _45040_ (.A(_14490_),
    .B(_14485_),
    .C(_14482_),
    .Y(_14491_));
 sky130_fd_sc_hd__nand2_4 _45041_ (.A(_14488_),
    .B(_14491_),
    .Y(_14492_));
 sky130_fd_sc_hd__a21oi_4 _45042_ (.A1(_14203_),
    .A2(_14210_),
    .B1(_14200_),
    .Y(_14493_));
 sky130_vsdinv _45043_ (.A(_14493_),
    .Y(_14494_));
 sky130_fd_sc_hd__a21boi_4 _45044_ (.A1(_14207_),
    .A2(_14243_),
    .B1_N(_14208_),
    .Y(_14495_));
 sky130_fd_sc_hd__nand2_4 _45045_ (.A(_13722_),
    .B(_14495_),
    .Y(_14496_));
 sky130_vsdinv _45046_ (.A(_14495_),
    .Y(_14497_));
 sky130_fd_sc_hd__nand3_4 _45047_ (.A(_14497_),
    .B(_13992_),
    .C(_13991_),
    .Y(_14498_));
 sky130_fd_sc_hd__buf_1 _45048_ (.A(_14248_),
    .X(_14499_));
 sky130_fd_sc_hd__nand3_4 _45049_ (.A(_14496_),
    .B(_14498_),
    .C(_14499_),
    .Y(_14500_));
 sky130_fd_sc_hd__a21o_4 _45050_ (.A1(_14496_),
    .A2(_14498_),
    .B1(_13998_),
    .X(_14501_));
 sky130_fd_sc_hd__nand3_4 _45051_ (.A(_14494_),
    .B(_14500_),
    .C(_14501_),
    .Y(_14502_));
 sky130_fd_sc_hd__nand2_4 _45052_ (.A(_14501_),
    .B(_14500_),
    .Y(_14503_));
 sky130_fd_sc_hd__nand2_4 _45053_ (.A(_14503_),
    .B(_14493_),
    .Y(_14504_));
 sky130_fd_sc_hd__a21boi_4 _45054_ (.A1(_14245_),
    .A2(_14499_),
    .B1_N(_14247_),
    .Y(_14505_));
 sky130_vsdinv _45055_ (.A(_14505_),
    .Y(_14506_));
 sky130_fd_sc_hd__a21o_4 _45056_ (.A1(_14502_),
    .A2(_14504_),
    .B1(_14506_),
    .X(_14507_));
 sky130_fd_sc_hd__nand3_4 _45057_ (.A(_14502_),
    .B(_14504_),
    .C(_14506_),
    .Y(_14508_));
 sky130_fd_sc_hd__nand2_4 _45058_ (.A(_14507_),
    .B(_14508_),
    .Y(_14509_));
 sky130_fd_sc_hd__maj3_4 _45059_ (.A(_14256_),
    .B(_14251_),
    .C(_14253_),
    .X(_14510_));
 sky130_fd_sc_hd__nand2_4 _45060_ (.A(_14509_),
    .B(_14510_),
    .Y(_14511_));
 sky130_vsdinv _45061_ (.A(_14510_),
    .Y(_14512_));
 sky130_fd_sc_hd__nand3_4 _45062_ (.A(_14512_),
    .B(_14507_),
    .C(_14508_),
    .Y(_14513_));
 sky130_fd_sc_hd__nand2_4 _45063_ (.A(_14511_),
    .B(_14513_),
    .Y(_14514_));
 sky130_fd_sc_hd__nand2_4 _45064_ (.A(_14514_),
    .B(_13745_),
    .Y(_14515_));
 sky130_fd_sc_hd__nand3_4 _45065_ (.A(_14511_),
    .B(_14513_),
    .C(_13747_),
    .Y(_14516_));
 sky130_fd_sc_hd__nand2_4 _45066_ (.A(_14515_),
    .B(_14516_),
    .Y(_14517_));
 sky130_fd_sc_hd__a21boi_4 _45067_ (.A1(_14221_),
    .A2(_14225_),
    .B1_N(_14223_),
    .Y(_14518_));
 sky130_fd_sc_hd__nand2_4 _45068_ (.A(_14517_),
    .B(_14518_),
    .Y(_14519_));
 sky130_fd_sc_hd__a21oi_4 _45069_ (.A1(_14216_),
    .A2(_14217_),
    .B1(_14219_),
    .Y(_14520_));
 sky130_fd_sc_hd__o21ai_4 _45070_ (.A1(_14224_),
    .A2(_14520_),
    .B1(_14223_),
    .Y(_14521_));
 sky130_fd_sc_hd__nand3_4 _45071_ (.A(_14521_),
    .B(_14515_),
    .C(_14516_),
    .Y(_14522_));
 sky130_fd_sc_hd__a21boi_4 _45072_ (.A1(_13756_),
    .A2(_14262_),
    .B1_N(_14260_),
    .Y(_14523_));
 sky130_vsdinv _45073_ (.A(_14523_),
    .Y(_14524_));
 sky130_fd_sc_hd__a21oi_4 _45074_ (.A1(_14519_),
    .A2(_14522_),
    .B1(_14524_),
    .Y(_14525_));
 sky130_vsdinv _45075_ (.A(_14525_),
    .Y(_14526_));
 sky130_fd_sc_hd__nand3_4 _45076_ (.A(_14519_),
    .B(_14524_),
    .C(_14522_),
    .Y(_14527_));
 sky130_fd_sc_hd__nand2_4 _45077_ (.A(_14526_),
    .B(_14527_),
    .Y(_14528_));
 sky130_fd_sc_hd__nand2_4 _45078_ (.A(_14492_),
    .B(_14528_),
    .Y(_14529_));
 sky130_vsdinv _45079_ (.A(_14527_),
    .Y(_14530_));
 sky130_fd_sc_hd__nor2_4 _45080_ (.A(_14525_),
    .B(_14530_),
    .Y(_14531_));
 sky130_fd_sc_hd__nand3_4 _45081_ (.A(_14531_),
    .B(_14488_),
    .C(_14491_),
    .Y(_14532_));
 sky130_fd_sc_hd__nand2_4 _45082_ (.A(_14529_),
    .B(_14532_),
    .Y(_14533_));
 sky130_fd_sc_hd__a21boi_4 _45083_ (.A1(_14282_),
    .A2(_14237_),
    .B1_N(_14239_),
    .Y(_14534_));
 sky130_fd_sc_hd__nand2_4 _45084_ (.A(_14533_),
    .B(_14534_),
    .Y(_14535_));
 sky130_fd_sc_hd__a21oi_4 _45085_ (.A1(_14233_),
    .A2(_14229_),
    .B1(_14238_),
    .Y(_14536_));
 sky130_fd_sc_hd__o21ai_4 _45086_ (.A1(_14278_),
    .A2(_14536_),
    .B1(_14239_),
    .Y(_14537_));
 sky130_fd_sc_hd__nand3_4 _45087_ (.A(_14537_),
    .B(_14529_),
    .C(_14532_),
    .Y(_14538_));
 sky130_fd_sc_hd__nand2_4 _45088_ (.A(_14535_),
    .B(_14538_),
    .Y(_14539_));
 sky130_fd_sc_hd__a21boi_4 _45089_ (.A1(_14269_),
    .A2(_14276_),
    .B1_N(_14271_),
    .Y(_14540_));
 sky130_fd_sc_hd__xor2_4 _45090_ (.A(_14291_),
    .B(_14540_),
    .X(_14541_));
 sky130_fd_sc_hd__nand2_4 _45091_ (.A(_14539_),
    .B(_14541_),
    .Y(_14542_));
 sky130_vsdinv _45092_ (.A(_14541_),
    .Y(_14543_));
 sky130_fd_sc_hd__nand3_4 _45093_ (.A(_14535_),
    .B(_14538_),
    .C(_14543_),
    .Y(_14544_));
 sky130_fd_sc_hd__nand2_4 _45094_ (.A(_14542_),
    .B(_14544_),
    .Y(_14545_));
 sky130_fd_sc_hd__a21boi_4 _45095_ (.A1(_14286_),
    .A2(_14295_),
    .B1_N(_14289_),
    .Y(_14546_));
 sky130_fd_sc_hd__nand2_4 _45096_ (.A(_14545_),
    .B(_14546_),
    .Y(_14547_));
 sky130_fd_sc_hd__nand2_4 _45097_ (.A(_14296_),
    .B(_14289_),
    .Y(_14548_));
 sky130_fd_sc_hd__nand3_4 _45098_ (.A(_14548_),
    .B(_14542_),
    .C(_14544_),
    .Y(_14549_));
 sky130_fd_sc_hd__nand2_4 _45099_ (.A(_14547_),
    .B(_14549_),
    .Y(_14550_));
 sky130_fd_sc_hd__a21oi_4 _45100_ (.A1(_14025_),
    .A2(_14020_),
    .B1(_14303_),
    .Y(_14551_));
 sky130_vsdinv _45101_ (.A(_14551_),
    .Y(_14552_));
 sky130_fd_sc_hd__nand2_4 _45102_ (.A(_14550_),
    .B(_14552_),
    .Y(_14553_));
 sky130_fd_sc_hd__nand3_4 _45103_ (.A(_14547_),
    .B(_14549_),
    .C(_14551_),
    .Y(_14554_));
 sky130_fd_sc_hd__nand2_4 _45104_ (.A(_14553_),
    .B(_14554_),
    .Y(_14555_));
 sky130_fd_sc_hd__a21boi_4 _45105_ (.A1(_14299_),
    .A2(_14304_),
    .B1_N(_14301_),
    .Y(_14556_));
 sky130_fd_sc_hd__nand2_4 _45106_ (.A(_14555_),
    .B(_14556_),
    .Y(_14557_));
 sky130_fd_sc_hd__nand2_4 _45107_ (.A(_14307_),
    .B(_14301_),
    .Y(_14558_));
 sky130_fd_sc_hd__nand3_4 _45108_ (.A(_14558_),
    .B(_14554_),
    .C(_14553_),
    .Y(_14559_));
 sky130_fd_sc_hd__nand2_4 _45109_ (.A(_14557_),
    .B(_14559_),
    .Y(_14560_));
 sky130_vsdinv _45110_ (.A(_14312_),
    .Y(_14561_));
 sky130_fd_sc_hd__a21oi_4 _45111_ (.A1(_14318_),
    .A2(_14310_),
    .B1(_14561_),
    .Y(_14562_));
 sky130_fd_sc_hd__xor2_4 _45112_ (.A(_14560_),
    .B(_14562_),
    .X(_01448_));
 sky130_fd_sc_hd__nand2_4 _45113_ (.A(_10584_),
    .B(_11105_),
    .Y(_14563_));
 sky130_fd_sc_hd__o21ai_4 _45114_ (.A1(_08835_),
    .A2(_13808_),
    .B1(_14563_),
    .Y(_14564_));
 sky130_fd_sc_hd__buf_1 _45115_ (.A(_11106_),
    .X(_14565_));
 sky130_fd_sc_hd__nand4_4 _45116_ (.A(_03304_),
    .B(_07286_),
    .C(_10959_),
    .D(_14565_),
    .Y(_14566_));
 sky130_fd_sc_hd__nand2_4 _45117_ (.A(_10989_),
    .B(_10955_),
    .Y(_14567_));
 sky130_vsdinv _45118_ (.A(_14567_),
    .Y(_14568_));
 sky130_fd_sc_hd__a21o_4 _45119_ (.A1(_14564_),
    .A2(_14566_),
    .B1(_14568_),
    .X(_14569_));
 sky130_fd_sc_hd__nand3_4 _45120_ (.A(_14564_),
    .B(_14568_),
    .C(_14566_),
    .Y(_14570_));
 sky130_fd_sc_hd__nand2_4 _45121_ (.A(_14569_),
    .B(_14570_),
    .Y(_14571_));
 sky130_fd_sc_hd__a21boi_4 _45122_ (.A1(_14322_),
    .A2(_14324_),
    .B1_N(_14325_),
    .Y(_14572_));
 sky130_fd_sc_hd__nand2_4 _45123_ (.A(_14571_),
    .B(_14572_),
    .Y(_14573_));
 sky130_vsdinv _45124_ (.A(_14572_),
    .Y(_14574_));
 sky130_fd_sc_hd__nand3_4 _45125_ (.A(_14574_),
    .B(_14570_),
    .C(_14569_),
    .Y(_14575_));
 sky130_fd_sc_hd__nand2_4 _45126_ (.A(_14096_),
    .B(_10512_),
    .Y(_14576_));
 sky130_fd_sc_hd__nand2_4 _45127_ (.A(_07302_),
    .B(_12093_),
    .Y(_14577_));
 sky130_fd_sc_hd__nand2_4 _45128_ (.A(_13331_),
    .B(_12092_),
    .Y(_14578_));
 sky130_fd_sc_hd__nand2_4 _45129_ (.A(_14577_),
    .B(_14578_),
    .Y(_14579_));
 sky130_fd_sc_hd__nand4_4 _45130_ (.A(_07306_),
    .B(_12458_),
    .C(_12409_),
    .D(_12410_),
    .Y(_14580_));
 sky130_fd_sc_hd__nand2_4 _45131_ (.A(_14579_),
    .B(_14580_),
    .Y(_14581_));
 sky130_fd_sc_hd__xor2_4 _45132_ (.A(_14576_),
    .B(_14581_),
    .X(_14582_));
 sky130_fd_sc_hd__a21o_4 _45133_ (.A1(_14573_),
    .A2(_14575_),
    .B1(_14582_),
    .X(_14583_));
 sky130_fd_sc_hd__nand3_4 _45134_ (.A(_14573_),
    .B(_14575_),
    .C(_14582_),
    .Y(_14584_));
 sky130_fd_sc_hd__nand2_4 _45135_ (.A(_14583_),
    .B(_14584_),
    .Y(_14585_));
 sky130_fd_sc_hd__maj3_4 _45136_ (.A(_14341_),
    .B(_14330_),
    .C(_14319_),
    .X(_14586_));
 sky130_fd_sc_hd__nand2_4 _45137_ (.A(_14585_),
    .B(_14586_),
    .Y(_14587_));
 sky130_fd_sc_hd__nand2_4 _45138_ (.A(_14343_),
    .B(_14329_),
    .Y(_14588_));
 sky130_fd_sc_hd__nand3_4 _45139_ (.A(_14588_),
    .B(_14584_),
    .C(_14583_),
    .Y(_14589_));
 sky130_fd_sc_hd__nand2_4 _45140_ (.A(_14587_),
    .B(_14589_),
    .Y(_14590_));
 sky130_fd_sc_hd__nand2_4 _45141_ (.A(_08042_),
    .B(_10305_),
    .Y(_14591_));
 sky130_fd_sc_hd__nand2_4 _45142_ (.A(_09070_),
    .B(_10481_),
    .Y(_14592_));
 sky130_fd_sc_hd__nand2_4 _45143_ (.A(_14591_),
    .B(_14592_),
    .Y(_14593_));
 sky130_fd_sc_hd__nand4_4 _45144_ (.A(_08051_),
    .B(_08052_),
    .C(_13011_),
    .D(_03596_),
    .Y(_14594_));
 sky130_fd_sc_hd__nand2_4 _45145_ (.A(_08056_),
    .B(_11473_),
    .Y(_14595_));
 sky130_vsdinv _45146_ (.A(_14595_),
    .Y(_14596_));
 sky130_fd_sc_hd__a21o_4 _45147_ (.A1(_14593_),
    .A2(_14594_),
    .B1(_14596_),
    .X(_14597_));
 sky130_fd_sc_hd__nand3_4 _45148_ (.A(_14593_),
    .B(_14594_),
    .C(_14596_),
    .Y(_14598_));
 sky130_fd_sc_hd__a21boi_4 _45149_ (.A1(_14335_),
    .A2(_14338_),
    .B1_N(_14336_),
    .Y(_14599_));
 sky130_fd_sc_hd__a21boi_4 _45150_ (.A1(_14597_),
    .A2(_14598_),
    .B1_N(_14599_),
    .Y(_14600_));
 sky130_vsdinv _45151_ (.A(_14600_),
    .Y(_14601_));
 sky130_vsdinv _45152_ (.A(_14599_),
    .Y(_14602_));
 sky130_fd_sc_hd__nand3_4 _45153_ (.A(_14602_),
    .B(_14597_),
    .C(_14598_),
    .Y(_14603_));
 sky130_fd_sc_hd__a21boi_4 _45154_ (.A1(_14352_),
    .A2(_14355_),
    .B1_N(_14353_),
    .Y(_14604_));
 sky130_vsdinv _45155_ (.A(_14604_),
    .Y(_14605_));
 sky130_fd_sc_hd__a21oi_4 _45156_ (.A1(_14601_),
    .A2(_14603_),
    .B1(_14605_),
    .Y(_14606_));
 sky130_vsdinv _45157_ (.A(_14606_),
    .Y(_14607_));
 sky130_fd_sc_hd__nand3_4 _45158_ (.A(_14601_),
    .B(_14605_),
    .C(_14603_),
    .Y(_14608_));
 sky130_fd_sc_hd__nand2_4 _45159_ (.A(_14607_),
    .B(_14608_),
    .Y(_14609_));
 sky130_fd_sc_hd__nand2_4 _45160_ (.A(_14590_),
    .B(_14609_),
    .Y(_14610_));
 sky130_vsdinv _45161_ (.A(_14609_),
    .Y(_14611_));
 sky130_fd_sc_hd__nand3_4 _45162_ (.A(_14611_),
    .B(_14589_),
    .C(_14587_),
    .Y(_14612_));
 sky130_fd_sc_hd__nand2_4 _45163_ (.A(_14610_),
    .B(_14612_),
    .Y(_14613_));
 sky130_fd_sc_hd__a21boi_4 _45164_ (.A1(_14346_),
    .A2(_14369_),
    .B1_N(_14348_),
    .Y(_14614_));
 sky130_fd_sc_hd__nand2_4 _45165_ (.A(_14613_),
    .B(_14614_),
    .Y(_14615_));
 sky130_vsdinv _45166_ (.A(_14614_),
    .Y(_14616_));
 sky130_fd_sc_hd__nand3_4 _45167_ (.A(_14616_),
    .B(_14612_),
    .C(_14610_),
    .Y(_14617_));
 sky130_fd_sc_hd__nand2_4 _45168_ (.A(_14615_),
    .B(_14617_),
    .Y(_14618_));
 sky130_fd_sc_hd__nand2_4 _45169_ (.A(_12220_),
    .B(_12467_),
    .Y(_14619_));
 sky130_fd_sc_hd__nand2_4 _45170_ (.A(_11593_),
    .B(_12466_),
    .Y(_14620_));
 sky130_fd_sc_hd__nand2_4 _45171_ (.A(_14619_),
    .B(_14620_),
    .Y(_14621_));
 sky130_fd_sc_hd__nand4_4 _45172_ (.A(_12220_),
    .B(_11593_),
    .C(_12466_),
    .D(_11173_),
    .Y(_14622_));
 sky130_fd_sc_hd__nand2_4 _45173_ (.A(_11595_),
    .B(_03564_),
    .Y(_14623_));
 sky130_vsdinv _45174_ (.A(_14623_),
    .Y(_14624_));
 sky130_fd_sc_hd__a21o_4 _45175_ (.A1(_14621_),
    .A2(_14622_),
    .B1(_14624_),
    .X(_14625_));
 sky130_fd_sc_hd__nand3_4 _45176_ (.A(_14621_),
    .B(_14622_),
    .C(_14624_),
    .Y(_14626_));
 sky130_fd_sc_hd__nand2_4 _45177_ (.A(_14625_),
    .B(_14626_),
    .Y(_14627_));
 sky130_fd_sc_hd__a21o_4 _45178_ (.A1(_14381_),
    .A2(_14385_),
    .B1(_14627_),
    .X(_14628_));
 sky130_fd_sc_hd__nand3_4 _45179_ (.A(_14627_),
    .B(_14381_),
    .C(_14385_),
    .Y(_14629_));
 sky130_fd_sc_hd__nand2_4 _45180_ (.A(_13114_),
    .B(_11514_),
    .Y(_14630_));
 sky130_fd_sc_hd__nand2_4 _45181_ (.A(_13943_),
    .B(_11516_),
    .Y(_14631_));
 sky130_fd_sc_hd__nand2_4 _45182_ (.A(_12821_),
    .B(_11186_),
    .Y(_14632_));
 sky130_fd_sc_hd__nand2_4 _45183_ (.A(_14631_),
    .B(_14632_),
    .Y(_14633_));
 sky130_fd_sc_hd__nand4_4 _45184_ (.A(_12533_),
    .B(_12233_),
    .C(_13884_),
    .D(_13885_),
    .Y(_14634_));
 sky130_fd_sc_hd__nand2_4 _45185_ (.A(_14633_),
    .B(_14634_),
    .Y(_14635_));
 sky130_fd_sc_hd__xor2_4 _45186_ (.A(_14630_),
    .B(_14635_),
    .X(_14636_));
 sky130_fd_sc_hd__a21o_4 _45187_ (.A1(_14628_),
    .A2(_14629_),
    .B1(_14636_),
    .X(_14637_));
 sky130_fd_sc_hd__nand3_4 _45188_ (.A(_14628_),
    .B(_14636_),
    .C(_14629_),
    .Y(_14638_));
 sky130_fd_sc_hd__a21boi_4 _45189_ (.A1(_14360_),
    .A2(_14364_),
    .B1_N(_14362_),
    .Y(_14639_));
 sky130_vsdinv _45190_ (.A(_14639_),
    .Y(_14640_));
 sky130_fd_sc_hd__a21oi_4 _45191_ (.A1(_14637_),
    .A2(_14638_),
    .B1(_14640_),
    .Y(_14641_));
 sky130_fd_sc_hd__nand3_4 _45192_ (.A(_14637_),
    .B(_14640_),
    .C(_14638_),
    .Y(_14642_));
 sky130_vsdinv _45193_ (.A(_14642_),
    .Y(_14643_));
 sky130_vsdinv _45194_ (.A(_14389_),
    .Y(_14644_));
 sky130_fd_sc_hd__a21oi_4 _45195_ (.A1(_14388_),
    .A2(_14396_),
    .B1(_14644_),
    .Y(_14645_));
 sky130_fd_sc_hd__o21ai_4 _45196_ (.A1(_14641_),
    .A2(_14643_),
    .B1(_14645_),
    .Y(_14646_));
 sky130_vsdinv _45197_ (.A(_14641_),
    .Y(_14647_));
 sky130_vsdinv _45198_ (.A(_14645_),
    .Y(_14648_));
 sky130_fd_sc_hd__nand3_4 _45199_ (.A(_14647_),
    .B(_14648_),
    .C(_14642_),
    .Y(_14649_));
 sky130_fd_sc_hd__nand2_4 _45200_ (.A(_14646_),
    .B(_14649_),
    .Y(_14650_));
 sky130_fd_sc_hd__nand2_4 _45201_ (.A(_14618_),
    .B(_14650_),
    .Y(_14651_));
 sky130_fd_sc_hd__nand4_4 _45202_ (.A(_14649_),
    .B(_14615_),
    .C(_14646_),
    .D(_14617_),
    .Y(_14652_));
 sky130_fd_sc_hd__nand2_4 _45203_ (.A(_14651_),
    .B(_14652_),
    .Y(_14653_));
 sky130_fd_sc_hd__a21boi_4 _45204_ (.A1(_14411_),
    .A2(_14373_),
    .B1_N(_14375_),
    .Y(_14654_));
 sky130_fd_sc_hd__nand2_4 _45205_ (.A(_14653_),
    .B(_14654_),
    .Y(_14655_));
 sky130_vsdinv _45206_ (.A(_14654_),
    .Y(_14656_));
 sky130_fd_sc_hd__nand3_4 _45207_ (.A(_14656_),
    .B(_14651_),
    .C(_14652_),
    .Y(_14657_));
 sky130_fd_sc_hd__nand2_4 _45208_ (.A(_14655_),
    .B(_14657_),
    .Y(_14658_));
 sky130_fd_sc_hd__nand2_4 _45209_ (.A(_03383_),
    .B(_07717_),
    .Y(_14659_));
 sky130_fd_sc_hd__nand2_4 _45210_ (.A(_11319_),
    .B(_10990_),
    .Y(_14660_));
 sky130_fd_sc_hd__nand2_4 _45211_ (.A(_14659_),
    .B(_14660_),
    .Y(_14661_));
 sky130_fd_sc_hd__nand4_4 _45212_ (.A(_12832_),
    .B(_13124_),
    .C(_07554_),
    .D(_07557_),
    .Y(_14662_));
 sky130_fd_sc_hd__nand2_4 _45213_ (.A(_11673_),
    .B(_08132_),
    .Y(_14663_));
 sky130_vsdinv _45214_ (.A(_14663_),
    .Y(_14664_));
 sky130_fd_sc_hd__a21o_4 _45215_ (.A1(_14661_),
    .A2(_14662_),
    .B1(_14664_),
    .X(_14665_));
 sky130_fd_sc_hd__nand3_4 _45216_ (.A(_14661_),
    .B(_14662_),
    .C(_14664_),
    .Y(_14666_));
 sky130_vsdinv _45217_ (.A(_14390_),
    .Y(_14667_));
 sky130_fd_sc_hd__a21boi_4 _45218_ (.A1(_14393_),
    .A2(_14667_),
    .B1_N(_14394_),
    .Y(_14668_));
 sky130_fd_sc_hd__a21boi_4 _45219_ (.A1(_14665_),
    .A2(_14666_),
    .B1_N(_14668_),
    .Y(_14669_));
 sky130_vsdinv _45220_ (.A(_14669_),
    .Y(_14670_));
 sky130_vsdinv _45221_ (.A(_14668_),
    .Y(_14671_));
 sky130_fd_sc_hd__nand3_4 _45222_ (.A(_14671_),
    .B(_14665_),
    .C(_14666_),
    .Y(_14672_));
 sky130_fd_sc_hd__nand2_4 _45223_ (.A(_14670_),
    .B(_14672_),
    .Y(_14673_));
 sky130_fd_sc_hd__a21o_4 _45224_ (.A1(_14425_),
    .A2(_14430_),
    .B1(_14673_),
    .X(_14674_));
 sky130_fd_sc_hd__a21boi_4 _45225_ (.A1(_14424_),
    .A2(_14428_),
    .B1_N(_14425_),
    .Y(_14675_));
 sky130_fd_sc_hd__nand2_4 _45226_ (.A(_14673_),
    .B(_14675_),
    .Y(_14676_));
 sky130_fd_sc_hd__nand2_4 _45227_ (.A(_14674_),
    .B(_14676_),
    .Y(_14677_));
 sky130_fd_sc_hd__maj3_4 _45228_ (.A(_14434_),
    .B(_14432_),
    .C(_14420_),
    .X(_14678_));
 sky130_fd_sc_hd__nand2_4 _45229_ (.A(_14677_),
    .B(_14678_),
    .Y(_14679_));
 sky130_vsdinv _45230_ (.A(_14678_),
    .Y(_14680_));
 sky130_fd_sc_hd__nand3_4 _45231_ (.A(_14674_),
    .B(_14676_),
    .C(_14680_),
    .Y(_14681_));
 sky130_fd_sc_hd__nand2_4 _45232_ (.A(_14679_),
    .B(_14681_),
    .Y(_14682_));
 sky130_fd_sc_hd__nand2_4 _45233_ (.A(_12308_),
    .B(_12523_),
    .Y(_14683_));
 sky130_fd_sc_hd__nand2_4 _45234_ (.A(_12310_),
    .B(_07051_),
    .Y(_14684_));
 sky130_fd_sc_hd__nand2_4 _45235_ (.A(_14683_),
    .B(_14684_),
    .Y(_14685_));
 sky130_fd_sc_hd__nand4_4 _45236_ (.A(_11989_),
    .B(_11991_),
    .C(_12527_),
    .D(_12528_),
    .Y(_14686_));
 sky130_fd_sc_hd__nand2_4 _45237_ (.A(_12315_),
    .B(_03511_),
    .Y(_14687_));
 sky130_vsdinv _45238_ (.A(_14687_),
    .Y(_14688_));
 sky130_fd_sc_hd__a21o_4 _45239_ (.A1(_14685_),
    .A2(_14686_),
    .B1(_14688_),
    .X(_14689_));
 sky130_fd_sc_hd__buf_1 _45240_ (.A(_14688_),
    .X(_14690_));
 sky130_fd_sc_hd__nand3_4 _45241_ (.A(_14685_),
    .B(_14686_),
    .C(_14690_),
    .Y(_14691_));
 sky130_fd_sc_hd__a21boi_4 _45242_ (.A1(_14446_),
    .A2(_14449_),
    .B1_N(_14447_),
    .Y(_14692_));
 sky130_fd_sc_hd__a21boi_4 _45243_ (.A1(_14689_),
    .A2(_14691_),
    .B1_N(_14692_),
    .Y(_14693_));
 sky130_fd_sc_hd__nand2_4 _45244_ (.A(_14689_),
    .B(_14691_),
    .Y(_14694_));
 sky130_fd_sc_hd__nor2_4 _45245_ (.A(_14692_),
    .B(_14694_),
    .Y(_14695_));
 sky130_fd_sc_hd__o21a_4 _45246_ (.A1(_14693_),
    .A2(_14695_),
    .B1(_14461_),
    .X(_14696_));
 sky130_fd_sc_hd__or3_4 _45247_ (.A(_14461_),
    .B(_14693_),
    .C(_14695_),
    .X(_14697_));
 sky130_vsdinv _45248_ (.A(_14697_),
    .Y(_14698_));
 sky130_fd_sc_hd__nor2_4 _45249_ (.A(_14696_),
    .B(_14698_),
    .Y(_14699_));
 sky130_vsdinv _45250_ (.A(_14699_),
    .Y(_14700_));
 sky130_fd_sc_hd__nand2_4 _45251_ (.A(_14682_),
    .B(_14700_),
    .Y(_14701_));
 sky130_fd_sc_hd__nand3_4 _45252_ (.A(_14679_),
    .B(_14699_),
    .C(_14681_),
    .Y(_14702_));
 sky130_fd_sc_hd__nand2_4 _45253_ (.A(_14701_),
    .B(_14702_),
    .Y(_14703_));
 sky130_fd_sc_hd__a21boi_4 _45254_ (.A1(_14401_),
    .A2(_14404_),
    .B1_N(_14402_),
    .Y(_14704_));
 sky130_fd_sc_hd__nand2_4 _45255_ (.A(_14703_),
    .B(_14704_),
    .Y(_14705_));
 sky130_vsdinv _45256_ (.A(_14704_),
    .Y(_14706_));
 sky130_fd_sc_hd__nand3_4 _45257_ (.A(_14706_),
    .B(_14701_),
    .C(_14702_),
    .Y(_14707_));
 sky130_fd_sc_hd__buf_1 _45258_ (.A(_14707_),
    .X(_14708_));
 sky130_fd_sc_hd__nand2_4 _45259_ (.A(_14705_),
    .B(_14708_),
    .Y(_14709_));
 sky130_fd_sc_hd__a21boi_4 _45260_ (.A1(_14440_),
    .A2(_14468_),
    .B1_N(_14442_),
    .Y(_14710_));
 sky130_fd_sc_hd__nand2_4 _45261_ (.A(_14709_),
    .B(_14710_),
    .Y(_14711_));
 sky130_vsdinv _45262_ (.A(_14710_),
    .Y(_14712_));
 sky130_fd_sc_hd__nand3_4 _45263_ (.A(_14705_),
    .B(_14712_),
    .C(_14707_),
    .Y(_14713_));
 sky130_fd_sc_hd__nand2_4 _45264_ (.A(_14711_),
    .B(_14713_),
    .Y(_14714_));
 sky130_fd_sc_hd__nand2_4 _45265_ (.A(_14658_),
    .B(_14714_),
    .Y(_14715_));
 sky130_fd_sc_hd__a21oi_4 _45266_ (.A1(_14705_),
    .A2(_14708_),
    .B1(_14712_),
    .Y(_14716_));
 sky130_vsdinv _45267_ (.A(_14713_),
    .Y(_14717_));
 sky130_fd_sc_hd__nor2_4 _45268_ (.A(_14716_),
    .B(_14717_),
    .Y(_14718_));
 sky130_fd_sc_hd__nand3_4 _45269_ (.A(_14718_),
    .B(_14657_),
    .C(_14655_),
    .Y(_14719_));
 sky130_fd_sc_hd__nand2_4 _45270_ (.A(_14715_),
    .B(_14719_),
    .Y(_14720_));
 sky130_fd_sc_hd__a21boi_4 _45271_ (.A1(_14484_),
    .A2(_14416_),
    .B1_N(_14418_),
    .Y(_14721_));
 sky130_fd_sc_hd__nand2_4 _45272_ (.A(_14720_),
    .B(_14721_),
    .Y(_14722_));
 sky130_vsdinv _45273_ (.A(_14721_),
    .Y(_14723_));
 sky130_fd_sc_hd__nand3_4 _45274_ (.A(_14723_),
    .B(_14715_),
    .C(_14719_),
    .Y(_14724_));
 sky130_fd_sc_hd__nand2_4 _45275_ (.A(_14722_),
    .B(_14724_),
    .Y(_14725_));
 sky130_fd_sc_hd__o21a_4 _45276_ (.A1(_13926_),
    .A2(_14456_),
    .B1(_14458_),
    .X(_14726_));
 sky130_vsdinv _45277_ (.A(_14726_),
    .Y(_14727_));
 sky130_fd_sc_hd__nand3_4 _45278_ (.A(_14727_),
    .B(_13992_),
    .C(_13991_),
    .Y(_14728_));
 sky130_fd_sc_hd__nand2_4 _45279_ (.A(_13718_),
    .B(_14726_),
    .Y(_14729_));
 sky130_fd_sc_hd__a21o_4 _45280_ (.A1(_14728_),
    .A2(_14729_),
    .B1(_13997_),
    .X(_14730_));
 sky130_fd_sc_hd__nand3_4 _45281_ (.A(_14728_),
    .B(_14729_),
    .C(_14248_),
    .Y(_14731_));
 sky130_fd_sc_hd__nand2_4 _45282_ (.A(_14730_),
    .B(_14731_),
    .Y(_14732_));
 sky130_vsdinv _45283_ (.A(_14732_),
    .Y(_14733_));
 sky130_fd_sc_hd__o21ai_4 _45284_ (.A1(_14453_),
    .A2(_14467_),
    .B1(_14733_),
    .Y(_14734_));
 sky130_fd_sc_hd__buf_1 _45285_ (.A(_14732_),
    .X(_14735_));
 sky130_fd_sc_hd__a21oi_4 _45286_ (.A1(_14464_),
    .A2(_14455_),
    .B1(_14453_),
    .Y(_14736_));
 sky130_fd_sc_hd__nand2_4 _45287_ (.A(_14735_),
    .B(_14736_),
    .Y(_14737_));
 sky130_fd_sc_hd__a21boi_4 _45288_ (.A1(_14496_),
    .A2(_14499_),
    .B1_N(_14498_),
    .Y(_14738_));
 sky130_vsdinv _45289_ (.A(_14738_),
    .Y(_14739_));
 sky130_fd_sc_hd__a21o_4 _45290_ (.A1(_14734_),
    .A2(_14737_),
    .B1(_14739_),
    .X(_14740_));
 sky130_fd_sc_hd__nand3_4 _45291_ (.A(_14734_),
    .B(_14737_),
    .C(_14739_),
    .Y(_14741_));
 sky130_fd_sc_hd__nand2_4 _45292_ (.A(_14740_),
    .B(_14741_),
    .Y(_14742_));
 sky130_fd_sc_hd__maj3_4 _45293_ (.A(_14505_),
    .B(_14503_),
    .C(_14493_),
    .X(_14743_));
 sky130_fd_sc_hd__nand2_4 _45294_ (.A(_14742_),
    .B(_14743_),
    .Y(_14744_));
 sky130_vsdinv _45295_ (.A(_14743_),
    .Y(_14745_));
 sky130_fd_sc_hd__nand3_4 _45296_ (.A(_14740_),
    .B(_14745_),
    .C(_14741_),
    .Y(_14746_));
 sky130_fd_sc_hd__nand2_4 _45297_ (.A(_14744_),
    .B(_14746_),
    .Y(_14747_));
 sky130_fd_sc_hd__nand2_4 _45298_ (.A(_14747_),
    .B(_13480_),
    .Y(_14748_));
 sky130_fd_sc_hd__nand3_4 _45299_ (.A(_14744_),
    .B(_13483_),
    .C(_14746_),
    .Y(_14749_));
 sky130_fd_sc_hd__nand2_4 _45300_ (.A(_14748_),
    .B(_14749_),
    .Y(_14750_));
 sky130_fd_sc_hd__a21boi_4 _45301_ (.A1(_14474_),
    .A2(_14477_),
    .B1_N(_14475_),
    .Y(_14751_));
 sky130_fd_sc_hd__nand2_4 _45302_ (.A(_14750_),
    .B(_14751_),
    .Y(_14752_));
 sky130_vsdinv _45303_ (.A(_14751_),
    .Y(_14753_));
 sky130_fd_sc_hd__nand3_4 _45304_ (.A(_14753_),
    .B(_14748_),
    .C(_14749_),
    .Y(_14754_));
 sky130_fd_sc_hd__buf_1 _45305_ (.A(_14754_),
    .X(_14755_));
 sky130_fd_sc_hd__nand2_4 _45306_ (.A(_14752_),
    .B(_14755_),
    .Y(_14756_));
 sky130_fd_sc_hd__buf_1 _45307_ (.A(_14015_),
    .X(_14757_));
 sky130_fd_sc_hd__a21boi_4 _45308_ (.A1(_14511_),
    .A2(_14757_),
    .B1_N(_14513_),
    .Y(_14758_));
 sky130_fd_sc_hd__nand2_4 _45309_ (.A(_14756_),
    .B(_14758_),
    .Y(_14759_));
 sky130_vsdinv _45310_ (.A(_14758_),
    .Y(_14760_));
 sky130_fd_sc_hd__nand3_4 _45311_ (.A(_14752_),
    .B(_14760_),
    .C(_14754_),
    .Y(_14761_));
 sky130_fd_sc_hd__nand2_4 _45312_ (.A(_14759_),
    .B(_14761_),
    .Y(_14762_));
 sky130_fd_sc_hd__nand2_4 _45313_ (.A(_14725_),
    .B(_14762_),
    .Y(_14763_));
 sky130_fd_sc_hd__a21oi_4 _45314_ (.A1(_14752_),
    .A2(_14755_),
    .B1(_14760_),
    .Y(_14764_));
 sky130_vsdinv _45315_ (.A(_14761_),
    .Y(_14765_));
 sky130_fd_sc_hd__nor2_4 _45316_ (.A(_14764_),
    .B(_14765_),
    .Y(_14766_));
 sky130_fd_sc_hd__nand3_4 _45317_ (.A(_14766_),
    .B(_14722_),
    .C(_14724_),
    .Y(_14767_));
 sky130_fd_sc_hd__nand2_4 _45318_ (.A(_14763_),
    .B(_14767_),
    .Y(_14768_));
 sky130_fd_sc_hd__a21boi_4 _45319_ (.A1(_14531_),
    .A2(_14488_),
    .B1_N(_14491_),
    .Y(_14769_));
 sky130_fd_sc_hd__nand2_4 _45320_ (.A(_14768_),
    .B(_14769_),
    .Y(_14770_));
 sky130_vsdinv _45321_ (.A(_14769_),
    .Y(_14771_));
 sky130_fd_sc_hd__nand3_4 _45322_ (.A(_14771_),
    .B(_14763_),
    .C(_14767_),
    .Y(_14772_));
 sky130_fd_sc_hd__nand2_4 _45323_ (.A(_14770_),
    .B(_14772_),
    .Y(_14773_));
 sky130_fd_sc_hd__a21boi_4 _45324_ (.A1(_14519_),
    .A2(_14524_),
    .B1_N(_14522_),
    .Y(_14774_));
 sky130_fd_sc_hd__xor2_4 _45325_ (.A(_14291_),
    .B(_14774_),
    .X(_14775_));
 sky130_fd_sc_hd__nand2_4 _45326_ (.A(_14773_),
    .B(_14775_),
    .Y(_14776_));
 sky130_vsdinv _45327_ (.A(_14775_),
    .Y(_14777_));
 sky130_fd_sc_hd__nand3_4 _45328_ (.A(_14770_),
    .B(_14772_),
    .C(_14777_),
    .Y(_14778_));
 sky130_fd_sc_hd__nand2_4 _45329_ (.A(_14776_),
    .B(_14778_),
    .Y(_14779_));
 sky130_fd_sc_hd__a21boi_4 _45330_ (.A1(_14535_),
    .A2(_14543_),
    .B1_N(_14538_),
    .Y(_14780_));
 sky130_fd_sc_hd__nand2_4 _45331_ (.A(_14779_),
    .B(_14780_),
    .Y(_14781_));
 sky130_vsdinv _45332_ (.A(_14780_),
    .Y(_14782_));
 sky130_fd_sc_hd__nand3_4 _45333_ (.A(_14782_),
    .B(_14778_),
    .C(_14776_),
    .Y(_14783_));
 sky130_fd_sc_hd__nand2_4 _45334_ (.A(_14781_),
    .B(_14783_),
    .Y(_14784_));
 sky130_fd_sc_hd__a21oi_4 _45335_ (.A1(_14277_),
    .A2(_14271_),
    .B1(_14050_),
    .Y(_14785_));
 sky130_vsdinv _45336_ (.A(_14785_),
    .Y(_14786_));
 sky130_fd_sc_hd__nand2_4 _45337_ (.A(_14784_),
    .B(_14786_),
    .Y(_14787_));
 sky130_fd_sc_hd__nand3_4 _45338_ (.A(_14781_),
    .B(_14785_),
    .C(_14783_),
    .Y(_14788_));
 sky130_fd_sc_hd__nand2_4 _45339_ (.A(_14787_),
    .B(_14788_),
    .Y(_14789_));
 sky130_fd_sc_hd__a21boi_4 _45340_ (.A1(_14547_),
    .A2(_14551_),
    .B1_N(_14549_),
    .Y(_14790_));
 sky130_fd_sc_hd__nand2_4 _45341_ (.A(_14789_),
    .B(_14790_),
    .Y(_14791_));
 sky130_vsdinv _45342_ (.A(_14790_),
    .Y(_14792_));
 sky130_fd_sc_hd__nand3_4 _45343_ (.A(_14792_),
    .B(_14787_),
    .C(_14788_),
    .Y(_14793_));
 sky130_fd_sc_hd__nand2_4 _45344_ (.A(_14791_),
    .B(_14793_),
    .Y(_14794_));
 sky130_fd_sc_hd__nand4_4 _45345_ (.A(_14312_),
    .B(_14310_),
    .C(_14557_),
    .D(_14559_),
    .Y(_14795_));
 sky130_fd_sc_hd__a21boi_4 _45346_ (.A1(_14561_),
    .A2(_14557_),
    .B1_N(_14559_),
    .Y(_14796_));
 sky130_fd_sc_hd__o21ai_4 _45347_ (.A1(_14317_),
    .A2(_14795_),
    .B1(_14796_),
    .Y(_14797_));
 sky130_vsdinv _45348_ (.A(_14795_),
    .Y(_14798_));
 sky130_fd_sc_hd__nand2_4 _45349_ (.A(_14314_),
    .B(_14798_),
    .Y(_14799_));
 sky130_fd_sc_hd__nor2_4 _45350_ (.A(_14799_),
    .B(_13805_),
    .Y(_14800_));
 sky130_fd_sc_hd__or2_4 _45351_ (.A(_14797_),
    .B(_14800_),
    .X(_14801_));
 sky130_fd_sc_hd__buf_1 _45352_ (.A(_14801_),
    .X(_14802_));
 sky130_fd_sc_hd__xnor2_4 _45353_ (.A(_14794_),
    .B(_14802_),
    .Y(_01449_));
 sky130_fd_sc_hd__a21oi_4 _45354_ (.A1(_14610_),
    .A2(_14612_),
    .B1(_14616_),
    .Y(_14803_));
 sky130_fd_sc_hd__o21ai_4 _45355_ (.A1(_14650_),
    .A2(_14803_),
    .B1(_14617_),
    .Y(_14804_));
 sky130_vsdinv _45356_ (.A(_14804_),
    .Y(_14805_));
 sky130_fd_sc_hd__a21boi_4 _45357_ (.A1(_14564_),
    .A2(_14568_),
    .B1_N(_14566_),
    .Y(_14806_));
 sky130_vsdinv _45358_ (.A(_14806_),
    .Y(_14807_));
 sky130_fd_sc_hd__nand2_4 _45359_ (.A(_13825_),
    .B(_11433_),
    .Y(_14808_));
 sky130_fd_sc_hd__o21ai_4 _45360_ (.A1(_08971_),
    .A2(_11432_),
    .B1(_14808_),
    .Y(_14809_));
 sky130_fd_sc_hd__nand2_4 _45361_ (.A(_07432_),
    .B(_10516_),
    .Y(_14810_));
 sky130_vsdinv _45362_ (.A(_14810_),
    .Y(_14811_));
 sky130_fd_sc_hd__nand4_4 _45363_ (.A(_03311_),
    .B(_10989_),
    .C(_10959_),
    .D(_14565_),
    .Y(_14812_));
 sky130_fd_sc_hd__nand3_4 _45364_ (.A(_14809_),
    .B(_14811_),
    .C(_14812_),
    .Y(_14813_));
 sky130_fd_sc_hd__nand2_4 _45365_ (.A(_14809_),
    .B(_14812_),
    .Y(_14814_));
 sky130_fd_sc_hd__nand2_4 _45366_ (.A(_14814_),
    .B(_14810_),
    .Y(_14815_));
 sky130_fd_sc_hd__nand3_4 _45367_ (.A(_14807_),
    .B(_14813_),
    .C(_14815_),
    .Y(_14816_));
 sky130_fd_sc_hd__nand2_4 _45368_ (.A(_14815_),
    .B(_14813_),
    .Y(_14817_));
 sky130_fd_sc_hd__nand2_4 _45369_ (.A(_14817_),
    .B(_14806_),
    .Y(_14818_));
 sky130_fd_sc_hd__nand2_4 _45370_ (.A(_14816_),
    .B(_14818_),
    .Y(_14819_));
 sky130_fd_sc_hd__nand2_4 _45371_ (.A(_13331_),
    .B(_10506_),
    .Y(_14820_));
 sky130_fd_sc_hd__nand2_4 _45372_ (.A(_07875_),
    .B(_10505_),
    .Y(_14821_));
 sky130_fd_sc_hd__nand2_4 _45373_ (.A(_14820_),
    .B(_14821_),
    .Y(_14822_));
 sky130_fd_sc_hd__nand4_4 _45374_ (.A(_13331_),
    .B(_11010_),
    .C(_10505_),
    .D(_10506_),
    .Y(_14823_));
 sky130_fd_sc_hd__nand2_4 _45375_ (.A(_03337_),
    .B(_12095_),
    .Y(_14824_));
 sky130_vsdinv _45376_ (.A(_14824_),
    .Y(_14825_));
 sky130_fd_sc_hd__a21oi_4 _45377_ (.A1(_14822_),
    .A2(_14823_),
    .B1(_14825_),
    .Y(_14826_));
 sky130_fd_sc_hd__nand3_4 _45378_ (.A(_14822_),
    .B(_14823_),
    .C(_14825_),
    .Y(_14827_));
 sky130_vsdinv _45379_ (.A(_14827_),
    .Y(_14828_));
 sky130_fd_sc_hd__nor2_4 _45380_ (.A(_14826_),
    .B(_14828_),
    .Y(_14829_));
 sky130_vsdinv _45381_ (.A(_14829_),
    .Y(_14830_));
 sky130_fd_sc_hd__nand2_4 _45382_ (.A(_14819_),
    .B(_14830_),
    .Y(_14831_));
 sky130_fd_sc_hd__nand3_4 _45383_ (.A(_14816_),
    .B(_14818_),
    .C(_14829_),
    .Y(_14832_));
 sky130_fd_sc_hd__nand2_4 _45384_ (.A(_14831_),
    .B(_14832_),
    .Y(_14833_));
 sky130_fd_sc_hd__a21boi_4 _45385_ (.A1(_14573_),
    .A2(_14582_),
    .B1_N(_14575_),
    .Y(_14834_));
 sky130_fd_sc_hd__nand2_4 _45386_ (.A(_14833_),
    .B(_14834_),
    .Y(_14835_));
 sky130_fd_sc_hd__nand2_4 _45387_ (.A(_14584_),
    .B(_14575_),
    .Y(_14836_));
 sky130_fd_sc_hd__nand3_4 _45388_ (.A(_14836_),
    .B(_14832_),
    .C(_14831_),
    .Y(_14837_));
 sky130_fd_sc_hd__nand2_4 _45389_ (.A(_14835_),
    .B(_14837_),
    .Y(_14838_));
 sky130_vsdinv _45390_ (.A(_14576_),
    .Y(_14839_));
 sky130_fd_sc_hd__a21boi_4 _45391_ (.A1(_14579_),
    .A2(_14839_),
    .B1_N(_14580_),
    .Y(_14840_));
 sky130_fd_sc_hd__nand2_4 _45392_ (.A(_10619_),
    .B(_11793_),
    .Y(_14841_));
 sky130_fd_sc_hd__nand2_4 _45393_ (.A(_08056_),
    .B(_13011_),
    .Y(_14842_));
 sky130_fd_sc_hd__nand2_4 _45394_ (.A(_14841_),
    .B(_14842_),
    .Y(_14843_));
 sky130_fd_sc_hd__nand4_4 _45395_ (.A(_03342_),
    .B(_10625_),
    .C(_11797_),
    .D(_11142_),
    .Y(_14844_));
 sky130_fd_sc_hd__nand2_4 _45396_ (.A(_13342_),
    .B(_09347_),
    .Y(_14845_));
 sky130_vsdinv _45397_ (.A(_14845_),
    .Y(_14846_));
 sky130_fd_sc_hd__a21o_4 _45398_ (.A1(_14843_),
    .A2(_14844_),
    .B1(_14846_),
    .X(_14847_));
 sky130_fd_sc_hd__nand3_4 _45399_ (.A(_14843_),
    .B(_14844_),
    .C(_14846_),
    .Y(_14848_));
 sky130_fd_sc_hd__nand2_4 _45400_ (.A(_14847_),
    .B(_14848_),
    .Y(_14849_));
 sky130_fd_sc_hd__or2_4 _45401_ (.A(_14840_),
    .B(_14849_),
    .X(_14850_));
 sky130_fd_sc_hd__nand2_4 _45402_ (.A(_14849_),
    .B(_14840_),
    .Y(_14851_));
 sky130_fd_sc_hd__a21boi_4 _45403_ (.A1(_14593_),
    .A2(_14596_),
    .B1_N(_14594_),
    .Y(_14852_));
 sky130_vsdinv _45404_ (.A(_14852_),
    .Y(_14853_));
 sky130_fd_sc_hd__a21oi_4 _45405_ (.A1(_14850_),
    .A2(_14851_),
    .B1(_14853_),
    .Y(_14854_));
 sky130_vsdinv _45406_ (.A(_14854_),
    .Y(_14855_));
 sky130_fd_sc_hd__nand3_4 _45407_ (.A(_14850_),
    .B(_14853_),
    .C(_14851_),
    .Y(_14856_));
 sky130_fd_sc_hd__nand2_4 _45408_ (.A(_14855_),
    .B(_14856_),
    .Y(_14857_));
 sky130_fd_sc_hd__nand2_4 _45409_ (.A(_14838_),
    .B(_14857_),
    .Y(_14858_));
 sky130_fd_sc_hd__nand4_4 _45410_ (.A(_14856_),
    .B(_14835_),
    .C(_14855_),
    .D(_14837_),
    .Y(_14859_));
 sky130_fd_sc_hd__nand2_4 _45411_ (.A(_14858_),
    .B(_14859_),
    .Y(_14860_));
 sky130_fd_sc_hd__a21boi_4 _45412_ (.A1(_14611_),
    .A2(_14587_),
    .B1_N(_14589_),
    .Y(_14861_));
 sky130_fd_sc_hd__nand2_4 _45413_ (.A(_14860_),
    .B(_14861_),
    .Y(_14862_));
 sky130_fd_sc_hd__a21oi_4 _45414_ (.A1(_14583_),
    .A2(_14584_),
    .B1(_14588_),
    .Y(_14863_));
 sky130_fd_sc_hd__o21ai_4 _45415_ (.A1(_14609_),
    .A2(_14863_),
    .B1(_14589_),
    .Y(_14864_));
 sky130_fd_sc_hd__nand3_4 _45416_ (.A(_14864_),
    .B(_14859_),
    .C(_14858_),
    .Y(_14865_));
 sky130_fd_sc_hd__nand2_4 _45417_ (.A(_14862_),
    .B(_14865_),
    .Y(_14866_));
 sky130_fd_sc_hd__buf_1 _45418_ (.A(_11824_),
    .X(_14867_));
 sky130_fd_sc_hd__nand2_4 _45419_ (.A(_08756_),
    .B(_14867_),
    .Y(_14868_));
 sky130_fd_sc_hd__buf_1 _45420_ (.A(_11829_),
    .X(_14869_));
 sky130_fd_sc_hd__nand2_4 _45421_ (.A(_14137_),
    .B(_14869_),
    .Y(_14870_));
 sky130_fd_sc_hd__nand2_4 _45422_ (.A(_14868_),
    .B(_14870_),
    .Y(_14871_));
 sky130_fd_sc_hd__buf_1 _45423_ (.A(_10884_),
    .X(_14872_));
 sky130_fd_sc_hd__buf_1 _45424_ (.A(_12157_),
    .X(_14873_));
 sky130_fd_sc_hd__nand4_4 _45425_ (.A(_08756_),
    .B(_14137_),
    .C(_14872_),
    .D(_14873_),
    .Y(_14874_));
 sky130_fd_sc_hd__nand2_4 _45426_ (.A(_13943_),
    .B(_13872_),
    .Y(_14875_));
 sky130_vsdinv _45427_ (.A(_14875_),
    .Y(_14876_));
 sky130_fd_sc_hd__a21o_4 _45428_ (.A1(_14871_),
    .A2(_14874_),
    .B1(_14876_),
    .X(_14877_));
 sky130_fd_sc_hd__nand3_4 _45429_ (.A(_14871_),
    .B(_14874_),
    .C(_14876_),
    .Y(_14878_));
 sky130_fd_sc_hd__nand2_4 _45430_ (.A(_14877_),
    .B(_14878_),
    .Y(_14879_));
 sky130_fd_sc_hd__a21o_4 _45431_ (.A1(_14622_),
    .A2(_14626_),
    .B1(_14879_),
    .X(_14880_));
 sky130_fd_sc_hd__nand3_4 _45432_ (.A(_14879_),
    .B(_14622_),
    .C(_14626_),
    .Y(_14881_));
 sky130_fd_sc_hd__buf_1 _45433_ (.A(_11317_),
    .X(_14882_));
 sky130_fd_sc_hd__nand2_4 _45434_ (.A(_14882_),
    .B(_03546_),
    .Y(_14883_));
 sky130_fd_sc_hd__buf_1 _45435_ (.A(_09580_),
    .X(_14884_));
 sky130_fd_sc_hd__nand2_4 _45436_ (.A(_14884_),
    .B(_13611_),
    .Y(_14885_));
 sky130_fd_sc_hd__o21ai_4 _45437_ (.A1(_03377_),
    .A2(_03559_),
    .B1(_14885_),
    .Y(_14886_));
 sky130_fd_sc_hd__nand4_4 _45438_ (.A(_12824_),
    .B(_13117_),
    .C(_13884_),
    .D(_13885_),
    .Y(_14887_));
 sky130_fd_sc_hd__nand2_4 _45439_ (.A(_14886_),
    .B(_14887_),
    .Y(_14888_));
 sky130_fd_sc_hd__xor2_4 _45440_ (.A(_14883_),
    .B(_14888_),
    .X(_14889_));
 sky130_fd_sc_hd__a21o_4 _45441_ (.A1(_14880_),
    .A2(_14881_),
    .B1(_14889_),
    .X(_14890_));
 sky130_fd_sc_hd__nand3_4 _45442_ (.A(_14880_),
    .B(_14889_),
    .C(_14881_),
    .Y(_14891_));
 sky130_fd_sc_hd__o21a_4 _45443_ (.A1(_14604_),
    .A2(_14600_),
    .B1(_14603_),
    .X(_14892_));
 sky130_vsdinv _45444_ (.A(_14892_),
    .Y(_14893_));
 sky130_fd_sc_hd__a21o_4 _45445_ (.A1(_14890_),
    .A2(_14891_),
    .B1(_14893_),
    .X(_14894_));
 sky130_fd_sc_hd__nand3_4 _45446_ (.A(_14890_),
    .B(_14893_),
    .C(_14891_),
    .Y(_14895_));
 sky130_fd_sc_hd__a21boi_4 _45447_ (.A1(_14636_),
    .A2(_14629_),
    .B1_N(_14628_),
    .Y(_14896_));
 sky130_vsdinv _45448_ (.A(_14896_),
    .Y(_14897_));
 sky130_fd_sc_hd__a21o_4 _45449_ (.A1(_14894_),
    .A2(_14895_),
    .B1(_14897_),
    .X(_14898_));
 sky130_fd_sc_hd__nand3_4 _45450_ (.A(_14894_),
    .B(_14897_),
    .C(_14895_),
    .Y(_14899_));
 sky130_fd_sc_hd__nand2_4 _45451_ (.A(_14898_),
    .B(_14899_),
    .Y(_14900_));
 sky130_fd_sc_hd__nand2_4 _45452_ (.A(_14866_),
    .B(_14900_),
    .Y(_14901_));
 sky130_fd_sc_hd__nand4_4 _45453_ (.A(_14899_),
    .B(_14862_),
    .C(_14865_),
    .D(_14898_),
    .Y(_14902_));
 sky130_fd_sc_hd__nand2_4 _45454_ (.A(_14901_),
    .B(_14902_),
    .Y(_14903_));
 sky130_fd_sc_hd__nand2_4 _45455_ (.A(_14805_),
    .B(_14903_),
    .Y(_14904_));
 sky130_fd_sc_hd__nand3_4 _45456_ (.A(_14804_),
    .B(_14902_),
    .C(_14901_),
    .Y(_14905_));
 sky130_fd_sc_hd__nand2_4 _45457_ (.A(_14904_),
    .B(_14905_),
    .Y(_14906_));
 sky130_fd_sc_hd__maj3_4 _45458_ (.A(_14631_),
    .B(_14632_),
    .C(_14630_),
    .X(_14907_));
 sky130_fd_sc_hd__nand2_4 _45459_ (.A(_10087_),
    .B(_08358_),
    .Y(_14908_));
 sky130_fd_sc_hd__nand2_4 _45460_ (.A(_11323_),
    .B(_08357_),
    .Y(_14909_));
 sky130_fd_sc_hd__nand2_4 _45461_ (.A(_14908_),
    .B(_14909_),
    .Y(_14910_));
 sky130_fd_sc_hd__nand4_4 _45462_ (.A(_13128_),
    .B(_10843_),
    .C(_07920_),
    .D(_07923_),
    .Y(_14911_));
 sky130_fd_sc_hd__nand2_4 _45463_ (.A(_11334_),
    .B(_07720_),
    .Y(_14912_));
 sky130_vsdinv _45464_ (.A(_14912_),
    .Y(_14913_));
 sky130_fd_sc_hd__a21o_4 _45465_ (.A1(_14910_),
    .A2(_14911_),
    .B1(_14913_),
    .X(_14914_));
 sky130_fd_sc_hd__nand3_4 _45466_ (.A(_14910_),
    .B(_14911_),
    .C(_14913_),
    .Y(_14915_));
 sky130_fd_sc_hd__nand2_4 _45467_ (.A(_14914_),
    .B(_14915_),
    .Y(_14916_));
 sky130_fd_sc_hd__or2_4 _45468_ (.A(_14907_),
    .B(_14916_),
    .X(_14917_));
 sky130_fd_sc_hd__nand2_4 _45469_ (.A(_14916_),
    .B(_14907_),
    .Y(_14918_));
 sky130_fd_sc_hd__a21boi_4 _45470_ (.A1(_14661_),
    .A2(_14664_),
    .B1_N(_14662_),
    .Y(_14919_));
 sky130_vsdinv _45471_ (.A(_14919_),
    .Y(_14920_));
 sky130_fd_sc_hd__a21o_4 _45472_ (.A1(_14917_),
    .A2(_14918_),
    .B1(_14920_),
    .X(_14921_));
 sky130_fd_sc_hd__nand3_4 _45473_ (.A(_14917_),
    .B(_14920_),
    .C(_14918_),
    .Y(_14922_));
 sky130_fd_sc_hd__nand2_4 _45474_ (.A(_14921_),
    .B(_14922_),
    .Y(_14923_));
 sky130_fd_sc_hd__o21a_4 _45475_ (.A1(_14675_),
    .A2(_14669_),
    .B1(_14672_),
    .X(_14924_));
 sky130_fd_sc_hd__nand2_4 _45476_ (.A(_14923_),
    .B(_14924_),
    .Y(_14925_));
 sky130_vsdinv _45477_ (.A(_14924_),
    .Y(_14926_));
 sky130_fd_sc_hd__nand3_4 _45478_ (.A(_14921_),
    .B(_14922_),
    .C(_14926_),
    .Y(_14927_));
 sky130_fd_sc_hd__nand2_4 _45479_ (.A(_14925_),
    .B(_14927_),
    .Y(_14928_));
 sky130_fd_sc_hd__a21boi_4 _45480_ (.A1(_14685_),
    .A2(_14690_),
    .B1_N(_14686_),
    .Y(_14929_));
 sky130_fd_sc_hd__nand2_4 _45481_ (.A(_11687_),
    .B(_07059_),
    .Y(_14930_));
 sky130_fd_sc_hd__o21ai_4 _45482_ (.A1(_03400_),
    .A2(_03526_),
    .B1(_14930_),
    .Y(_14931_));
 sky130_fd_sc_hd__nand4_4 _45483_ (.A(_11690_),
    .B(_12909_),
    .C(_12527_),
    .D(_12528_),
    .Y(_14932_));
 sky130_fd_sc_hd__a21o_4 _45484_ (.A1(_14931_),
    .A2(_14932_),
    .B1(_14688_),
    .X(_14933_));
 sky130_fd_sc_hd__nand3_4 _45485_ (.A(_14931_),
    .B(_14690_),
    .C(_14932_),
    .Y(_14934_));
 sky130_fd_sc_hd__nand2_4 _45486_ (.A(_14933_),
    .B(_14934_),
    .Y(_14935_));
 sky130_fd_sc_hd__nor2_4 _45487_ (.A(_14929_),
    .B(_14935_),
    .Y(_14936_));
 sky130_vsdinv _45488_ (.A(_14936_),
    .Y(_14937_));
 sky130_fd_sc_hd__nand2_4 _45489_ (.A(_14935_),
    .B(_14929_),
    .Y(_14938_));
 sky130_fd_sc_hd__a21oi_4 _45490_ (.A1(_14937_),
    .A2(_14938_),
    .B1(_14463_),
    .Y(_14939_));
 sky130_fd_sc_hd__nand3_4 _45491_ (.A(_14937_),
    .B(_14462_),
    .C(_14938_),
    .Y(_14940_));
 sky130_vsdinv _45492_ (.A(_14940_),
    .Y(_14941_));
 sky130_fd_sc_hd__nor2_4 _45493_ (.A(_14939_),
    .B(_14941_),
    .Y(_14942_));
 sky130_vsdinv _45494_ (.A(_14942_),
    .Y(_14943_));
 sky130_fd_sc_hd__nand2_4 _45495_ (.A(_14928_),
    .B(_14943_),
    .Y(_14944_));
 sky130_fd_sc_hd__nand3_4 _45496_ (.A(_14925_),
    .B(_14942_),
    .C(_14927_),
    .Y(_14945_));
 sky130_fd_sc_hd__nand2_4 _45497_ (.A(_14944_),
    .B(_14945_),
    .Y(_14946_));
 sky130_fd_sc_hd__o21ai_4 _45498_ (.A1(_14645_),
    .A2(_14641_),
    .B1(_14642_),
    .Y(_14947_));
 sky130_vsdinv _45499_ (.A(_14947_),
    .Y(_14948_));
 sky130_fd_sc_hd__nand2_4 _45500_ (.A(_14946_),
    .B(_14948_),
    .Y(_14949_));
 sky130_fd_sc_hd__nand3_4 _45501_ (.A(_14944_),
    .B(_14947_),
    .C(_14945_),
    .Y(_14950_));
 sky130_fd_sc_hd__a21boi_4 _45502_ (.A1(_14679_),
    .A2(_14699_),
    .B1_N(_14681_),
    .Y(_14951_));
 sky130_vsdinv _45503_ (.A(_14951_),
    .Y(_14952_));
 sky130_fd_sc_hd__a21oi_4 _45504_ (.A1(_14949_),
    .A2(_14950_),
    .B1(_14952_),
    .Y(_14953_));
 sky130_vsdinv _45505_ (.A(_14953_),
    .Y(_14954_));
 sky130_fd_sc_hd__nand3_4 _45506_ (.A(_14949_),
    .B(_14952_),
    .C(_14950_),
    .Y(_14955_));
 sky130_fd_sc_hd__nand2_4 _45507_ (.A(_14954_),
    .B(_14955_),
    .Y(_14956_));
 sky130_fd_sc_hd__nand2_4 _45508_ (.A(_14906_),
    .B(_14956_),
    .Y(_14957_));
 sky130_vsdinv _45509_ (.A(_14955_),
    .Y(_14958_));
 sky130_fd_sc_hd__nor2_4 _45510_ (.A(_14953_),
    .B(_14958_),
    .Y(_14959_));
 sky130_fd_sc_hd__nand3_4 _45511_ (.A(_14959_),
    .B(_14905_),
    .C(_14904_),
    .Y(_14960_));
 sky130_fd_sc_hd__nand2_4 _45512_ (.A(_14957_),
    .B(_14960_),
    .Y(_14961_));
 sky130_fd_sc_hd__a21boi_4 _45513_ (.A1(_14718_),
    .A2(_14655_),
    .B1_N(_14657_),
    .Y(_14962_));
 sky130_fd_sc_hd__nand2_4 _45514_ (.A(_14961_),
    .B(_14962_),
    .Y(_14963_));
 sky130_fd_sc_hd__a21boi_4 _45515_ (.A1(_14651_),
    .A2(_14652_),
    .B1_N(_14654_),
    .Y(_14964_));
 sky130_fd_sc_hd__o21ai_4 _45516_ (.A1(_14714_),
    .A2(_14964_),
    .B1(_14657_),
    .Y(_14965_));
 sky130_fd_sc_hd__nand3_4 _45517_ (.A(_14965_),
    .B(_14960_),
    .C(_14957_),
    .Y(_14966_));
 sky130_fd_sc_hd__nand2_4 _45518_ (.A(_14963_),
    .B(_14966_),
    .Y(_14967_));
 sky130_fd_sc_hd__buf_1 _45519_ (.A(_14732_),
    .X(_14968_));
 sky130_fd_sc_hd__maj3_4 _45520_ (.A(_14736_),
    .B(_14968_),
    .C(_14738_),
    .X(_14969_));
 sky130_vsdinv _45521_ (.A(_14969_),
    .Y(_14970_));
 sky130_vsdinv _45522_ (.A(_14693_),
    .Y(_14971_));
 sky130_fd_sc_hd__a21oi_4 _45523_ (.A1(_14971_),
    .A2(_14462_),
    .B1(_14695_),
    .Y(_14972_));
 sky130_vsdinv _45524_ (.A(_14972_),
    .Y(_14973_));
 sky130_fd_sc_hd__nand3_4 _45525_ (.A(_14973_),
    .B(_14731_),
    .C(_14730_),
    .Y(_14974_));
 sky130_fd_sc_hd__nand2_4 _45526_ (.A(_14968_),
    .B(_14972_),
    .Y(_14975_));
 sky130_fd_sc_hd__a21boi_4 _45527_ (.A1(_14248_),
    .A2(_14729_),
    .B1_N(_14728_),
    .Y(_14976_));
 sky130_vsdinv _45528_ (.A(_14976_),
    .Y(_14977_));
 sky130_fd_sc_hd__a21o_4 _45529_ (.A1(_14974_),
    .A2(_14975_),
    .B1(_14977_),
    .X(_14978_));
 sky130_fd_sc_hd__buf_1 _45530_ (.A(_14977_),
    .X(_14979_));
 sky130_fd_sc_hd__nand3_4 _45531_ (.A(_14974_),
    .B(_14975_),
    .C(_14979_),
    .Y(_14980_));
 sky130_fd_sc_hd__nand3_4 _45532_ (.A(_14970_),
    .B(_14978_),
    .C(_14980_),
    .Y(_14981_));
 sky130_fd_sc_hd__nand2_4 _45533_ (.A(_14978_),
    .B(_14980_),
    .Y(_14982_));
 sky130_fd_sc_hd__nand2_4 _45534_ (.A(_14982_),
    .B(_14969_),
    .Y(_14983_));
 sky130_fd_sc_hd__nand2_4 _45535_ (.A(_14981_),
    .B(_14983_),
    .Y(_14984_));
 sky130_fd_sc_hd__nand2_4 _45536_ (.A(_14984_),
    .B(_13745_),
    .Y(_14985_));
 sky130_fd_sc_hd__nand3_4 _45537_ (.A(_14981_),
    .B(_14983_),
    .C(_13747_),
    .Y(_14986_));
 sky130_fd_sc_hd__nand2_4 _45538_ (.A(_14985_),
    .B(_14986_),
    .Y(_14987_));
 sky130_fd_sc_hd__a21boi_4 _45539_ (.A1(_14705_),
    .A2(_14712_),
    .B1_N(_14708_),
    .Y(_14988_));
 sky130_fd_sc_hd__nand2_4 _45540_ (.A(_14987_),
    .B(_14988_),
    .Y(_14989_));
 sky130_fd_sc_hd__a21oi_4 _45541_ (.A1(_14701_),
    .A2(_14702_),
    .B1(_14706_),
    .Y(_14990_));
 sky130_fd_sc_hd__o21ai_4 _45542_ (.A1(_14710_),
    .A2(_14990_),
    .B1(_14708_),
    .Y(_14991_));
 sky130_fd_sc_hd__nand3_4 _45543_ (.A(_14991_),
    .B(_14986_),
    .C(_14985_),
    .Y(_14992_));
 sky130_fd_sc_hd__nand2_4 _45544_ (.A(_14989_),
    .B(_14992_),
    .Y(_14993_));
 sky130_fd_sc_hd__a21boi_4 _45545_ (.A1(_14744_),
    .A2(_14273_),
    .B1_N(_14746_),
    .Y(_14994_));
 sky130_fd_sc_hd__nand2_4 _45546_ (.A(_14993_),
    .B(_14994_),
    .Y(_14995_));
 sky130_vsdinv _45547_ (.A(_14994_),
    .Y(_14996_));
 sky130_fd_sc_hd__nand3_4 _45548_ (.A(_14989_),
    .B(_14992_),
    .C(_14996_),
    .Y(_14997_));
 sky130_fd_sc_hd__nand2_4 _45549_ (.A(_14995_),
    .B(_14997_),
    .Y(_14998_));
 sky130_fd_sc_hd__nand2_4 _45550_ (.A(_14967_),
    .B(_14998_),
    .Y(_14999_));
 sky130_vsdinv _45551_ (.A(_14998_),
    .Y(_15000_));
 sky130_fd_sc_hd__nand3_4 _45552_ (.A(_15000_),
    .B(_14966_),
    .C(_14963_),
    .Y(_15001_));
 sky130_fd_sc_hd__nand2_4 _45553_ (.A(_14999_),
    .B(_15001_),
    .Y(_15002_));
 sky130_fd_sc_hd__a21boi_4 _45554_ (.A1(_14766_),
    .A2(_14722_),
    .B1_N(_14724_),
    .Y(_15003_));
 sky130_fd_sc_hd__nand2_4 _45555_ (.A(_15002_),
    .B(_15003_),
    .Y(_15004_));
 sky130_fd_sc_hd__a21boi_4 _45556_ (.A1(_14715_),
    .A2(_14719_),
    .B1_N(_14721_),
    .Y(_15005_));
 sky130_fd_sc_hd__o21ai_4 _45557_ (.A1(_14762_),
    .A2(_15005_),
    .B1(_14724_),
    .Y(_15006_));
 sky130_fd_sc_hd__nand3_4 _45558_ (.A(_15006_),
    .B(_14999_),
    .C(_15001_),
    .Y(_15007_));
 sky130_fd_sc_hd__nand2_4 _45559_ (.A(_15004_),
    .B(_15007_),
    .Y(_15008_));
 sky130_fd_sc_hd__a21boi_4 _45560_ (.A1(_14752_),
    .A2(_14760_),
    .B1_N(_14755_),
    .Y(_15009_));
 sky130_fd_sc_hd__xor2_4 _45561_ (.A(_13776_),
    .B(_15009_),
    .X(_15010_));
 sky130_fd_sc_hd__nand2_4 _45562_ (.A(_15008_),
    .B(_15010_),
    .Y(_15011_));
 sky130_vsdinv _45563_ (.A(_15010_),
    .Y(_15012_));
 sky130_fd_sc_hd__nand3_4 _45564_ (.A(_15004_),
    .B(_15007_),
    .C(_15012_),
    .Y(_15013_));
 sky130_fd_sc_hd__nand2_4 _45565_ (.A(_15011_),
    .B(_15013_),
    .Y(_15014_));
 sky130_fd_sc_hd__a21boi_4 _45566_ (.A1(_14770_),
    .A2(_14777_),
    .B1_N(_14772_),
    .Y(_15015_));
 sky130_fd_sc_hd__nand2_4 _45567_ (.A(_15014_),
    .B(_15015_),
    .Y(_15016_));
 sky130_fd_sc_hd__nand2_4 _45568_ (.A(_14778_),
    .B(_14772_),
    .Y(_15017_));
 sky130_fd_sc_hd__nand3_4 _45569_ (.A(_15017_),
    .B(_15011_),
    .C(_15013_),
    .Y(_15018_));
 sky130_fd_sc_hd__nand2_4 _45570_ (.A(_15016_),
    .B(_15018_),
    .Y(_15019_));
 sky130_fd_sc_hd__a21oi_4 _45571_ (.A1(_14527_),
    .A2(_14522_),
    .B1(_14303_),
    .Y(_15020_));
 sky130_vsdinv _45572_ (.A(_15020_),
    .Y(_15021_));
 sky130_fd_sc_hd__nand2_4 _45573_ (.A(_15019_),
    .B(_15021_),
    .Y(_15022_));
 sky130_fd_sc_hd__nand3_4 _45574_ (.A(_15016_),
    .B(_15018_),
    .C(_15020_),
    .Y(_15023_));
 sky130_fd_sc_hd__nand2_4 _45575_ (.A(_15022_),
    .B(_15023_),
    .Y(_15024_));
 sky130_fd_sc_hd__a21boi_4 _45576_ (.A1(_14781_),
    .A2(_14785_),
    .B1_N(_14783_),
    .Y(_15025_));
 sky130_fd_sc_hd__nand2_4 _45577_ (.A(_15024_),
    .B(_15025_),
    .Y(_15026_));
 sky130_fd_sc_hd__nand2_4 _45578_ (.A(_14788_),
    .B(_14783_),
    .Y(_15027_));
 sky130_fd_sc_hd__nand3_4 _45579_ (.A(_15027_),
    .B(_15022_),
    .C(_15023_),
    .Y(_15028_));
 sky130_fd_sc_hd__nand2_4 _45580_ (.A(_15026_),
    .B(_15028_),
    .Y(_15029_));
 sky130_fd_sc_hd__a21boi_4 _45581_ (.A1(_14802_),
    .A2(_14791_),
    .B1_N(_14793_),
    .Y(_15030_));
 sky130_fd_sc_hd__xor2_4 _45582_ (.A(_15029_),
    .B(_15030_),
    .X(_01450_));
 sky130_fd_sc_hd__nand2_4 _45583_ (.A(_03315_),
    .B(_14565_),
    .Y(_15031_));
 sky130_fd_sc_hd__o21ai_4 _45584_ (.A1(_03319_),
    .A2(_03629_),
    .B1(_15031_),
    .Y(_15032_));
 sky130_fd_sc_hd__buf_1 _45585_ (.A(_03628_),
    .X(_15033_));
 sky130_fd_sc_hd__nand4_4 _45586_ (.A(_03315_),
    .B(_07858_),
    .C(_15033_),
    .D(_11384_),
    .Y(_15034_));
 sky130_fd_sc_hd__nand2_4 _45587_ (.A(_07621_),
    .B(_03620_),
    .Y(_15035_));
 sky130_vsdinv _45588_ (.A(_15035_),
    .Y(_15036_));
 sky130_fd_sc_hd__a21o_4 _45589_ (.A1(_15032_),
    .A2(_15034_),
    .B1(_15036_),
    .X(_15037_));
 sky130_fd_sc_hd__nand3_4 _45590_ (.A(_15032_),
    .B(_15034_),
    .C(_15036_),
    .Y(_15038_));
 sky130_fd_sc_hd__nand2_4 _45591_ (.A(_15037_),
    .B(_15038_),
    .Y(_15039_));
 sky130_fd_sc_hd__a21boi_4 _45592_ (.A1(_14809_),
    .A2(_14811_),
    .B1_N(_14812_),
    .Y(_15040_));
 sky130_fd_sc_hd__nand2_4 _45593_ (.A(_15039_),
    .B(_15040_),
    .Y(_15041_));
 sky130_vsdinv _45594_ (.A(_15040_),
    .Y(_15042_));
 sky130_fd_sc_hd__nand3_4 _45595_ (.A(_15042_),
    .B(_15037_),
    .C(_15038_),
    .Y(_15043_));
 sky130_fd_sc_hd__nand2_4 _45596_ (.A(_15041_),
    .B(_15043_),
    .Y(_15044_));
 sky130_fd_sc_hd__nand2_4 _45597_ (.A(_14096_),
    .B(_12404_),
    .Y(_15045_));
 sky130_fd_sc_hd__nand2_4 _45598_ (.A(_07630_),
    .B(_12406_),
    .Y(_15046_));
 sky130_fd_sc_hd__nand2_4 _45599_ (.A(_15045_),
    .B(_15046_),
    .Y(_15047_));
 sky130_fd_sc_hd__nand4_4 _45600_ (.A(_07627_),
    .B(_11015_),
    .C(_12409_),
    .D(_12410_),
    .Y(_15048_));
 sky130_fd_sc_hd__nand2_4 _45601_ (.A(_13340_),
    .B(_10512_),
    .Y(_15049_));
 sky130_vsdinv _45602_ (.A(_15049_),
    .Y(_15050_));
 sky130_fd_sc_hd__a21oi_4 _45603_ (.A1(_15047_),
    .A2(_15048_),
    .B1(_15050_),
    .Y(_15051_));
 sky130_fd_sc_hd__nand3_4 _45604_ (.A(_15047_),
    .B(_15048_),
    .C(_15050_),
    .Y(_15052_));
 sky130_vsdinv _45605_ (.A(_15052_),
    .Y(_15053_));
 sky130_fd_sc_hd__nor2_4 _45606_ (.A(_15051_),
    .B(_15053_),
    .Y(_15054_));
 sky130_vsdinv _45607_ (.A(_15054_),
    .Y(_15055_));
 sky130_fd_sc_hd__nand2_4 _45608_ (.A(_15044_),
    .B(_15055_),
    .Y(_15056_));
 sky130_fd_sc_hd__nand3_4 _45609_ (.A(_15041_),
    .B(_15054_),
    .C(_15043_),
    .Y(_15057_));
 sky130_fd_sc_hd__nand2_4 _45610_ (.A(_15056_),
    .B(_15057_),
    .Y(_15058_));
 sky130_fd_sc_hd__a21boi_4 _45611_ (.A1(_14829_),
    .A2(_14818_),
    .B1_N(_14816_),
    .Y(_15059_));
 sky130_fd_sc_hd__nand2_4 _45612_ (.A(_15058_),
    .B(_15059_),
    .Y(_15060_));
 sky130_vsdinv _45613_ (.A(_15059_),
    .Y(_15061_));
 sky130_fd_sc_hd__nand3_4 _45614_ (.A(_15061_),
    .B(_15057_),
    .C(_15056_),
    .Y(_15062_));
 sky130_fd_sc_hd__nand2_4 _45615_ (.A(_15060_),
    .B(_15062_),
    .Y(_15063_));
 sky130_fd_sc_hd__nand2_4 _45616_ (.A(_11242_),
    .B(_13298_),
    .Y(_15064_));
 sky130_fd_sc_hd__nand2_4 _45617_ (.A(_13342_),
    .B(_12111_),
    .Y(_15065_));
 sky130_fd_sc_hd__nand2_4 _45618_ (.A(_15064_),
    .B(_15065_),
    .Y(_15066_));
 sky130_fd_sc_hd__nand4_4 _45619_ (.A(_08309_),
    .B(_08315_),
    .C(_12430_),
    .D(_12115_),
    .Y(_15067_));
 sky130_fd_sc_hd__nand2_4 _45620_ (.A(_08755_),
    .B(_13303_),
    .Y(_15068_));
 sky130_vsdinv _45621_ (.A(_15068_),
    .Y(_15069_));
 sky130_fd_sc_hd__a21o_4 _45622_ (.A1(_15066_),
    .A2(_15067_),
    .B1(_15069_),
    .X(_15070_));
 sky130_fd_sc_hd__nand3_4 _45623_ (.A(_15066_),
    .B(_15067_),
    .C(_15069_),
    .Y(_15071_));
 sky130_fd_sc_hd__a21boi_4 _45624_ (.A1(_14822_),
    .A2(_14825_),
    .B1_N(_14823_),
    .Y(_15072_));
 sky130_fd_sc_hd__a21boi_4 _45625_ (.A1(_15070_),
    .A2(_15071_),
    .B1_N(_15072_),
    .Y(_15073_));
 sky130_vsdinv _45626_ (.A(_15073_),
    .Y(_15074_));
 sky130_vsdinv _45627_ (.A(_15072_),
    .Y(_15075_));
 sky130_fd_sc_hd__nand3_4 _45628_ (.A(_15075_),
    .B(_15070_),
    .C(_15071_),
    .Y(_15076_));
 sky130_fd_sc_hd__a21boi_4 _45629_ (.A1(_14843_),
    .A2(_14846_),
    .B1_N(_14844_),
    .Y(_15077_));
 sky130_vsdinv _45630_ (.A(_15077_),
    .Y(_15078_));
 sky130_fd_sc_hd__a21oi_4 _45631_ (.A1(_15074_),
    .A2(_15076_),
    .B1(_15078_),
    .Y(_15079_));
 sky130_fd_sc_hd__nand3_4 _45632_ (.A(_15074_),
    .B(_15078_),
    .C(_15076_),
    .Y(_15080_));
 sky130_vsdinv _45633_ (.A(_15080_),
    .Y(_15081_));
 sky130_fd_sc_hd__nor2_4 _45634_ (.A(_15079_),
    .B(_15081_),
    .Y(_15082_));
 sky130_vsdinv _45635_ (.A(_15082_),
    .Y(_15083_));
 sky130_fd_sc_hd__nand2_4 _45636_ (.A(_15063_),
    .B(_15083_),
    .Y(_15084_));
 sky130_fd_sc_hd__nand3_4 _45637_ (.A(_15060_),
    .B(_15062_),
    .C(_15082_),
    .Y(_15085_));
 sky130_fd_sc_hd__nand2_4 _45638_ (.A(_15084_),
    .B(_15085_),
    .Y(_15086_));
 sky130_fd_sc_hd__o21a_4 _45639_ (.A1(_14857_),
    .A2(_14838_),
    .B1(_14837_),
    .X(_15087_));
 sky130_fd_sc_hd__nand2_4 _45640_ (.A(_15086_),
    .B(_15087_),
    .Y(_15088_));
 sky130_fd_sc_hd__nand2_4 _45641_ (.A(_14859_),
    .B(_14837_),
    .Y(_15089_));
 sky130_fd_sc_hd__nand3_4 _45642_ (.A(_15089_),
    .B(_15085_),
    .C(_15084_),
    .Y(_15090_));
 sky130_fd_sc_hd__nand2_4 _45643_ (.A(_15088_),
    .B(_15090_),
    .Y(_15091_));
 sky130_fd_sc_hd__nand2_4 _45644_ (.A(_13376_),
    .B(_12157_),
    .Y(_15092_));
 sky130_fd_sc_hd__nand2_4 _45645_ (.A(_12817_),
    .B(_12156_),
    .Y(_15093_));
 sky130_fd_sc_hd__nand2_4 _45646_ (.A(_15092_),
    .B(_15093_),
    .Y(_15094_));
 sky130_fd_sc_hd__nand4_4 _45647_ (.A(_11595_),
    .B(_10785_),
    .C(_03570_),
    .D(_12467_),
    .Y(_15095_));
 sky130_fd_sc_hd__nand2_4 _45648_ (.A(_09578_),
    .B(_10540_),
    .Y(_15096_));
 sky130_vsdinv _45649_ (.A(_15096_),
    .Y(_15097_));
 sky130_fd_sc_hd__a21o_4 _45650_ (.A1(_15094_),
    .A2(_15095_),
    .B1(_15097_),
    .X(_15098_));
 sky130_fd_sc_hd__nand3_4 _45651_ (.A(_15094_),
    .B(_15095_),
    .C(_15097_),
    .Y(_15099_));
 sky130_fd_sc_hd__nand2_4 _45652_ (.A(_15098_),
    .B(_15099_),
    .Y(_15100_));
 sky130_fd_sc_hd__a21o_4 _45653_ (.A1(_14874_),
    .A2(_14878_),
    .B1(_15100_),
    .X(_15101_));
 sky130_fd_sc_hd__nand3_4 _45654_ (.A(_15100_),
    .B(_14874_),
    .C(_14878_),
    .Y(_15102_));
 sky130_fd_sc_hd__nand2_4 _45655_ (.A(_14426_),
    .B(_12456_),
    .Y(_15103_));
 sky130_fd_sc_hd__nand2_4 _45656_ (.A(_11949_),
    .B(_11187_),
    .Y(_15104_));
 sky130_fd_sc_hd__nand2_4 _45657_ (.A(_13127_),
    .B(_11518_),
    .Y(_15105_));
 sky130_fd_sc_hd__xnor2_4 _45658_ (.A(_15104_),
    .B(_15105_),
    .Y(_15106_));
 sky130_fd_sc_hd__xor2_4 _45659_ (.A(_15103_),
    .B(_15106_),
    .X(_15107_));
 sky130_fd_sc_hd__a21o_4 _45660_ (.A1(_15101_),
    .A2(_15102_),
    .B1(_15107_),
    .X(_15108_));
 sky130_fd_sc_hd__nand3_4 _45661_ (.A(_15107_),
    .B(_15101_),
    .C(_15102_),
    .Y(_15109_));
 sky130_fd_sc_hd__maj3_4 _45662_ (.A(_14852_),
    .B(_14849_),
    .C(_14840_),
    .X(_15110_));
 sky130_vsdinv _45663_ (.A(_15110_),
    .Y(_15111_));
 sky130_fd_sc_hd__a21o_4 _45664_ (.A1(_15108_),
    .A2(_15109_),
    .B1(_15111_),
    .X(_15112_));
 sky130_fd_sc_hd__nand3_4 _45665_ (.A(_15108_),
    .B(_15111_),
    .C(_15109_),
    .Y(_15113_));
 sky130_fd_sc_hd__a21boi_4 _45666_ (.A1(_14889_),
    .A2(_14881_),
    .B1_N(_14880_),
    .Y(_15114_));
 sky130_vsdinv _45667_ (.A(_15114_),
    .Y(_15115_));
 sky130_fd_sc_hd__a21oi_4 _45668_ (.A1(_15112_),
    .A2(_15113_),
    .B1(_15115_),
    .Y(_15116_));
 sky130_vsdinv _45669_ (.A(_15116_),
    .Y(_15117_));
 sky130_fd_sc_hd__nand3_4 _45670_ (.A(_15112_),
    .B(_15115_),
    .C(_15113_),
    .Y(_15118_));
 sky130_fd_sc_hd__nand2_4 _45671_ (.A(_15117_),
    .B(_15118_),
    .Y(_15119_));
 sky130_fd_sc_hd__nand2_4 _45672_ (.A(_15091_),
    .B(_15119_),
    .Y(_15120_));
 sky130_vsdinv _45673_ (.A(_15118_),
    .Y(_15121_));
 sky130_fd_sc_hd__nor2_4 _45674_ (.A(_15116_),
    .B(_15121_),
    .Y(_15122_));
 sky130_fd_sc_hd__nand3_4 _45675_ (.A(_15122_),
    .B(_15090_),
    .C(_15088_),
    .Y(_15123_));
 sky130_fd_sc_hd__nand2_4 _45676_ (.A(_15120_),
    .B(_15123_),
    .Y(_15124_));
 sky130_fd_sc_hd__o21a_4 _45677_ (.A1(_14900_),
    .A2(_14866_),
    .B1(_14865_),
    .X(_15125_));
 sky130_fd_sc_hd__nand2_4 _45678_ (.A(_15124_),
    .B(_15125_),
    .Y(_15126_));
 sky130_fd_sc_hd__nand2_4 _45679_ (.A(_14902_),
    .B(_14865_),
    .Y(_15127_));
 sky130_fd_sc_hd__nand3_4 _45680_ (.A(_15127_),
    .B(_15123_),
    .C(_15120_),
    .Y(_15128_));
 sky130_fd_sc_hd__nand2_4 _45681_ (.A(_15126_),
    .B(_15128_),
    .Y(_15129_));
 sky130_vsdinv _45682_ (.A(_14883_),
    .Y(_15130_));
 sky130_fd_sc_hd__nand3_4 _45683_ (.A(_14886_),
    .B(_14887_),
    .C(_15130_),
    .Y(_15131_));
 sky130_fd_sc_hd__buf_1 _45684_ (.A(_12878_),
    .X(_15132_));
 sky130_fd_sc_hd__nand2_4 _45685_ (.A(_15132_),
    .B(_11873_),
    .Y(_15133_));
 sky130_fd_sc_hd__nand2_4 _45686_ (.A(_03397_),
    .B(_11872_),
    .Y(_15134_));
 sky130_fd_sc_hd__nand2_4 _45687_ (.A(_15133_),
    .B(_15134_),
    .Y(_15135_));
 sky130_fd_sc_hd__buf_1 _45688_ (.A(_11323_),
    .X(_15136_));
 sky130_fd_sc_hd__nand4_4 _45689_ (.A(_15136_),
    .B(_13410_),
    .C(_03537_),
    .D(_03542_),
    .Y(_15137_));
 sky130_fd_sc_hd__nand2_4 _45690_ (.A(_10837_),
    .B(_07337_),
    .Y(_15138_));
 sky130_vsdinv _45691_ (.A(_15138_),
    .Y(_15139_));
 sky130_fd_sc_hd__a21o_4 _45692_ (.A1(_15135_),
    .A2(_15137_),
    .B1(_15139_),
    .X(_15140_));
 sky130_fd_sc_hd__nand3_4 _45693_ (.A(_15135_),
    .B(_15137_),
    .C(_15139_),
    .Y(_15141_));
 sky130_fd_sc_hd__nand2_4 _45694_ (.A(_15140_),
    .B(_15141_),
    .Y(_15142_));
 sky130_fd_sc_hd__a21o_4 _45695_ (.A1(_14887_),
    .A2(_15131_),
    .B1(_15142_),
    .X(_15143_));
 sky130_fd_sc_hd__a21boi_4 _45696_ (.A1(_14886_),
    .A2(_15130_),
    .B1_N(_14887_),
    .Y(_15144_));
 sky130_fd_sc_hd__nand2_4 _45697_ (.A(_15142_),
    .B(_15144_),
    .Y(_15145_));
 sky130_fd_sc_hd__a21boi_4 _45698_ (.A1(_14910_),
    .A2(_14913_),
    .B1_N(_14911_),
    .Y(_15146_));
 sky130_vsdinv _45699_ (.A(_15146_),
    .Y(_15147_));
 sky130_fd_sc_hd__a21o_4 _45700_ (.A1(_15143_),
    .A2(_15145_),
    .B1(_15147_),
    .X(_15148_));
 sky130_fd_sc_hd__nand3_4 _45701_ (.A(_15143_),
    .B(_15147_),
    .C(_15145_),
    .Y(_15149_));
 sky130_fd_sc_hd__maj3_4 _45702_ (.A(_14919_),
    .B(_14916_),
    .C(_14907_),
    .X(_15150_));
 sky130_vsdinv _45703_ (.A(_15150_),
    .Y(_15151_));
 sky130_fd_sc_hd__a21o_4 _45704_ (.A1(_15148_),
    .A2(_15149_),
    .B1(_15151_),
    .X(_15152_));
 sky130_fd_sc_hd__nand3_4 _45705_ (.A(_15151_),
    .B(_15148_),
    .C(_15149_),
    .Y(_15153_));
 sky130_fd_sc_hd__o21a_4 _45706_ (.A1(_12527_),
    .A2(_07523_),
    .B1(_11692_),
    .X(_15154_));
 sky130_fd_sc_hd__nand3_4 _45707_ (.A(_12910_),
    .B(_03519_),
    .C(_11905_),
    .Y(_15155_));
 sky130_fd_sc_hd__a21o_4 _45708_ (.A1(_15154_),
    .A2(_15155_),
    .B1(_14687_),
    .X(_15156_));
 sky130_fd_sc_hd__nand3_4 _45709_ (.A(_15154_),
    .B(_14687_),
    .C(_15155_),
    .Y(_15157_));
 sky130_fd_sc_hd__a21boi_4 _45710_ (.A1(_14931_),
    .A2(_14690_),
    .B1_N(_14932_),
    .Y(_15158_));
 sky130_vsdinv _45711_ (.A(_15158_),
    .Y(_15159_));
 sky130_fd_sc_hd__a21o_4 _45712_ (.A1(_15156_),
    .A2(_15157_),
    .B1(_15159_),
    .X(_15160_));
 sky130_fd_sc_hd__nand3_4 _45713_ (.A(_15159_),
    .B(_15156_),
    .C(_15157_),
    .Y(_15161_));
 sky130_fd_sc_hd__nand2_4 _45714_ (.A(_15160_),
    .B(_15161_),
    .Y(_15162_));
 sky130_fd_sc_hd__xor2_4 _45715_ (.A(_14464_),
    .B(_15162_),
    .X(_15163_));
 sky130_fd_sc_hd__a21o_4 _45716_ (.A1(_15152_),
    .A2(_15153_),
    .B1(_15163_),
    .X(_15164_));
 sky130_fd_sc_hd__nand3_4 _45717_ (.A(_15152_),
    .B(_15163_),
    .C(_15153_),
    .Y(_15165_));
 sky130_fd_sc_hd__nand2_4 _45718_ (.A(_14899_),
    .B(_14895_),
    .Y(_15166_));
 sky130_fd_sc_hd__a21oi_4 _45719_ (.A1(_15164_),
    .A2(_15165_),
    .B1(_15166_),
    .Y(_15167_));
 sky130_fd_sc_hd__nand3_4 _45720_ (.A(_15166_),
    .B(_15164_),
    .C(_15165_),
    .Y(_15168_));
 sky130_vsdinv _45721_ (.A(_15168_),
    .Y(_15169_));
 sky130_fd_sc_hd__a21boi_4 _45722_ (.A1(_14925_),
    .A2(_14942_),
    .B1_N(_14927_),
    .Y(_15170_));
 sky130_fd_sc_hd__o21ai_4 _45723_ (.A1(_15167_),
    .A2(_15169_),
    .B1(_15170_),
    .Y(_15171_));
 sky130_vsdinv _45724_ (.A(_15167_),
    .Y(_15172_));
 sky130_vsdinv _45725_ (.A(_15170_),
    .Y(_15173_));
 sky130_fd_sc_hd__nand3_4 _45726_ (.A(_15172_),
    .B(_15173_),
    .C(_15168_),
    .Y(_15174_));
 sky130_fd_sc_hd__nand2_4 _45727_ (.A(_15171_),
    .B(_15174_),
    .Y(_15175_));
 sky130_fd_sc_hd__nand2_4 _45728_ (.A(_15129_),
    .B(_15175_),
    .Y(_15176_));
 sky130_fd_sc_hd__nand4_4 _45729_ (.A(_15174_),
    .B(_15126_),
    .C(_15171_),
    .D(_15128_),
    .Y(_15177_));
 sky130_fd_sc_hd__nand2_4 _45730_ (.A(_15176_),
    .B(_15177_),
    .Y(_15178_));
 sky130_vsdinv _45731_ (.A(_14905_),
    .Y(_15179_));
 sky130_fd_sc_hd__a21oi_4 _45732_ (.A1(_14959_),
    .A2(_14904_),
    .B1(_15179_),
    .Y(_15180_));
 sky130_fd_sc_hd__nand2_4 _45733_ (.A(_15178_),
    .B(_15180_),
    .Y(_15181_));
 sky130_fd_sc_hd__a21o_4 _45734_ (.A1(_14959_),
    .A2(_14904_),
    .B1(_15179_),
    .X(_15182_));
 sky130_fd_sc_hd__nand3_4 _45735_ (.A(_15182_),
    .B(_15177_),
    .C(_15176_),
    .Y(_15183_));
 sky130_fd_sc_hd__nand2_4 _45736_ (.A(_15181_),
    .B(_15183_),
    .Y(_15184_));
 sky130_fd_sc_hd__a21o_4 _45737_ (.A1(_14940_),
    .A2(_14937_),
    .B1(_14968_),
    .X(_15185_));
 sky130_fd_sc_hd__a21oi_4 _45738_ (.A1(_14938_),
    .A2(_14464_),
    .B1(_14936_),
    .Y(_15186_));
 sky130_fd_sc_hd__nand2_4 _45739_ (.A(_14735_),
    .B(_15186_),
    .Y(_15187_));
 sky130_fd_sc_hd__a21o_4 _45740_ (.A1(_15185_),
    .A2(_15187_),
    .B1(_14979_),
    .X(_15188_));
 sky130_fd_sc_hd__nand3_4 _45741_ (.A(_15185_),
    .B(_14979_),
    .C(_15187_),
    .Y(_15189_));
 sky130_fd_sc_hd__nand2_4 _45742_ (.A(_15188_),
    .B(_15189_),
    .Y(_15190_));
 sky130_fd_sc_hd__a21boi_4 _45743_ (.A1(_14975_),
    .A2(_14979_),
    .B1_N(_14974_),
    .Y(_15191_));
 sky130_fd_sc_hd__nand2_4 _45744_ (.A(_15190_),
    .B(_15191_),
    .Y(_15192_));
 sky130_vsdinv _45745_ (.A(_15191_),
    .Y(_15193_));
 sky130_fd_sc_hd__nand3_4 _45746_ (.A(_15188_),
    .B(_15193_),
    .C(_15189_),
    .Y(_15194_));
 sky130_fd_sc_hd__nand2_4 _45747_ (.A(_15192_),
    .B(_15194_),
    .Y(_15195_));
 sky130_fd_sc_hd__nand2_4 _45748_ (.A(_15195_),
    .B(_13480_),
    .Y(_15196_));
 sky130_fd_sc_hd__nand3_4 _45749_ (.A(_15192_),
    .B(_13747_),
    .C(_15194_),
    .Y(_15197_));
 sky130_fd_sc_hd__nand2_4 _45750_ (.A(_15196_),
    .B(_15197_),
    .Y(_15198_));
 sky130_fd_sc_hd__a21boi_4 _45751_ (.A1(_14949_),
    .A2(_14952_),
    .B1_N(_14950_),
    .Y(_15199_));
 sky130_fd_sc_hd__nand2_4 _45752_ (.A(_15198_),
    .B(_15199_),
    .Y(_15200_));
 sky130_vsdinv _45753_ (.A(_15199_),
    .Y(_15201_));
 sky130_fd_sc_hd__nand3_4 _45754_ (.A(_15201_),
    .B(_15197_),
    .C(_15196_),
    .Y(_15202_));
 sky130_fd_sc_hd__buf_1 _45755_ (.A(_15202_),
    .X(_15203_));
 sky130_fd_sc_hd__a21boi_4 _45756_ (.A1(_14757_),
    .A2(_14983_),
    .B1_N(_14981_),
    .Y(_15204_));
 sky130_vsdinv _45757_ (.A(_15204_),
    .Y(_15205_));
 sky130_fd_sc_hd__a21o_4 _45758_ (.A1(_15200_),
    .A2(_15203_),
    .B1(_15205_),
    .X(_15206_));
 sky130_fd_sc_hd__nand3_4 _45759_ (.A(_15200_),
    .B(_15202_),
    .C(_15205_),
    .Y(_15207_));
 sky130_fd_sc_hd__nand2_4 _45760_ (.A(_15206_),
    .B(_15207_),
    .Y(_15208_));
 sky130_fd_sc_hd__nand2_4 _45761_ (.A(_15184_),
    .B(_15208_),
    .Y(_15209_));
 sky130_fd_sc_hd__a21oi_4 _45762_ (.A1(_15200_),
    .A2(_15203_),
    .B1(_15205_),
    .Y(_15210_));
 sky130_vsdinv _45763_ (.A(_15207_),
    .Y(_15211_));
 sky130_fd_sc_hd__nor2_4 _45764_ (.A(_15210_),
    .B(_15211_),
    .Y(_15212_));
 sky130_fd_sc_hd__nand3_4 _45765_ (.A(_15212_),
    .B(_15181_),
    .C(_15183_),
    .Y(_15213_));
 sky130_fd_sc_hd__nand2_4 _45766_ (.A(_15209_),
    .B(_15213_),
    .Y(_15214_));
 sky130_vsdinv _45767_ (.A(_14966_),
    .Y(_15215_));
 sky130_fd_sc_hd__a21oi_4 _45768_ (.A1(_15000_),
    .A2(_14963_),
    .B1(_15215_),
    .Y(_15216_));
 sky130_fd_sc_hd__nand2_4 _45769_ (.A(_15214_),
    .B(_15216_),
    .Y(_15217_));
 sky130_fd_sc_hd__a21o_4 _45770_ (.A1(_15000_),
    .A2(_14963_),
    .B1(_15215_),
    .X(_15218_));
 sky130_fd_sc_hd__nand3_4 _45771_ (.A(_15218_),
    .B(_15213_),
    .C(_15209_),
    .Y(_15219_));
 sky130_fd_sc_hd__nand2_4 _45772_ (.A(_15217_),
    .B(_15219_),
    .Y(_15220_));
 sky130_fd_sc_hd__a21boi_4 _45773_ (.A1(_14989_),
    .A2(_14996_),
    .B1_N(_14992_),
    .Y(_15221_));
 sky130_fd_sc_hd__xor2_4 _45774_ (.A(_14291_),
    .B(_15221_),
    .X(_15222_));
 sky130_fd_sc_hd__nand2_4 _45775_ (.A(_15220_),
    .B(_15222_),
    .Y(_15223_));
 sky130_vsdinv _45776_ (.A(_15222_),
    .Y(_15224_));
 sky130_fd_sc_hd__nand3_4 _45777_ (.A(_15217_),
    .B(_15219_),
    .C(_15224_),
    .Y(_15225_));
 sky130_fd_sc_hd__nand2_4 _45778_ (.A(_15223_),
    .B(_15225_),
    .Y(_15226_));
 sky130_fd_sc_hd__a21boi_4 _45779_ (.A1(_15004_),
    .A2(_15012_),
    .B1_N(_15007_),
    .Y(_15227_));
 sky130_fd_sc_hd__nand2_4 _45780_ (.A(_15226_),
    .B(_15227_),
    .Y(_15228_));
 sky130_vsdinv _45781_ (.A(_15227_),
    .Y(_15229_));
 sky130_fd_sc_hd__nand3_4 _45782_ (.A(_15229_),
    .B(_15223_),
    .C(_15225_),
    .Y(_15230_));
 sky130_fd_sc_hd__nand2_4 _45783_ (.A(_15228_),
    .B(_15230_),
    .Y(_15231_));
 sky130_fd_sc_hd__a21oi_4 _45784_ (.A1(_14761_),
    .A2(_14755_),
    .B1(_14050_),
    .Y(_15232_));
 sky130_vsdinv _45785_ (.A(_15232_),
    .Y(_15233_));
 sky130_fd_sc_hd__nand2_4 _45786_ (.A(_15231_),
    .B(_15233_),
    .Y(_15234_));
 sky130_fd_sc_hd__nand3_4 _45787_ (.A(_15228_),
    .B(_15230_),
    .C(_15232_),
    .Y(_15235_));
 sky130_fd_sc_hd__nand2_4 _45788_ (.A(_15234_),
    .B(_15235_),
    .Y(_15236_));
 sky130_fd_sc_hd__a21boi_4 _45789_ (.A1(_15016_),
    .A2(_15020_),
    .B1_N(_15018_),
    .Y(_15237_));
 sky130_fd_sc_hd__nand2_4 _45790_ (.A(_15236_),
    .B(_15237_),
    .Y(_15238_));
 sky130_vsdinv _45791_ (.A(_15237_),
    .Y(_15239_));
 sky130_fd_sc_hd__nand3_4 _45792_ (.A(_15239_),
    .B(_15234_),
    .C(_15235_),
    .Y(_15240_));
 sky130_fd_sc_hd__nand2_4 _45793_ (.A(_15238_),
    .B(_15240_),
    .Y(_15241_));
 sky130_fd_sc_hd__nor2_4 _45794_ (.A(_15029_),
    .B(_14794_),
    .Y(_15242_));
 sky130_fd_sc_hd__o21ai_4 _45795_ (.A1(_14797_),
    .A2(_14800_),
    .B1(_15242_),
    .Y(_15243_));
 sky130_fd_sc_hd__nand2_4 _45796_ (.A(_14793_),
    .B(_15028_),
    .Y(_15244_));
 sky130_fd_sc_hd__nand2_4 _45797_ (.A(_15244_),
    .B(_15026_),
    .Y(_15245_));
 sky130_fd_sc_hd__nand2_4 _45798_ (.A(_15243_),
    .B(_15245_),
    .Y(_15246_));
 sky130_fd_sc_hd__xnor2_4 _45799_ (.A(_15241_),
    .B(_15246_),
    .Y(_01451_));
 sky130_fd_sc_hd__a21boi_4 _45800_ (.A1(_15032_),
    .A2(_15036_),
    .B1_N(_15034_),
    .Y(_15247_));
 sky130_vsdinv _45801_ (.A(_15247_),
    .Y(_15248_));
 sky130_fd_sc_hd__buf_1 _45802_ (.A(_13808_),
    .X(_15249_));
 sky130_fd_sc_hd__buf_1 _45803_ (.A(_11438_),
    .X(_15250_));
 sky130_fd_sc_hd__nand2_4 _45804_ (.A(_07295_),
    .B(_15250_),
    .Y(_15251_));
 sky130_fd_sc_hd__o21ai_4 _45805_ (.A1(_11513_),
    .A2(_15249_),
    .B1(_15251_),
    .Y(_15252_));
 sky130_fd_sc_hd__buf_1 _45806_ (.A(_14565_),
    .X(_15253_));
 sky130_fd_sc_hd__nand4_4 _45807_ (.A(_03319_),
    .B(_07295_),
    .C(_15250_),
    .D(_15253_),
    .Y(_15254_));
 sky130_fd_sc_hd__nand2_4 _45808_ (.A(_13042_),
    .B(_10517_),
    .Y(_15255_));
 sky130_vsdinv _45809_ (.A(_15255_),
    .Y(_15256_));
 sky130_fd_sc_hd__a21o_4 _45810_ (.A1(_15252_),
    .A2(_15254_),
    .B1(_15256_),
    .X(_15257_));
 sky130_fd_sc_hd__nand3_4 _45811_ (.A(_15252_),
    .B(_15254_),
    .C(_15256_),
    .Y(_15258_));
 sky130_fd_sc_hd__nand3_4 _45812_ (.A(_15248_),
    .B(_15257_),
    .C(_15258_),
    .Y(_15259_));
 sky130_fd_sc_hd__nand2_4 _45813_ (.A(_15257_),
    .B(_15258_),
    .Y(_15260_));
 sky130_fd_sc_hd__nand2_4 _45814_ (.A(_15260_),
    .B(_15247_),
    .Y(_15261_));
 sky130_fd_sc_hd__nand2_4 _45815_ (.A(_11910_),
    .B(_10513_),
    .Y(_15262_));
 sky130_fd_sc_hd__buf_1 _45816_ (.A(_03613_),
    .X(_15263_));
 sky130_fd_sc_hd__nand2_4 _45817_ (.A(_13054_),
    .B(_15263_),
    .Y(_15264_));
 sky130_fd_sc_hd__nand2_4 _45818_ (.A(_11022_),
    .B(_03607_),
    .Y(_15265_));
 sky130_fd_sc_hd__nand2_4 _45819_ (.A(_15264_),
    .B(_15265_),
    .Y(_15266_));
 sky130_fd_sc_hd__buf_1 _45820_ (.A(_12406_),
    .X(_15267_));
 sky130_fd_sc_hd__buf_1 _45821_ (.A(_12404_),
    .X(_15268_));
 sky130_fd_sc_hd__nand4_4 _45822_ (.A(_13054_),
    .B(_11022_),
    .C(_15267_),
    .D(_15268_),
    .Y(_15269_));
 sky130_fd_sc_hd__nand2_4 _45823_ (.A(_15266_),
    .B(_15269_),
    .Y(_15270_));
 sky130_fd_sc_hd__xor2_4 _45824_ (.A(_15262_),
    .B(_15270_),
    .X(_15271_));
 sky130_fd_sc_hd__a21o_4 _45825_ (.A1(_15259_),
    .A2(_15261_),
    .B1(_15271_),
    .X(_15272_));
 sky130_fd_sc_hd__nand3_4 _45826_ (.A(_15259_),
    .B(_15261_),
    .C(_15271_),
    .Y(_15273_));
 sky130_fd_sc_hd__nand2_4 _45827_ (.A(_15272_),
    .B(_15273_),
    .Y(_15274_));
 sky130_vsdinv _45828_ (.A(_15043_),
    .Y(_15275_));
 sky130_fd_sc_hd__a21oi_4 _45829_ (.A1(_15041_),
    .A2(_15054_),
    .B1(_15275_),
    .Y(_15276_));
 sky130_fd_sc_hd__nand2_4 _45830_ (.A(_15274_),
    .B(_15276_),
    .Y(_15277_));
 sky130_vsdinv _45831_ (.A(_15276_),
    .Y(_15278_));
 sky130_fd_sc_hd__nand3_4 _45832_ (.A(_15278_),
    .B(_15272_),
    .C(_15273_),
    .Y(_15279_));
 sky130_fd_sc_hd__nand2_4 _45833_ (.A(_15277_),
    .B(_15279_),
    .Y(_15280_));
 sky130_fd_sc_hd__a21boi_4 _45834_ (.A1(_15047_),
    .A2(_15050_),
    .B1_N(_15048_),
    .Y(_15281_));
 sky130_fd_sc_hd__nand2_4 _45835_ (.A(_13342_),
    .B(_13298_),
    .Y(_15282_));
 sky130_fd_sc_hd__nand2_4 _45836_ (.A(_09830_),
    .B(_12427_),
    .Y(_15283_));
 sky130_fd_sc_hd__nand2_4 _45837_ (.A(_15282_),
    .B(_15283_),
    .Y(_15284_));
 sky130_fd_sc_hd__nand4_4 _45838_ (.A(_08528_),
    .B(_08531_),
    .C(_12430_),
    .D(_12115_),
    .Y(_15285_));
 sky130_fd_sc_hd__nand2_4 _45839_ (.A(_11249_),
    .B(_13303_),
    .Y(_15286_));
 sky130_vsdinv _45840_ (.A(_15286_),
    .Y(_15287_));
 sky130_fd_sc_hd__a21o_4 _45841_ (.A1(_15284_),
    .A2(_15285_),
    .B1(_15287_),
    .X(_15288_));
 sky130_fd_sc_hd__nand3_4 _45842_ (.A(_15284_),
    .B(_15285_),
    .C(_15287_),
    .Y(_15289_));
 sky130_fd_sc_hd__nand2_4 _45843_ (.A(_15288_),
    .B(_15289_),
    .Y(_15290_));
 sky130_fd_sc_hd__nor2_4 _45844_ (.A(_15281_),
    .B(_15290_),
    .Y(_15291_));
 sky130_vsdinv _45845_ (.A(_15291_),
    .Y(_15292_));
 sky130_fd_sc_hd__nand2_4 _45846_ (.A(_15290_),
    .B(_15281_),
    .Y(_15293_));
 sky130_fd_sc_hd__a21boi_4 _45847_ (.A1(_15066_),
    .A2(_15069_),
    .B1_N(_15067_),
    .Y(_15294_));
 sky130_vsdinv _45848_ (.A(_15294_),
    .Y(_15295_));
 sky130_fd_sc_hd__a21oi_4 _45849_ (.A1(_15292_),
    .A2(_15293_),
    .B1(_15295_),
    .Y(_15296_));
 sky130_fd_sc_hd__nand3_4 _45850_ (.A(_15292_),
    .B(_15295_),
    .C(_15293_),
    .Y(_15297_));
 sky130_vsdinv _45851_ (.A(_15297_),
    .Y(_15298_));
 sky130_fd_sc_hd__nor2_4 _45852_ (.A(_15296_),
    .B(_15298_),
    .Y(_15299_));
 sky130_vsdinv _45853_ (.A(_15299_),
    .Y(_15300_));
 sky130_fd_sc_hd__nand2_4 _45854_ (.A(_15280_),
    .B(_15300_),
    .Y(_15301_));
 sky130_fd_sc_hd__nand3_4 _45855_ (.A(_15277_),
    .B(_15279_),
    .C(_15299_),
    .Y(_15302_));
 sky130_fd_sc_hd__nand2_4 _45856_ (.A(_15301_),
    .B(_15302_),
    .Y(_15303_));
 sky130_fd_sc_hd__a21boi_4 _45857_ (.A1(_15060_),
    .A2(_15082_),
    .B1_N(_15062_),
    .Y(_15304_));
 sky130_fd_sc_hd__nand2_4 _45858_ (.A(_15303_),
    .B(_15304_),
    .Y(_15305_));
 sky130_vsdinv _45859_ (.A(_15304_),
    .Y(_15306_));
 sky130_fd_sc_hd__nand3_4 _45860_ (.A(_15306_),
    .B(_15301_),
    .C(_15302_),
    .Y(_15307_));
 sky130_fd_sc_hd__nand2_4 _45861_ (.A(_15305_),
    .B(_15307_),
    .Y(_15308_));
 sky130_fd_sc_hd__a21boi_4 _45862_ (.A1(_15094_),
    .A2(_15097_),
    .B1_N(_15095_),
    .Y(_15309_));
 sky130_fd_sc_hd__nand2_4 _45863_ (.A(_12530_),
    .B(_12467_),
    .Y(_15310_));
 sky130_fd_sc_hd__nand2_4 _45864_ (.A(_13112_),
    .B(_03570_),
    .Y(_15311_));
 sky130_fd_sc_hd__nand2_4 _45865_ (.A(_15310_),
    .B(_15311_),
    .Y(_15312_));
 sky130_fd_sc_hd__nand4_4 _45866_ (.A(_13943_),
    .B(_12821_),
    .C(_08632_),
    .D(_14377_),
    .Y(_15313_));
 sky130_fd_sc_hd__nand2_4 _45867_ (.A(_11949_),
    .B(_13872_),
    .Y(_15314_));
 sky130_vsdinv _45868_ (.A(_15314_),
    .Y(_15315_));
 sky130_fd_sc_hd__a21o_4 _45869_ (.A1(_15312_),
    .A2(_15313_),
    .B1(_15315_),
    .X(_15316_));
 sky130_fd_sc_hd__nand3_4 _45870_ (.A(_15312_),
    .B(_15313_),
    .C(_15315_),
    .Y(_15317_));
 sky130_fd_sc_hd__nand2_4 _45871_ (.A(_15316_),
    .B(_15317_),
    .Y(_15318_));
 sky130_fd_sc_hd__nor2_4 _45872_ (.A(_15309_),
    .B(_15318_),
    .Y(_15319_));
 sky130_vsdinv _45873_ (.A(_15319_),
    .Y(_15320_));
 sky130_fd_sc_hd__nand2_4 _45874_ (.A(_15318_),
    .B(_15309_),
    .Y(_15321_));
 sky130_fd_sc_hd__nand2_4 _45875_ (.A(_15136_),
    .B(_11514_),
    .Y(_15322_));
 sky130_fd_sc_hd__nand2_4 _45876_ (.A(_14882_),
    .B(_13055_),
    .Y(_15323_));
 sky130_fd_sc_hd__nand2_4 _45877_ (.A(_12279_),
    .B(_11521_),
    .Y(_15324_));
 sky130_fd_sc_hd__xnor2_4 _45878_ (.A(_15323_),
    .B(_15324_),
    .Y(_15325_));
 sky130_fd_sc_hd__xor2_4 _45879_ (.A(_15322_),
    .B(_15325_),
    .X(_15326_));
 sky130_fd_sc_hd__a21o_4 _45880_ (.A1(_15320_),
    .A2(_15321_),
    .B1(_15326_),
    .X(_15327_));
 sky130_fd_sc_hd__nand3_4 _45881_ (.A(_15326_),
    .B(_15321_),
    .C(_15320_),
    .Y(_15328_));
 sky130_fd_sc_hd__o21a_4 _45882_ (.A1(_15077_),
    .A2(_15073_),
    .B1(_15076_),
    .X(_15329_));
 sky130_vsdinv _45883_ (.A(_15329_),
    .Y(_15330_));
 sky130_fd_sc_hd__a21o_4 _45884_ (.A1(_15327_),
    .A2(_15328_),
    .B1(_15330_),
    .X(_15331_));
 sky130_fd_sc_hd__nand3_4 _45885_ (.A(_15327_),
    .B(_15330_),
    .C(_15328_),
    .Y(_15332_));
 sky130_fd_sc_hd__a21boi_4 _45886_ (.A1(_15107_),
    .A2(_15102_),
    .B1_N(_15101_),
    .Y(_15333_));
 sky130_vsdinv _45887_ (.A(_15333_),
    .Y(_15334_));
 sky130_fd_sc_hd__a21oi_4 _45888_ (.A1(_15331_),
    .A2(_15332_),
    .B1(_15334_),
    .Y(_15335_));
 sky130_vsdinv _45889_ (.A(_15335_),
    .Y(_15336_));
 sky130_fd_sc_hd__nand3_4 _45890_ (.A(_15331_),
    .B(_15334_),
    .C(_15332_),
    .Y(_15337_));
 sky130_fd_sc_hd__nand2_4 _45891_ (.A(_15336_),
    .B(_15337_),
    .Y(_15338_));
 sky130_fd_sc_hd__nand2_4 _45892_ (.A(_15308_),
    .B(_15338_),
    .Y(_15339_));
 sky130_vsdinv _45893_ (.A(_15337_),
    .Y(_15340_));
 sky130_fd_sc_hd__nor2_4 _45894_ (.A(_15335_),
    .B(_15340_),
    .Y(_15341_));
 sky130_fd_sc_hd__nand3_4 _45895_ (.A(_15341_),
    .B(_15307_),
    .C(_15305_),
    .Y(_15342_));
 sky130_fd_sc_hd__nand2_4 _45896_ (.A(_15339_),
    .B(_15342_),
    .Y(_15343_));
 sky130_vsdinv _45897_ (.A(_15090_),
    .Y(_15344_));
 sky130_fd_sc_hd__a21oi_4 _45898_ (.A1(_15122_),
    .A2(_15088_),
    .B1(_15344_),
    .Y(_15345_));
 sky130_fd_sc_hd__nand2_4 _45899_ (.A(_15343_),
    .B(_15345_),
    .Y(_15346_));
 sky130_fd_sc_hd__a21o_4 _45900_ (.A1(_15122_),
    .A2(_15088_),
    .B1(_15344_),
    .X(_15347_));
 sky130_fd_sc_hd__nand3_4 _45901_ (.A(_15347_),
    .B(_15339_),
    .C(_15342_),
    .Y(_15348_));
 sky130_fd_sc_hd__nand2_4 _45902_ (.A(_15346_),
    .B(_15348_),
    .Y(_15349_));
 sky130_vsdinv _45903_ (.A(_15113_),
    .Y(_15350_));
 sky130_fd_sc_hd__a21oi_4 _45904_ (.A1(_15112_),
    .A2(_15115_),
    .B1(_15350_),
    .Y(_15351_));
 sky130_vsdinv _45905_ (.A(_15351_),
    .Y(_15352_));
 sky130_fd_sc_hd__maj3_4 _45906_ (.A(_15104_),
    .B(_15105_),
    .C(_15103_),
    .X(_15353_));
 sky130_fd_sc_hd__nand2_4 _45907_ (.A(_11675_),
    .B(_07717_),
    .Y(_15354_));
 sky130_fd_sc_hd__nand2_4 _45908_ (.A(_11684_),
    .B(_03536_),
    .Y(_15355_));
 sky130_fd_sc_hd__nand2_4 _45909_ (.A(_15354_),
    .B(_15355_),
    .Y(_15356_));
 sky130_fd_sc_hd__nand4_4 _45910_ (.A(_11989_),
    .B(_11991_),
    .C(_07554_),
    .D(_07557_),
    .Y(_15357_));
 sky130_fd_sc_hd__nand2_4 _45911_ (.A(_03405_),
    .B(_07561_),
    .Y(_15358_));
 sky130_vsdinv _45912_ (.A(_15358_),
    .Y(_15359_));
 sky130_fd_sc_hd__buf_1 _45913_ (.A(_15359_),
    .X(_15360_));
 sky130_fd_sc_hd__a21o_4 _45914_ (.A1(_15356_),
    .A2(_15357_),
    .B1(_15360_),
    .X(_15361_));
 sky130_fd_sc_hd__nand3_4 _45915_ (.A(_15356_),
    .B(_15357_),
    .C(_15360_),
    .Y(_15362_));
 sky130_fd_sc_hd__nand2_4 _45916_ (.A(_15361_),
    .B(_15362_),
    .Y(_15363_));
 sky130_fd_sc_hd__nor2_4 _45917_ (.A(_15353_),
    .B(_15363_),
    .Y(_15364_));
 sky130_vsdinv _45918_ (.A(_15364_),
    .Y(_15365_));
 sky130_fd_sc_hd__nand2_4 _45919_ (.A(_15363_),
    .B(_15353_),
    .Y(_15366_));
 sky130_fd_sc_hd__a21boi_4 _45920_ (.A1(_15135_),
    .A2(_15139_),
    .B1_N(_15137_),
    .Y(_15367_));
 sky130_vsdinv _45921_ (.A(_15367_),
    .Y(_15368_));
 sky130_fd_sc_hd__a21o_4 _45922_ (.A1(_15365_),
    .A2(_15366_),
    .B1(_15368_),
    .X(_15369_));
 sky130_fd_sc_hd__nand3_4 _45923_ (.A(_15365_),
    .B(_15368_),
    .C(_15366_),
    .Y(_15370_));
 sky130_fd_sc_hd__nand2_4 _45924_ (.A(_15369_),
    .B(_15370_),
    .Y(_15371_));
 sky130_fd_sc_hd__maj3_4 _45925_ (.A(_15146_),
    .B(_15142_),
    .C(_15144_),
    .X(_15372_));
 sky130_fd_sc_hd__nand2_4 _45926_ (.A(_15371_),
    .B(_15372_),
    .Y(_15373_));
 sky130_fd_sc_hd__nand4_4 _45927_ (.A(_03407_),
    .B(_08598_),
    .C(_11907_),
    .D(_12221_),
    .Y(_15374_));
 sky130_fd_sc_hd__o21a_4 _45928_ (.A1(_14688_),
    .A2(_15154_),
    .B1(_15374_),
    .X(_15375_));
 sky130_fd_sc_hd__a21o_4 _45929_ (.A1(_14459_),
    .A2(_14460_),
    .B1(_15375_),
    .X(_15376_));
 sky130_fd_sc_hd__nand3_4 _45930_ (.A(_14459_),
    .B(_14460_),
    .C(_15375_),
    .Y(_15377_));
 sky130_fd_sc_hd__and2_4 _45931_ (.A(_15376_),
    .B(_15377_),
    .X(_15378_));
 sky130_fd_sc_hd__buf_1 _45932_ (.A(_15378_),
    .X(_15379_));
 sky130_vsdinv _45933_ (.A(_15372_),
    .Y(_15380_));
 sky130_fd_sc_hd__nand3_4 _45934_ (.A(_15369_),
    .B(_15380_),
    .C(_15370_),
    .Y(_15381_));
 sky130_fd_sc_hd__nand3_4 _45935_ (.A(_15373_),
    .B(_15379_),
    .C(_15381_),
    .Y(_15382_));
 sky130_fd_sc_hd__buf_1 _45936_ (.A(_15378_),
    .X(_15383_));
 sky130_fd_sc_hd__a21o_4 _45937_ (.A1(_15373_),
    .A2(_15381_),
    .B1(_15383_),
    .X(_15384_));
 sky130_fd_sc_hd__nand3_4 _45938_ (.A(_15352_),
    .B(_15382_),
    .C(_15384_),
    .Y(_15385_));
 sky130_fd_sc_hd__nand2_4 _45939_ (.A(_15384_),
    .B(_15382_),
    .Y(_15386_));
 sky130_fd_sc_hd__nand2_4 _45940_ (.A(_15386_),
    .B(_15351_),
    .Y(_15387_));
 sky130_fd_sc_hd__a21boi_4 _45941_ (.A1(_15152_),
    .A2(_15163_),
    .B1_N(_15153_),
    .Y(_15388_));
 sky130_vsdinv _45942_ (.A(_15388_),
    .Y(_15389_));
 sky130_fd_sc_hd__a21oi_4 _45943_ (.A1(_15385_),
    .A2(_15387_),
    .B1(_15389_),
    .Y(_15390_));
 sky130_vsdinv _45944_ (.A(_15390_),
    .Y(_15391_));
 sky130_fd_sc_hd__nand3_4 _45945_ (.A(_15385_),
    .B(_15387_),
    .C(_15389_),
    .Y(_15392_));
 sky130_fd_sc_hd__nand2_4 _45946_ (.A(_15391_),
    .B(_15392_),
    .Y(_15393_));
 sky130_fd_sc_hd__nand2_4 _45947_ (.A(_15349_),
    .B(_15393_),
    .Y(_15394_));
 sky130_vsdinv _45948_ (.A(_15392_),
    .Y(_15395_));
 sky130_fd_sc_hd__nor2_4 _45949_ (.A(_15390_),
    .B(_15395_),
    .Y(_15396_));
 sky130_fd_sc_hd__nand3_4 _45950_ (.A(_15396_),
    .B(_15346_),
    .C(_15348_),
    .Y(_15397_));
 sky130_fd_sc_hd__nand2_4 _45951_ (.A(_15394_),
    .B(_15397_),
    .Y(_15398_));
 sky130_fd_sc_hd__a21oi_4 _45952_ (.A1(_15120_),
    .A2(_15123_),
    .B1(_15127_),
    .Y(_15399_));
 sky130_fd_sc_hd__o21a_4 _45953_ (.A1(_15399_),
    .A2(_15175_),
    .B1(_15128_),
    .X(_15400_));
 sky130_fd_sc_hd__nand2_4 _45954_ (.A(_15398_),
    .B(_15400_),
    .Y(_15401_));
 sky130_fd_sc_hd__o21ai_4 _45955_ (.A1(_15399_),
    .A2(_15175_),
    .B1(_15128_),
    .Y(_15402_));
 sky130_fd_sc_hd__nand3_4 _45956_ (.A(_15402_),
    .B(_15394_),
    .C(_15397_),
    .Y(_15403_));
 sky130_fd_sc_hd__nand2_4 _45957_ (.A(_15401_),
    .B(_15403_),
    .Y(_15404_));
 sky130_fd_sc_hd__nand2_4 _45958_ (.A(_15162_),
    .B(_14463_),
    .Y(_15405_));
 sky130_fd_sc_hd__a21o_4 _45959_ (.A1(_15405_),
    .A2(_15374_),
    .B1(_14732_),
    .X(_15406_));
 sky130_fd_sc_hd__nand3_4 _45960_ (.A(_14968_),
    .B(_15405_),
    .C(_15374_),
    .Y(_15407_));
 sky130_fd_sc_hd__nand2_4 _45961_ (.A(_15406_),
    .B(_15407_),
    .Y(_15408_));
 sky130_fd_sc_hd__nand2_4 _45962_ (.A(_15408_),
    .B(_14976_),
    .Y(_15409_));
 sky130_fd_sc_hd__buf_1 _45963_ (.A(_14977_),
    .X(_15410_));
 sky130_fd_sc_hd__nand3_4 _45964_ (.A(_15406_),
    .B(_15407_),
    .C(_15410_),
    .Y(_15411_));
 sky130_fd_sc_hd__nand2_4 _45965_ (.A(_15409_),
    .B(_15411_),
    .Y(_15412_));
 sky130_fd_sc_hd__maj3_4 _45966_ (.A(_14976_),
    .B(_14735_),
    .C(_15186_),
    .X(_15413_));
 sky130_fd_sc_hd__nand2_4 _45967_ (.A(_15412_),
    .B(_15413_),
    .Y(_15414_));
 sky130_vsdinv _45968_ (.A(_15413_),
    .Y(_15415_));
 sky130_fd_sc_hd__nand3_4 _45969_ (.A(_15415_),
    .B(_15411_),
    .C(_15409_),
    .Y(_15416_));
 sky130_fd_sc_hd__a21o_4 _45970_ (.A1(_15414_),
    .A2(_15416_),
    .B1(_13483_),
    .X(_15417_));
 sky130_fd_sc_hd__nand3_4 _45971_ (.A(_15414_),
    .B(_15416_),
    .C(_14273_),
    .Y(_15418_));
 sky130_fd_sc_hd__nand2_4 _45972_ (.A(_15417_),
    .B(_15418_),
    .Y(_15419_));
 sky130_fd_sc_hd__o21ai_4 _45973_ (.A1(_15170_),
    .A2(_15167_),
    .B1(_15168_),
    .Y(_15420_));
 sky130_vsdinv _45974_ (.A(_15420_),
    .Y(_15421_));
 sky130_fd_sc_hd__nand2_4 _45975_ (.A(_15419_),
    .B(_15421_),
    .Y(_15422_));
 sky130_fd_sc_hd__nand3_4 _45976_ (.A(_15420_),
    .B(_15417_),
    .C(_15418_),
    .Y(_15423_));
 sky130_fd_sc_hd__nand2_4 _45977_ (.A(_15422_),
    .B(_15423_),
    .Y(_15424_));
 sky130_fd_sc_hd__a21boi_4 _45978_ (.A1(_15192_),
    .A2(_13756_),
    .B1_N(_15194_),
    .Y(_15425_));
 sky130_fd_sc_hd__nand2_4 _45979_ (.A(_15424_),
    .B(_15425_),
    .Y(_15426_));
 sky130_vsdinv _45980_ (.A(_15425_),
    .Y(_15427_));
 sky130_fd_sc_hd__nand3_4 _45981_ (.A(_15422_),
    .B(_15427_),
    .C(_15423_),
    .Y(_15428_));
 sky130_fd_sc_hd__nand2_4 _45982_ (.A(_15426_),
    .B(_15428_),
    .Y(_15429_));
 sky130_fd_sc_hd__nand2_4 _45983_ (.A(_15404_),
    .B(_15429_),
    .Y(_15430_));
 sky130_vsdinv _45984_ (.A(_15429_),
    .Y(_15431_));
 sky130_fd_sc_hd__nand3_4 _45985_ (.A(_15431_),
    .B(_15403_),
    .C(_15401_),
    .Y(_15432_));
 sky130_fd_sc_hd__nand2_4 _45986_ (.A(_15430_),
    .B(_15432_),
    .Y(_15433_));
 sky130_fd_sc_hd__a21boi_4 _45987_ (.A1(_15212_),
    .A2(_15181_),
    .B1_N(_15183_),
    .Y(_15434_));
 sky130_fd_sc_hd__nand2_4 _45988_ (.A(_15433_),
    .B(_15434_),
    .Y(_15435_));
 sky130_vsdinv _45989_ (.A(_15181_),
    .Y(_15436_));
 sky130_fd_sc_hd__o21ai_4 _45990_ (.A1(_15208_),
    .A2(_15436_),
    .B1(_15183_),
    .Y(_15437_));
 sky130_fd_sc_hd__nand3_4 _45991_ (.A(_15437_),
    .B(_15430_),
    .C(_15432_),
    .Y(_15438_));
 sky130_fd_sc_hd__nand2_4 _45992_ (.A(_15435_),
    .B(_15438_),
    .Y(_15439_));
 sky130_fd_sc_hd__buf_8 _45993_ (.A(_13776_),
    .X(_15440_));
 sky130_fd_sc_hd__a21boi_4 _45994_ (.A1(_15200_),
    .A2(_15205_),
    .B1_N(_15203_),
    .Y(_15441_));
 sky130_fd_sc_hd__xor2_4 _45995_ (.A(_15440_),
    .B(_15441_),
    .X(_15442_));
 sky130_fd_sc_hd__nand2_4 _45996_ (.A(_15439_),
    .B(_15442_),
    .Y(_15443_));
 sky130_vsdinv _45997_ (.A(_15442_),
    .Y(_15444_));
 sky130_fd_sc_hd__nand3_4 _45998_ (.A(_15435_),
    .B(_15438_),
    .C(_15444_),
    .Y(_15445_));
 sky130_fd_sc_hd__nand2_4 _45999_ (.A(_15443_),
    .B(_15445_),
    .Y(_15446_));
 sky130_fd_sc_hd__nand2_4 _46000_ (.A(_15225_),
    .B(_15219_),
    .Y(_15447_));
 sky130_vsdinv _46001_ (.A(_15447_),
    .Y(_15448_));
 sky130_fd_sc_hd__nand2_4 _46002_ (.A(_15446_),
    .B(_15448_),
    .Y(_15449_));
 sky130_fd_sc_hd__nand3_4 _46003_ (.A(_15447_),
    .B(_15443_),
    .C(_15445_),
    .Y(_15450_));
 sky130_fd_sc_hd__nand2_4 _46004_ (.A(_15449_),
    .B(_15450_),
    .Y(_15451_));
 sky130_fd_sc_hd__buf_1 _46005_ (.A(_14303_),
    .X(_15452_));
 sky130_fd_sc_hd__a21oi_4 _46006_ (.A1(_14997_),
    .A2(_14992_),
    .B1(_15452_),
    .Y(_15453_));
 sky130_vsdinv _46007_ (.A(_15453_),
    .Y(_15454_));
 sky130_fd_sc_hd__nand2_4 _46008_ (.A(_15451_),
    .B(_15454_),
    .Y(_15455_));
 sky130_fd_sc_hd__nand3_4 _46009_ (.A(_15449_),
    .B(_15453_),
    .C(_15450_),
    .Y(_15456_));
 sky130_fd_sc_hd__nand2_4 _46010_ (.A(_15455_),
    .B(_15456_),
    .Y(_15457_));
 sky130_fd_sc_hd__nand2_4 _46011_ (.A(_15235_),
    .B(_15230_),
    .Y(_15458_));
 sky130_vsdinv _46012_ (.A(_15458_),
    .Y(_15459_));
 sky130_fd_sc_hd__nand2_4 _46013_ (.A(_15457_),
    .B(_15459_),
    .Y(_15460_));
 sky130_fd_sc_hd__nand3_4 _46014_ (.A(_15458_),
    .B(_15455_),
    .C(_15456_),
    .Y(_15461_));
 sky130_fd_sc_hd__nand2_4 _46015_ (.A(_15460_),
    .B(_15461_),
    .Y(_15462_));
 sky130_vsdinv _46016_ (.A(_15240_),
    .Y(_15463_));
 sky130_fd_sc_hd__a21oi_4 _46017_ (.A1(_15246_),
    .A2(_15238_),
    .B1(_15463_),
    .Y(_15464_));
 sky130_fd_sc_hd__xor2_4 _46018_ (.A(_15462_),
    .B(_15464_),
    .X(_01452_));
 sky130_fd_sc_hd__buf_1 _46019_ (.A(_10958_),
    .X(_15465_));
 sky130_fd_sc_hd__nand2_4 _46020_ (.A(_14096_),
    .B(_15465_),
    .Y(_15466_));
 sky130_fd_sc_hd__o21ai_4 _46021_ (.A1(_07625_),
    .A2(_13808_),
    .B1(_15466_),
    .Y(_15467_));
 sky130_fd_sc_hd__nand4_4 _46022_ (.A(_03326_),
    .B(_11014_),
    .C(_15465_),
    .D(_11384_),
    .Y(_15468_));
 sky130_fd_sc_hd__nand2_4 _46023_ (.A(_11871_),
    .B(_03620_),
    .Y(_15469_));
 sky130_vsdinv _46024_ (.A(_15469_),
    .Y(_15470_));
 sky130_fd_sc_hd__a21o_4 _46025_ (.A1(_15467_),
    .A2(_15468_),
    .B1(_15470_),
    .X(_15471_));
 sky130_fd_sc_hd__nand3_4 _46026_ (.A(_15467_),
    .B(_15468_),
    .C(_15470_),
    .Y(_15472_));
 sky130_fd_sc_hd__nand2_4 _46027_ (.A(_15471_),
    .B(_15472_),
    .Y(_15473_));
 sky130_fd_sc_hd__a21o_4 _46028_ (.A1(_15254_),
    .A2(_15258_),
    .B1(_15473_),
    .X(_15474_));
 sky130_fd_sc_hd__nand3_4 _46029_ (.A(_15473_),
    .B(_15254_),
    .C(_15258_),
    .Y(_15475_));
 sky130_fd_sc_hd__nand2_4 _46030_ (.A(_08528_),
    .B(_10509_),
    .Y(_15476_));
 sky130_fd_sc_hd__nand2_4 _46031_ (.A(_13051_),
    .B(_15263_),
    .Y(_15477_));
 sky130_fd_sc_hd__buf_1 _46032_ (.A(_11776_),
    .X(_15478_));
 sky130_fd_sc_hd__nand2_4 _46033_ (.A(_11904_),
    .B(_15478_),
    .Y(_15479_));
 sky130_fd_sc_hd__nand2_4 _46034_ (.A(_15477_),
    .B(_15479_),
    .Y(_15480_));
 sky130_fd_sc_hd__nand4_4 _46035_ (.A(_13051_),
    .B(_11243_),
    .C(_03607_),
    .D(_15263_),
    .Y(_15481_));
 sky130_fd_sc_hd__nand2_4 _46036_ (.A(_15480_),
    .B(_15481_),
    .Y(_15482_));
 sky130_fd_sc_hd__xor2_4 _46037_ (.A(_15476_),
    .B(_15482_),
    .X(_15483_));
 sky130_fd_sc_hd__a21o_4 _46038_ (.A1(_15474_),
    .A2(_15475_),
    .B1(_15483_),
    .X(_15484_));
 sky130_fd_sc_hd__nand3_4 _46039_ (.A(_15474_),
    .B(_15475_),
    .C(_15483_),
    .Y(_15485_));
 sky130_fd_sc_hd__nand2_4 _46040_ (.A(_15484_),
    .B(_15485_),
    .Y(_15486_));
 sky130_fd_sc_hd__a21o_4 _46041_ (.A1(_15259_),
    .A2(_15273_),
    .B1(_15486_),
    .X(_15487_));
 sky130_fd_sc_hd__nand3_4 _46042_ (.A(_15486_),
    .B(_15259_),
    .C(_15273_),
    .Y(_15488_));
 sky130_fd_sc_hd__a21boi_4 _46043_ (.A1(_15284_),
    .A2(_15287_),
    .B1_N(_15285_),
    .Y(_15489_));
 sky130_vsdinv _46044_ (.A(_15262_),
    .Y(_15490_));
 sky130_fd_sc_hd__a21boi_4 _46045_ (.A1(_15266_),
    .A2(_15490_),
    .B1_N(_15269_),
    .Y(_15491_));
 sky130_fd_sc_hd__nand2_4 _46046_ (.A(_12533_),
    .B(_03583_),
    .Y(_15492_));
 sky130_vsdinv _46047_ (.A(_15492_),
    .Y(_15493_));
 sky130_fd_sc_hd__buf_1 _46048_ (.A(_10305_),
    .X(_15494_));
 sky130_fd_sc_hd__nand2_4 _46049_ (.A(_13088_),
    .B(_15494_),
    .Y(_15495_));
 sky130_fd_sc_hd__buf_1 _46050_ (.A(_09831_),
    .X(_15496_));
 sky130_fd_sc_hd__nand2_4 _46051_ (.A(_15496_),
    .B(_03588_),
    .Y(_15497_));
 sky130_fd_sc_hd__nand2_4 _46052_ (.A(_15495_),
    .B(_15497_),
    .Y(_15498_));
 sky130_fd_sc_hd__buf_1 _46053_ (.A(_12431_),
    .X(_15499_));
 sky130_fd_sc_hd__nand4_4 _46054_ (.A(_14140_),
    .B(_14137_),
    .C(_13842_),
    .D(_15499_),
    .Y(_15500_));
 sky130_fd_sc_hd__nand2_4 _46055_ (.A(_15498_),
    .B(_15500_),
    .Y(_15501_));
 sky130_fd_sc_hd__xor2_4 _46056_ (.A(_15493_),
    .B(_15501_),
    .X(_15502_));
 sky130_fd_sc_hd__xnor2_4 _46057_ (.A(_15491_),
    .B(_15502_),
    .Y(_15503_));
 sky130_fd_sc_hd__xor2_4 _46058_ (.A(_15489_),
    .B(_15503_),
    .X(_15504_));
 sky130_fd_sc_hd__a21o_4 _46059_ (.A1(_15487_),
    .A2(_15488_),
    .B1(_15504_),
    .X(_15505_));
 sky130_fd_sc_hd__nand3_4 _46060_ (.A(_15487_),
    .B(_15504_),
    .C(_15488_),
    .Y(_15506_));
 sky130_fd_sc_hd__nand2_4 _46061_ (.A(_15505_),
    .B(_15506_),
    .Y(_15507_));
 sky130_fd_sc_hd__a21boi_4 _46062_ (.A1(_15277_),
    .A2(_15299_),
    .B1_N(_15279_),
    .Y(_15508_));
 sky130_fd_sc_hd__nand2_4 _46063_ (.A(_15507_),
    .B(_15508_),
    .Y(_15509_));
 sky130_vsdinv _46064_ (.A(_15508_),
    .Y(_15510_));
 sky130_fd_sc_hd__nand3_4 _46065_ (.A(_15505_),
    .B(_15510_),
    .C(_15506_),
    .Y(_15511_));
 sky130_fd_sc_hd__a21boi_4 _46066_ (.A1(_15312_),
    .A2(_15315_),
    .B1_N(_15313_),
    .Y(_15512_));
 sky130_fd_sc_hd__nand2_4 _46067_ (.A(_11639_),
    .B(_11502_),
    .Y(_15513_));
 sky130_fd_sc_hd__o21ai_4 _46068_ (.A1(_03376_),
    .A2(_03577_),
    .B1(_15513_),
    .Y(_15514_));
 sky130_fd_sc_hd__nand4_4 _46069_ (.A(_11893_),
    .B(_10084_),
    .C(_08632_),
    .D(_11173_),
    .Y(_15515_));
 sky130_fd_sc_hd__nand2_4 _46070_ (.A(_11951_),
    .B(_03564_),
    .Y(_15516_));
 sky130_vsdinv _46071_ (.A(_15516_),
    .Y(_15517_));
 sky130_fd_sc_hd__a21o_4 _46072_ (.A1(_15514_),
    .A2(_15515_),
    .B1(_15517_),
    .X(_15518_));
 sky130_fd_sc_hd__nand3_4 _46073_ (.A(_15514_),
    .B(_15515_),
    .C(_15517_),
    .Y(_15519_));
 sky130_fd_sc_hd__nand2_4 _46074_ (.A(_15518_),
    .B(_15519_),
    .Y(_15520_));
 sky130_fd_sc_hd__nor2_4 _46075_ (.A(_15512_),
    .B(_15520_),
    .Y(_15521_));
 sky130_vsdinv _46076_ (.A(_15521_),
    .Y(_15522_));
 sky130_fd_sc_hd__nand2_4 _46077_ (.A(_15520_),
    .B(_15512_),
    .Y(_15523_));
 sky130_fd_sc_hd__nand2_4 _46078_ (.A(_13169_),
    .B(_07980_),
    .Y(_15524_));
 sky130_fd_sc_hd__nand2_4 _46079_ (.A(_14426_),
    .B(_11187_),
    .Y(_15525_));
 sky130_fd_sc_hd__nand2_4 _46080_ (.A(_15132_),
    .B(_11518_),
    .Y(_15526_));
 sky130_fd_sc_hd__xnor2_4 _46081_ (.A(_15525_),
    .B(_15526_),
    .Y(_15527_));
 sky130_fd_sc_hd__xor2_4 _46082_ (.A(_15524_),
    .B(_15527_),
    .X(_15528_));
 sky130_fd_sc_hd__a21o_4 _46083_ (.A1(_15522_),
    .A2(_15523_),
    .B1(_15528_),
    .X(_15529_));
 sky130_fd_sc_hd__nand3_4 _46084_ (.A(_15522_),
    .B(_15528_),
    .C(_15523_),
    .Y(_15530_));
 sky130_fd_sc_hd__nand2_4 _46085_ (.A(_15529_),
    .B(_15530_),
    .Y(_15531_));
 sky130_fd_sc_hd__a21o_4 _46086_ (.A1(_15292_),
    .A2(_15297_),
    .B1(_15531_),
    .X(_15532_));
 sky130_fd_sc_hd__nand3_4 _46087_ (.A(_15531_),
    .B(_15292_),
    .C(_15297_),
    .Y(_15533_));
 sky130_fd_sc_hd__a21oi_4 _46088_ (.A1(_15326_),
    .A2(_15321_),
    .B1(_15319_),
    .Y(_15534_));
 sky130_vsdinv _46089_ (.A(_15534_),
    .Y(_15535_));
 sky130_fd_sc_hd__a21o_4 _46090_ (.A1(_15532_),
    .A2(_15533_),
    .B1(_15535_),
    .X(_15536_));
 sky130_fd_sc_hd__nand3_4 _46091_ (.A(_15532_),
    .B(_15535_),
    .C(_15533_),
    .Y(_15537_));
 sky130_fd_sc_hd__nand2_4 _46092_ (.A(_15536_),
    .B(_15537_),
    .Y(_15538_));
 sky130_fd_sc_hd__a21bo_4 _46093_ (.A1(_15509_),
    .A2(_15511_),
    .B1_N(_15538_),
    .X(_15539_));
 sky130_fd_sc_hd__nand4_4 _46094_ (.A(_15537_),
    .B(_15509_),
    .C(_15536_),
    .D(_15511_),
    .Y(_15540_));
 sky130_fd_sc_hd__nand2_4 _46095_ (.A(_15539_),
    .B(_15540_),
    .Y(_15541_));
 sky130_fd_sc_hd__a21boi_4 _46096_ (.A1(_15341_),
    .A2(_15305_),
    .B1_N(_15307_),
    .Y(_15542_));
 sky130_fd_sc_hd__nand2_4 _46097_ (.A(_15541_),
    .B(_15542_),
    .Y(_15543_));
 sky130_vsdinv _46098_ (.A(_15542_),
    .Y(_15544_));
 sky130_fd_sc_hd__nand3_4 _46099_ (.A(_15539_),
    .B(_15544_),
    .C(_15540_),
    .Y(_15545_));
 sky130_fd_sc_hd__nand2_4 _46100_ (.A(_15543_),
    .B(_15545_),
    .Y(_15546_));
 sky130_fd_sc_hd__maj3_4 _46101_ (.A(_15323_),
    .B(_15324_),
    .C(_15322_),
    .X(_15547_));
 sky130_fd_sc_hd__nand2_4 _46102_ (.A(_11337_),
    .B(_13644_),
    .Y(_15548_));
 sky130_fd_sc_hd__nand2_4 _46103_ (.A(_11339_),
    .B(_08571_),
    .Y(_15549_));
 sky130_fd_sc_hd__nand2_4 _46104_ (.A(_15548_),
    .B(_15549_),
    .Y(_15550_));
 sky130_fd_sc_hd__nand4_4 _46105_ (.A(_10837_),
    .B(_03407_),
    .C(_13089_),
    .D(_12190_),
    .Y(_15551_));
 sky130_fd_sc_hd__a21o_4 _46106_ (.A1(_15550_),
    .A2(_15551_),
    .B1(_15360_),
    .X(_15552_));
 sky130_fd_sc_hd__buf_1 _46107_ (.A(_15360_),
    .X(_15553_));
 sky130_fd_sc_hd__nand3_4 _46108_ (.A(_15550_),
    .B(_15551_),
    .C(_15553_),
    .Y(_15554_));
 sky130_fd_sc_hd__nand2_4 _46109_ (.A(_15552_),
    .B(_15554_),
    .Y(_15555_));
 sky130_fd_sc_hd__or2_4 _46110_ (.A(_15547_),
    .B(_15555_),
    .X(_15556_));
 sky130_fd_sc_hd__nand2_4 _46111_ (.A(_15555_),
    .B(_15547_),
    .Y(_15557_));
 sky130_fd_sc_hd__a21boi_4 _46112_ (.A1(_15356_),
    .A2(_15553_),
    .B1_N(_15357_),
    .Y(_15558_));
 sky130_vsdinv _46113_ (.A(_15558_),
    .Y(_15559_));
 sky130_fd_sc_hd__a21o_4 _46114_ (.A1(_15556_),
    .A2(_15557_),
    .B1(_15559_),
    .X(_15560_));
 sky130_fd_sc_hd__nand3_4 _46115_ (.A(_15556_),
    .B(_15557_),
    .C(_15559_),
    .Y(_15561_));
 sky130_fd_sc_hd__a21oi_4 _46116_ (.A1(_15366_),
    .A2(_15368_),
    .B1(_15364_),
    .Y(_15562_));
 sky130_vsdinv _46117_ (.A(_15562_),
    .Y(_15563_));
 sky130_fd_sc_hd__a21o_4 _46118_ (.A1(_15560_),
    .A2(_15561_),
    .B1(_15563_),
    .X(_15564_));
 sky130_fd_sc_hd__nand3_4 _46119_ (.A(_15560_),
    .B(_15561_),
    .C(_15563_),
    .Y(_15565_));
 sky130_fd_sc_hd__a21o_4 _46120_ (.A1(_15564_),
    .A2(_15565_),
    .B1(_15383_),
    .X(_15566_));
 sky130_fd_sc_hd__nand3_4 _46121_ (.A(_15564_),
    .B(_15379_),
    .C(_15565_),
    .Y(_15567_));
 sky130_fd_sc_hd__nand2_4 _46122_ (.A(_15566_),
    .B(_15567_),
    .Y(_15568_));
 sky130_fd_sc_hd__a21o_4 _46123_ (.A1(_15332_),
    .A2(_15337_),
    .B1(_15568_),
    .X(_15569_));
 sky130_fd_sc_hd__nand3_4 _46124_ (.A(_15568_),
    .B(_15332_),
    .C(_15337_),
    .Y(_15570_));
 sky130_fd_sc_hd__buf_1 _46125_ (.A(_15383_),
    .X(_15571_));
 sky130_fd_sc_hd__a21boi_4 _46126_ (.A1(_15373_),
    .A2(_15571_),
    .B1_N(_15381_),
    .Y(_15572_));
 sky130_vsdinv _46127_ (.A(_15572_),
    .Y(_15573_));
 sky130_fd_sc_hd__a21o_4 _46128_ (.A1(_15569_),
    .A2(_15570_),
    .B1(_15573_),
    .X(_15574_));
 sky130_fd_sc_hd__nand3_4 _46129_ (.A(_15569_),
    .B(_15573_),
    .C(_15570_),
    .Y(_15575_));
 sky130_fd_sc_hd__nand2_4 _46130_ (.A(_15574_),
    .B(_15575_),
    .Y(_15576_));
 sky130_fd_sc_hd__nand2_4 _46131_ (.A(_15546_),
    .B(_15576_),
    .Y(_15577_));
 sky130_vsdinv _46132_ (.A(_15576_),
    .Y(_15578_));
 sky130_fd_sc_hd__nand3_4 _46133_ (.A(_15543_),
    .B(_15578_),
    .C(_15545_),
    .Y(_15579_));
 sky130_fd_sc_hd__nand2_4 _46134_ (.A(_15577_),
    .B(_15579_),
    .Y(_15580_));
 sky130_fd_sc_hd__a21boi_4 _46135_ (.A1(_15396_),
    .A2(_15346_),
    .B1_N(_15348_),
    .Y(_15581_));
 sky130_fd_sc_hd__nand2_4 _46136_ (.A(_15580_),
    .B(_15581_),
    .Y(_15582_));
 sky130_vsdinv _46137_ (.A(_15581_),
    .Y(_15583_));
 sky130_fd_sc_hd__nand3_4 _46138_ (.A(_15577_),
    .B(_15583_),
    .C(_15579_),
    .Y(_15584_));
 sky130_fd_sc_hd__nand2_4 _46139_ (.A(_15582_),
    .B(_15584_),
    .Y(_15585_));
 sky130_fd_sc_hd__and2_4 _46140_ (.A(_15377_),
    .B(_15374_),
    .X(_15586_));
 sky130_fd_sc_hd__nand2_4 _46141_ (.A(_14735_),
    .B(_15586_),
    .Y(_15587_));
 sky130_vsdinv _46142_ (.A(_15586_),
    .Y(_15588_));
 sky130_fd_sc_hd__nand3_4 _46143_ (.A(_15588_),
    .B(_14730_),
    .C(_14731_),
    .Y(_15589_));
 sky130_fd_sc_hd__nand3_4 _46144_ (.A(_15587_),
    .B(_15410_),
    .C(_15589_),
    .Y(_15590_));
 sky130_fd_sc_hd__a21o_4 _46145_ (.A1(_15587_),
    .A2(_15589_),
    .B1(_15410_),
    .X(_15591_));
 sky130_fd_sc_hd__a21boi_4 _46146_ (.A1(_15410_),
    .A2(_15407_),
    .B1_N(_15406_),
    .Y(_15592_));
 sky130_vsdinv _46147_ (.A(_15592_),
    .Y(_15593_));
 sky130_fd_sc_hd__a21o_4 _46148_ (.A1(_15590_),
    .A2(_15591_),
    .B1(_15593_),
    .X(_15594_));
 sky130_fd_sc_hd__nand3_4 _46149_ (.A(_15593_),
    .B(_15590_),
    .C(_15591_),
    .Y(_15595_));
 sky130_fd_sc_hd__a21o_4 _46150_ (.A1(_15594_),
    .A2(_15595_),
    .B1(_13483_),
    .X(_15596_));
 sky130_fd_sc_hd__nand3_4 _46151_ (.A(_15594_),
    .B(_14273_),
    .C(_15595_),
    .Y(_15597_));
 sky130_fd_sc_hd__a21boi_4 _46152_ (.A1(_15389_),
    .A2(_15387_),
    .B1_N(_15385_),
    .Y(_15598_));
 sky130_vsdinv _46153_ (.A(_15598_),
    .Y(_15599_));
 sky130_fd_sc_hd__a21o_4 _46154_ (.A1(_15596_),
    .A2(_15597_),
    .B1(_15599_),
    .X(_15600_));
 sky130_fd_sc_hd__nand3_4 _46155_ (.A(_15596_),
    .B(_15599_),
    .C(_15597_),
    .Y(_15601_));
 sky130_fd_sc_hd__a21boi_4 _46156_ (.A1(_15414_),
    .A2(_14757_),
    .B1_N(_15416_),
    .Y(_15602_));
 sky130_vsdinv _46157_ (.A(_15602_),
    .Y(_15603_));
 sky130_fd_sc_hd__a21o_4 _46158_ (.A1(_15600_),
    .A2(_15601_),
    .B1(_15603_),
    .X(_15604_));
 sky130_fd_sc_hd__nand3_4 _46159_ (.A(_15600_),
    .B(_15603_),
    .C(_15601_),
    .Y(_15605_));
 sky130_fd_sc_hd__nand2_4 _46160_ (.A(_15604_),
    .B(_15605_),
    .Y(_15606_));
 sky130_fd_sc_hd__nand2_4 _46161_ (.A(_15585_),
    .B(_15606_),
    .Y(_15607_));
 sky130_vsdinv _46162_ (.A(_15606_),
    .Y(_15608_));
 sky130_fd_sc_hd__nand3_4 _46163_ (.A(_15582_),
    .B(_15608_),
    .C(_15584_),
    .Y(_15609_));
 sky130_fd_sc_hd__nand2_4 _46164_ (.A(_15607_),
    .B(_15609_),
    .Y(_15610_));
 sky130_fd_sc_hd__a21boi_4 _46165_ (.A1(_15431_),
    .A2(_15401_),
    .B1_N(_15403_),
    .Y(_15611_));
 sky130_fd_sc_hd__nand2_4 _46166_ (.A(_15610_),
    .B(_15611_),
    .Y(_15612_));
 sky130_vsdinv _46167_ (.A(_15611_),
    .Y(_15613_));
 sky130_fd_sc_hd__nand3_4 _46168_ (.A(_15607_),
    .B(_15609_),
    .C(_15613_),
    .Y(_15614_));
 sky130_fd_sc_hd__nand2_4 _46169_ (.A(_15612_),
    .B(_15614_),
    .Y(_15615_));
 sky130_fd_sc_hd__a21boi_4 _46170_ (.A1(_15422_),
    .A2(_15427_),
    .B1_N(_15423_),
    .Y(_15616_));
 sky130_fd_sc_hd__xor2_4 _46171_ (.A(_15440_),
    .B(_15616_),
    .X(_15617_));
 sky130_fd_sc_hd__nand2_4 _46172_ (.A(_15615_),
    .B(_15617_),
    .Y(_15618_));
 sky130_vsdinv _46173_ (.A(_15617_),
    .Y(_15619_));
 sky130_fd_sc_hd__nand3_4 _46174_ (.A(_15612_),
    .B(_15619_),
    .C(_15614_),
    .Y(_15620_));
 sky130_fd_sc_hd__nand2_4 _46175_ (.A(_15618_),
    .B(_15620_),
    .Y(_15621_));
 sky130_fd_sc_hd__a21boi_4 _46176_ (.A1(_15435_),
    .A2(_15444_),
    .B1_N(_15438_),
    .Y(_15622_));
 sky130_fd_sc_hd__nand2_4 _46177_ (.A(_15621_),
    .B(_15622_),
    .Y(_15623_));
 sky130_vsdinv _46178_ (.A(_15622_),
    .Y(_15624_));
 sky130_fd_sc_hd__nand3_4 _46179_ (.A(_15618_),
    .B(_15620_),
    .C(_15624_),
    .Y(_15625_));
 sky130_fd_sc_hd__nand2_4 _46180_ (.A(_15623_),
    .B(_15625_),
    .Y(_15626_));
 sky130_fd_sc_hd__buf_1 _46181_ (.A(_14050_),
    .X(_15627_));
 sky130_fd_sc_hd__a21oi_4 _46182_ (.A1(_15207_),
    .A2(_15203_),
    .B1(_15627_),
    .Y(_15628_));
 sky130_vsdinv _46183_ (.A(_15628_),
    .Y(_15629_));
 sky130_fd_sc_hd__nand2_4 _46184_ (.A(_15626_),
    .B(_15629_),
    .Y(_15630_));
 sky130_fd_sc_hd__nand3_4 _46185_ (.A(_15623_),
    .B(_15628_),
    .C(_15625_),
    .Y(_15631_));
 sky130_fd_sc_hd__nand2_4 _46186_ (.A(_15456_),
    .B(_15450_),
    .Y(_15632_));
 sky130_fd_sc_hd__a21oi_4 _46187_ (.A1(_15630_),
    .A2(_15631_),
    .B1(_15632_),
    .Y(_15633_));
 sky130_fd_sc_hd__nand3_4 _46188_ (.A(_15630_),
    .B(_15631_),
    .C(_15632_),
    .Y(_15634_));
 sky130_vsdinv _46189_ (.A(_15634_),
    .Y(_15635_));
 sky130_fd_sc_hd__nor2_4 _46190_ (.A(_15633_),
    .B(_15635_),
    .Y(_15636_));
 sky130_fd_sc_hd__nor2_4 _46191_ (.A(_15241_),
    .B(_15462_),
    .Y(_15637_));
 sky130_fd_sc_hd__nand2_4 _46192_ (.A(_15637_),
    .B(_15242_),
    .Y(_15638_));
 sky130_fd_sc_hd__nor2_4 _46193_ (.A(_14799_),
    .B(_15638_),
    .Y(_15639_));
 sky130_fd_sc_hd__nand4_4 _46194_ (.A(_14793_),
    .B(_14791_),
    .C(_15028_),
    .D(_15026_),
    .Y(_15640_));
 sky130_fd_sc_hd__nand4_4 _46195_ (.A(_15240_),
    .B(_15460_),
    .C(_15238_),
    .D(_15461_),
    .Y(_15641_));
 sky130_fd_sc_hd__nor2_4 _46196_ (.A(_15640_),
    .B(_15641_),
    .Y(_15642_));
 sky130_fd_sc_hd__nand2_4 _46197_ (.A(_14797_),
    .B(_15642_),
    .Y(_15643_));
 sky130_fd_sc_hd__a21boi_4 _46198_ (.A1(_15463_),
    .A2(_15460_),
    .B1_N(_15461_),
    .Y(_15644_));
 sky130_fd_sc_hd__o21a_4 _46199_ (.A1(_15245_),
    .A2(_15641_),
    .B1(_15644_),
    .X(_15645_));
 sky130_fd_sc_hd__nand2_4 _46200_ (.A(_15643_),
    .B(_15645_),
    .Y(_15646_));
 sky130_fd_sc_hd__a21oi_4 _46201_ (.A1(_13802_),
    .A2(_15639_),
    .B1(_15646_),
    .Y(_15647_));
 sky130_fd_sc_hd__nand4_4 _46202_ (.A(_14314_),
    .B(_15637_),
    .C(_14798_),
    .D(_15242_),
    .Y(_15648_));
 sky130_fd_sc_hd__nor2_4 _46203_ (.A(_13803_),
    .B(_15648_),
    .Y(_15649_));
 sky130_fd_sc_hd__nand2_4 _46204_ (.A(_11426_),
    .B(_15649_),
    .Y(_15650_));
 sky130_fd_sc_hd__nand2_4 _46205_ (.A(_15647_),
    .B(_15650_),
    .Y(_15651_));
 sky130_fd_sc_hd__buf_8 _46206_ (.A(_15651_),
    .X(_15652_));
 sky130_fd_sc_hd__xor2_4 _46207_ (.A(_15636_),
    .B(_15652_),
    .X(_01453_));
 sky130_fd_sc_hd__a21boi_4 _46208_ (.A1(_15543_),
    .A2(_15578_),
    .B1_N(_15545_),
    .Y(_15653_));
 sky130_vsdinv _46209_ (.A(_15653_),
    .Y(_15654_));
 sky130_fd_sc_hd__a21boi_4 _46210_ (.A1(_15488_),
    .A2(_15504_),
    .B1_N(_15487_),
    .Y(_15655_));
 sky130_vsdinv _46211_ (.A(_15655_),
    .Y(_15656_));
 sky130_fd_sc_hd__nand2_4 _46212_ (.A(_11871_),
    .B(_15033_),
    .Y(_15657_));
 sky130_fd_sc_hd__o21ai_4 _46213_ (.A1(_13042_),
    .A2(_03634_),
    .B1(_15657_),
    .Y(_15658_));
 sky130_fd_sc_hd__buf_4 _46214_ (.A(_10959_),
    .X(_15659_));
 sky130_fd_sc_hd__nand4_4 _46215_ (.A(_03333_),
    .B(_12189_),
    .C(_15659_),
    .D(_15253_),
    .Y(_15660_));
 sky130_fd_sc_hd__nand2_4 _46216_ (.A(_12192_),
    .B(_10517_),
    .Y(_15661_));
 sky130_vsdinv _46217_ (.A(_15661_),
    .Y(_15662_));
 sky130_fd_sc_hd__a21o_4 _46218_ (.A1(_15658_),
    .A2(_15660_),
    .B1(_15662_),
    .X(_15663_));
 sky130_fd_sc_hd__nand3_4 _46219_ (.A(_15658_),
    .B(_15660_),
    .C(_15662_),
    .Y(_15664_));
 sky130_fd_sc_hd__a21boi_4 _46220_ (.A1(_15467_),
    .A2(_15470_),
    .B1_N(_15468_),
    .Y(_15665_));
 sky130_fd_sc_hd__a21boi_4 _46221_ (.A1(_15663_),
    .A2(_15664_),
    .B1_N(_15665_),
    .Y(_15666_));
 sky130_vsdinv _46222_ (.A(_15666_),
    .Y(_15667_));
 sky130_vsdinv _46223_ (.A(_15665_),
    .Y(_15668_));
 sky130_fd_sc_hd__nand3_4 _46224_ (.A(_15668_),
    .B(_15663_),
    .C(_15664_),
    .Y(_15669_));
 sky130_fd_sc_hd__nand2_4 _46225_ (.A(_11242_),
    .B(_11777_),
    .Y(_15670_));
 sky130_fd_sc_hd__nand2_4 _46226_ (.A(_11030_),
    .B(_11776_),
    .Y(_15671_));
 sky130_fd_sc_hd__nand2_4 _46227_ (.A(_15670_),
    .B(_15671_),
    .Y(_15672_));
 sky130_fd_sc_hd__nand4_4 _46228_ (.A(_11033_),
    .B(_11034_),
    .C(_12406_),
    .D(_12404_),
    .Y(_15673_));
 sky130_fd_sc_hd__nand2_4 _46229_ (.A(_08755_),
    .B(_12095_),
    .Y(_15674_));
 sky130_vsdinv _46230_ (.A(_15674_),
    .Y(_15675_));
 sky130_fd_sc_hd__a21o_4 _46231_ (.A1(_15672_),
    .A2(_15673_),
    .B1(_15675_),
    .X(_15676_));
 sky130_fd_sc_hd__nand3_4 _46232_ (.A(_15672_),
    .B(_15673_),
    .C(_15675_),
    .Y(_15677_));
 sky130_fd_sc_hd__and2_4 _46233_ (.A(_15676_),
    .B(_15677_),
    .X(_15678_));
 sky130_fd_sc_hd__a21o_4 _46234_ (.A1(_15667_),
    .A2(_15669_),
    .B1(_15678_),
    .X(_15679_));
 sky130_fd_sc_hd__nand3_4 _46235_ (.A(_15667_),
    .B(_15669_),
    .C(_15678_),
    .Y(_15680_));
 sky130_fd_sc_hd__a21boi_4 _46236_ (.A1(_15475_),
    .A2(_15483_),
    .B1_N(_15474_),
    .Y(_15681_));
 sky130_fd_sc_hd__a21boi_4 _46237_ (.A1(_15679_),
    .A2(_15680_),
    .B1_N(_15681_),
    .Y(_15682_));
 sky130_vsdinv _46238_ (.A(_15682_),
    .Y(_15683_));
 sky130_vsdinv _46239_ (.A(_15681_),
    .Y(_15684_));
 sky130_fd_sc_hd__nand3_4 _46240_ (.A(_15684_),
    .B(_15679_),
    .C(_15680_),
    .Y(_15685_));
 sky130_fd_sc_hd__a21boi_4 _46241_ (.A1(_15498_),
    .A2(_15493_),
    .B1_N(_15500_),
    .Y(_15686_));
 sky130_vsdinv _46242_ (.A(_15476_),
    .Y(_15687_));
 sky130_fd_sc_hd__a21boi_4 _46243_ (.A1(_15480_),
    .A2(_15687_),
    .B1_N(_15481_),
    .Y(_15688_));
 sky130_fd_sc_hd__nand2_4 _46244_ (.A(_11249_),
    .B(_13298_),
    .Y(_15689_));
 sky130_fd_sc_hd__nand2_4 _46245_ (.A(_10666_),
    .B(_12111_),
    .Y(_15690_));
 sky130_fd_sc_hd__nand2_4 _46246_ (.A(_15689_),
    .B(_15690_),
    .Y(_15691_));
 sky130_fd_sc_hd__nand4_4 _46247_ (.A(_10783_),
    .B(_11287_),
    .C(_12114_),
    .D(_12115_),
    .Y(_15692_));
 sky130_fd_sc_hd__nand2_4 _46248_ (.A(_11635_),
    .B(_13303_),
    .Y(_15693_));
 sky130_vsdinv _46249_ (.A(_15693_),
    .Y(_15694_));
 sky130_fd_sc_hd__a21o_4 _46250_ (.A1(_15691_),
    .A2(_15692_),
    .B1(_15694_),
    .X(_15695_));
 sky130_fd_sc_hd__nand3_4 _46251_ (.A(_15691_),
    .B(_15692_),
    .C(_15694_),
    .Y(_15696_));
 sky130_fd_sc_hd__nand2_4 _46252_ (.A(_15695_),
    .B(_15696_),
    .Y(_15697_));
 sky130_fd_sc_hd__or2_4 _46253_ (.A(_15688_),
    .B(_15697_),
    .X(_15698_));
 sky130_fd_sc_hd__nand2_4 _46254_ (.A(_15697_),
    .B(_15688_),
    .Y(_15699_));
 sky130_fd_sc_hd__nand2_4 _46255_ (.A(_15698_),
    .B(_15699_),
    .Y(_15700_));
 sky130_fd_sc_hd__xor2_4 _46256_ (.A(_15686_),
    .B(_15700_),
    .X(_15701_));
 sky130_fd_sc_hd__a21o_4 _46257_ (.A1(_15683_),
    .A2(_15685_),
    .B1(_15701_),
    .X(_15702_));
 sky130_fd_sc_hd__nand3_4 _46258_ (.A(_15683_),
    .B(_15685_),
    .C(_15701_),
    .Y(_15703_));
 sky130_fd_sc_hd__nand3_4 _46259_ (.A(_15656_),
    .B(_15702_),
    .C(_15703_),
    .Y(_15704_));
 sky130_fd_sc_hd__nand2_4 _46260_ (.A(_15702_),
    .B(_15703_),
    .Y(_15705_));
 sky130_fd_sc_hd__nand2_4 _46261_ (.A(_15705_),
    .B(_15655_),
    .Y(_15706_));
 sky130_fd_sc_hd__maj3_4 _46262_ (.A(_15489_),
    .B(_15502_),
    .C(_15491_),
    .X(_15707_));
 sky130_fd_sc_hd__nand2_4 _46263_ (.A(_12277_),
    .B(_14872_),
    .Y(_15708_));
 sky130_fd_sc_hd__o21ai_4 _46264_ (.A1(_03380_),
    .A2(_03578_),
    .B1(_15708_),
    .Y(_15709_));
 sky130_fd_sc_hd__nand4_4 _46265_ (.A(_14884_),
    .B(_14882_),
    .C(_14872_),
    .D(_14873_),
    .Y(_15710_));
 sky130_fd_sc_hd__nand2_4 _46266_ (.A(_12279_),
    .B(_12754_),
    .Y(_15711_));
 sky130_vsdinv _46267_ (.A(_15711_),
    .Y(_15712_));
 sky130_fd_sc_hd__a21o_4 _46268_ (.A1(_15709_),
    .A2(_15710_),
    .B1(_15712_),
    .X(_15713_));
 sky130_fd_sc_hd__nand3_4 _46269_ (.A(_15709_),
    .B(_15710_),
    .C(_15712_),
    .Y(_15714_));
 sky130_fd_sc_hd__a21boi_4 _46270_ (.A1(_15514_),
    .A2(_15517_),
    .B1_N(_15515_),
    .Y(_15715_));
 sky130_vsdinv _46271_ (.A(_15715_),
    .Y(_15716_));
 sky130_fd_sc_hd__a21o_4 _46272_ (.A1(_15713_),
    .A2(_15714_),
    .B1(_15716_),
    .X(_15717_));
 sky130_fd_sc_hd__nand3_4 _46273_ (.A(_15716_),
    .B(_15713_),
    .C(_15714_),
    .Y(_15718_));
 sky130_fd_sc_hd__nand2_4 _46274_ (.A(_10838_),
    .B(_03546_),
    .Y(_15719_));
 sky130_fd_sc_hd__buf_1 _46275_ (.A(_10843_),
    .X(_15720_));
 sky130_fd_sc_hd__nand2_4 _46276_ (.A(_15720_),
    .B(_11523_),
    .Y(_15721_));
 sky130_fd_sc_hd__nand2_4 _46277_ (.A(_10847_),
    .B(_13611_),
    .Y(_15722_));
 sky130_fd_sc_hd__xnor2_4 _46278_ (.A(_15721_),
    .B(_15722_),
    .Y(_15723_));
 sky130_fd_sc_hd__xor2_4 _46279_ (.A(_15719_),
    .B(_15723_),
    .X(_15724_));
 sky130_fd_sc_hd__a21o_4 _46280_ (.A1(_15717_),
    .A2(_15718_),
    .B1(_15724_),
    .X(_15725_));
 sky130_fd_sc_hd__nand3_4 _46281_ (.A(_15724_),
    .B(_15717_),
    .C(_15718_),
    .Y(_15726_));
 sky130_fd_sc_hd__nand2_4 _46282_ (.A(_15725_),
    .B(_15726_),
    .Y(_15727_));
 sky130_fd_sc_hd__or2_4 _46283_ (.A(_15707_),
    .B(_15727_),
    .X(_15728_));
 sky130_fd_sc_hd__a21boi_4 _46284_ (.A1(_15725_),
    .A2(_15726_),
    .B1_N(_15707_),
    .Y(_15729_));
 sky130_vsdinv _46285_ (.A(_15729_),
    .Y(_15730_));
 sky130_fd_sc_hd__a21oi_4 _46286_ (.A1(_15528_),
    .A2(_15523_),
    .B1(_15521_),
    .Y(_15731_));
 sky130_vsdinv _46287_ (.A(_15731_),
    .Y(_15732_));
 sky130_fd_sc_hd__a21o_4 _46288_ (.A1(_15728_),
    .A2(_15730_),
    .B1(_15732_),
    .X(_15733_));
 sky130_fd_sc_hd__nand3_4 _46289_ (.A(_15728_),
    .B(_15730_),
    .C(_15732_),
    .Y(_15734_));
 sky130_fd_sc_hd__nand2_4 _46290_ (.A(_15733_),
    .B(_15734_),
    .Y(_15735_));
 sky130_vsdinv _46291_ (.A(_15735_),
    .Y(_15736_));
 sky130_fd_sc_hd__a21o_4 _46292_ (.A1(_15704_),
    .A2(_15706_),
    .B1(_15736_),
    .X(_15737_));
 sky130_fd_sc_hd__nand3_4 _46293_ (.A(_15704_),
    .B(_15706_),
    .C(_15736_),
    .Y(_15738_));
 sky130_fd_sc_hd__nand2_4 _46294_ (.A(_15737_),
    .B(_15738_),
    .Y(_15739_));
 sky130_fd_sc_hd__maj3_4 _46295_ (.A(_15507_),
    .B(_15538_),
    .C(_15508_),
    .X(_15740_));
 sky130_fd_sc_hd__nand2_4 _46296_ (.A(_15739_),
    .B(_15740_),
    .Y(_15741_));
 sky130_fd_sc_hd__nand2_4 _46297_ (.A(_15540_),
    .B(_15511_),
    .Y(_15742_));
 sky130_fd_sc_hd__nand3_4 _46298_ (.A(_15742_),
    .B(_15737_),
    .C(_15738_),
    .Y(_15743_));
 sky130_fd_sc_hd__nand2_4 _46299_ (.A(_11339_),
    .B(_07709_),
    .Y(_15744_));
 sky130_fd_sc_hd__nand2_4 _46300_ (.A(_15549_),
    .B(_15744_),
    .Y(_15745_));
 sky130_fd_sc_hd__nand3_4 _46301_ (.A(_11691_),
    .B(_08568_),
    .C(_07556_),
    .Y(_15746_));
 sky130_fd_sc_hd__nand3_4 _46302_ (.A(_15745_),
    .B(_15359_),
    .C(_15746_),
    .Y(_15747_));
 sky130_fd_sc_hd__a21o_4 _46303_ (.A1(_15745_),
    .A2(_15746_),
    .B1(_15359_),
    .X(_15748_));
 sky130_fd_sc_hd__maj3_4 _46304_ (.A(_15525_),
    .B(_15526_),
    .C(_15524_),
    .X(_15749_));
 sky130_vsdinv _46305_ (.A(_15749_),
    .Y(_15750_));
 sky130_fd_sc_hd__a21o_4 _46306_ (.A1(_15747_),
    .A2(_15748_),
    .B1(_15750_),
    .X(_15751_));
 sky130_fd_sc_hd__nand3_4 _46307_ (.A(_15750_),
    .B(_15747_),
    .C(_15748_),
    .Y(_15752_));
 sky130_fd_sc_hd__a21boi_4 _46308_ (.A1(_15550_),
    .A2(_15553_),
    .B1_N(_15551_),
    .Y(_15753_));
 sky130_vsdinv _46309_ (.A(_15753_),
    .Y(_15754_));
 sky130_fd_sc_hd__a21o_4 _46310_ (.A1(_15751_),
    .A2(_15752_),
    .B1(_15754_),
    .X(_15755_));
 sky130_fd_sc_hd__nand3_4 _46311_ (.A(_15751_),
    .B(_15752_),
    .C(_15754_),
    .Y(_15756_));
 sky130_fd_sc_hd__maj3_4 _46312_ (.A(_15547_),
    .B(_15555_),
    .C(_15558_),
    .X(_15757_));
 sky130_vsdinv _46313_ (.A(_15757_),
    .Y(_15758_));
 sky130_fd_sc_hd__a21o_4 _46314_ (.A1(_15755_),
    .A2(_15756_),
    .B1(_15758_),
    .X(_15759_));
 sky130_fd_sc_hd__nand3_4 _46315_ (.A(_15755_),
    .B(_15758_),
    .C(_15756_),
    .Y(_15760_));
 sky130_fd_sc_hd__a21o_4 _46316_ (.A1(_15759_),
    .A2(_15760_),
    .B1(_15379_),
    .X(_15761_));
 sky130_fd_sc_hd__buf_1 _46317_ (.A(_15383_),
    .X(_15762_));
 sky130_fd_sc_hd__nand3_4 _46318_ (.A(_15759_),
    .B(_15762_),
    .C(_15760_),
    .Y(_15763_));
 sky130_fd_sc_hd__nand2_4 _46319_ (.A(_15761_),
    .B(_15763_),
    .Y(_15764_));
 sky130_fd_sc_hd__a21o_4 _46320_ (.A1(_15532_),
    .A2(_15537_),
    .B1(_15764_),
    .X(_15765_));
 sky130_fd_sc_hd__nand3_4 _46321_ (.A(_15764_),
    .B(_15532_),
    .C(_15537_),
    .Y(_15766_));
 sky130_fd_sc_hd__buf_1 _46322_ (.A(_15379_),
    .X(_15767_));
 sky130_fd_sc_hd__a21boi_4 _46323_ (.A1(_15564_),
    .A2(_15767_),
    .B1_N(_15565_),
    .Y(_15768_));
 sky130_vsdinv _46324_ (.A(_15768_),
    .Y(_15769_));
 sky130_fd_sc_hd__a21o_4 _46325_ (.A1(_15765_),
    .A2(_15766_),
    .B1(_15769_),
    .X(_15770_));
 sky130_fd_sc_hd__nand3_4 _46326_ (.A(_15765_),
    .B(_15769_),
    .C(_15766_),
    .Y(_15771_));
 sky130_fd_sc_hd__and2_4 _46327_ (.A(_15770_),
    .B(_15771_),
    .X(_15772_));
 sky130_fd_sc_hd__nand3_4 _46328_ (.A(_15741_),
    .B(_15743_),
    .C(_15772_),
    .Y(_15773_));
 sky130_fd_sc_hd__nand2_4 _46329_ (.A(_15741_),
    .B(_15743_),
    .Y(_15774_));
 sky130_vsdinv _46330_ (.A(_15772_),
    .Y(_15775_));
 sky130_fd_sc_hd__nand2_4 _46331_ (.A(_15774_),
    .B(_15775_),
    .Y(_15776_));
 sky130_fd_sc_hd__nand3_4 _46332_ (.A(_15654_),
    .B(_15773_),
    .C(_15776_),
    .Y(_15777_));
 sky130_fd_sc_hd__nand2_4 _46333_ (.A(_15776_),
    .B(_15773_),
    .Y(_15778_));
 sky130_fd_sc_hd__nand2_4 _46334_ (.A(_15778_),
    .B(_15653_),
    .Y(_15779_));
 sky130_fd_sc_hd__nand2_4 _46335_ (.A(_15777_),
    .B(_15779_),
    .Y(_15780_));
 sky130_fd_sc_hd__nand4_4 _46336_ (.A(_13719_),
    .B(_15588_),
    .C(_14499_),
    .D(_14727_),
    .Y(_15781_));
 sky130_fd_sc_hd__nand2_4 _46337_ (.A(_15597_),
    .B(_15781_),
    .Y(_15782_));
 sky130_fd_sc_hd__nand4_4 _46338_ (.A(_13994_),
    .B(_15586_),
    .C(_13996_),
    .D(_14726_),
    .Y(_15783_));
 sky130_fd_sc_hd__nand2_4 _46339_ (.A(_15781_),
    .B(_15783_),
    .Y(_15784_));
 sky130_fd_sc_hd__xnor2_4 _46340_ (.A(_15784_),
    .B(_13478_),
    .Y(_15785_));
 sky130_vsdinv _46341_ (.A(_15785_),
    .Y(_15786_));
 sky130_fd_sc_hd__buf_1 _46342_ (.A(_15786_),
    .X(_15787_));
 sky130_fd_sc_hd__a21o_4 _46343_ (.A1(_15575_),
    .A2(_15569_),
    .B1(_15787_),
    .X(_15788_));
 sky130_fd_sc_hd__nand3_4 _46344_ (.A(_15575_),
    .B(_15569_),
    .C(_15787_),
    .Y(_15789_));
 sky130_fd_sc_hd__nand2_4 _46345_ (.A(_15788_),
    .B(_15789_),
    .Y(_15790_));
 sky130_fd_sc_hd__xor2_4 _46346_ (.A(_15782_),
    .B(_15790_),
    .X(_15791_));
 sky130_fd_sc_hd__nand2_4 _46347_ (.A(_15780_),
    .B(_15791_),
    .Y(_15792_));
 sky130_vsdinv _46348_ (.A(_15791_),
    .Y(_15793_));
 sky130_fd_sc_hd__nand3_4 _46349_ (.A(_15793_),
    .B(_15777_),
    .C(_15779_),
    .Y(_15794_));
 sky130_fd_sc_hd__nand2_4 _46350_ (.A(_15792_),
    .B(_15794_),
    .Y(_15795_));
 sky130_fd_sc_hd__nand2_4 _46351_ (.A(_15609_),
    .B(_15584_),
    .Y(_15796_));
 sky130_vsdinv _46352_ (.A(_15796_),
    .Y(_15797_));
 sky130_fd_sc_hd__nand2_4 _46353_ (.A(_15795_),
    .B(_15797_),
    .Y(_15798_));
 sky130_fd_sc_hd__nand3_4 _46354_ (.A(_15796_),
    .B(_15792_),
    .C(_15794_),
    .Y(_15799_));
 sky130_fd_sc_hd__nand2_4 _46355_ (.A(_15798_),
    .B(_15799_),
    .Y(_15800_));
 sky130_fd_sc_hd__buf_1 _46356_ (.A(_15440_),
    .X(_15801_));
 sky130_fd_sc_hd__a21boi_4 _46357_ (.A1(_15600_),
    .A2(_15603_),
    .B1_N(_15601_),
    .Y(_15802_));
 sky130_fd_sc_hd__xor2_4 _46358_ (.A(_15801_),
    .B(_15802_),
    .X(_15803_));
 sky130_fd_sc_hd__nand2_4 _46359_ (.A(_15800_),
    .B(_15803_),
    .Y(_15804_));
 sky130_vsdinv _46360_ (.A(_15803_),
    .Y(_15805_));
 sky130_fd_sc_hd__nand3_4 _46361_ (.A(_15798_),
    .B(_15799_),
    .C(_15805_),
    .Y(_15806_));
 sky130_fd_sc_hd__nand2_4 _46362_ (.A(_15804_),
    .B(_15806_),
    .Y(_15807_));
 sky130_fd_sc_hd__a21boi_4 _46363_ (.A1(_15612_),
    .A2(_15619_),
    .B1_N(_15614_),
    .Y(_15808_));
 sky130_fd_sc_hd__nand2_4 _46364_ (.A(_15807_),
    .B(_15808_),
    .Y(_15809_));
 sky130_vsdinv _46365_ (.A(_15808_),
    .Y(_15810_));
 sky130_fd_sc_hd__nand3_4 _46366_ (.A(_15810_),
    .B(_15806_),
    .C(_15804_),
    .Y(_15811_));
 sky130_fd_sc_hd__nand2_4 _46367_ (.A(_15809_),
    .B(_15811_),
    .Y(_15812_));
 sky130_fd_sc_hd__a21oi_4 _46368_ (.A1(_15428_),
    .A2(_15423_),
    .B1(_15627_),
    .Y(_15813_));
 sky130_vsdinv _46369_ (.A(_15813_),
    .Y(_15814_));
 sky130_fd_sc_hd__nand2_4 _46370_ (.A(_15812_),
    .B(_15814_),
    .Y(_15815_));
 sky130_fd_sc_hd__nand3_4 _46371_ (.A(_15809_),
    .B(_15811_),
    .C(_15813_),
    .Y(_15816_));
 sky130_fd_sc_hd__a21oi_4 _46372_ (.A1(_15618_),
    .A2(_15620_),
    .B1(_15624_),
    .Y(_15817_));
 sky130_fd_sc_hd__o21ai_4 _46373_ (.A1(_15629_),
    .A2(_15817_),
    .B1(_15625_),
    .Y(_15818_));
 sky130_fd_sc_hd__a21oi_4 _46374_ (.A1(_15815_),
    .A2(_15816_),
    .B1(_15818_),
    .Y(_15819_));
 sky130_fd_sc_hd__nand3_4 _46375_ (.A(_15815_),
    .B(_15818_),
    .C(_15816_),
    .Y(_15820_));
 sky130_vsdinv _46376_ (.A(_15820_),
    .Y(_15821_));
 sky130_fd_sc_hd__nor2_4 _46377_ (.A(_15819_),
    .B(_15821_),
    .Y(_15822_));
 sky130_fd_sc_hd__a21oi_4 _46378_ (.A1(_15652_),
    .A2(_15636_),
    .B1(_15635_),
    .Y(_15823_));
 sky130_fd_sc_hd__xnor2_4 _46379_ (.A(_15822_),
    .B(_15823_),
    .Y(_01454_));
 sky130_fd_sc_hd__a21boi_4 _46380_ (.A1(_15706_),
    .A2(_15736_),
    .B1_N(_15704_),
    .Y(_15824_));
 sky130_vsdinv _46381_ (.A(_15824_),
    .Y(_15825_));
 sky130_fd_sc_hd__nand2_4 _46382_ (.A(_08307_),
    .B(_15465_),
    .Y(_15826_));
 sky130_fd_sc_hd__o21ai_4 _46383_ (.A1(_12189_),
    .A2(_03634_),
    .B1(_15826_),
    .Y(_15827_));
 sky130_fd_sc_hd__nand4_4 _46384_ (.A(_03338_),
    .B(_10624_),
    .C(_15465_),
    .D(_11384_),
    .Y(_15828_));
 sky130_fd_sc_hd__nand2_4 _46385_ (.A(_08309_),
    .B(_10517_),
    .Y(_15829_));
 sky130_vsdinv _46386_ (.A(_15829_),
    .Y(_15830_));
 sky130_fd_sc_hd__a21o_4 _46387_ (.A1(_15827_),
    .A2(_15828_),
    .B1(_15830_),
    .X(_15831_));
 sky130_fd_sc_hd__nand3_4 _46388_ (.A(_15827_),
    .B(_15828_),
    .C(_15830_),
    .Y(_15832_));
 sky130_fd_sc_hd__a21boi_4 _46389_ (.A1(_15658_),
    .A2(_15662_),
    .B1_N(_15660_),
    .Y(_15833_));
 sky130_fd_sc_hd__a21boi_4 _46390_ (.A1(_15831_),
    .A2(_15832_),
    .B1_N(_15833_),
    .Y(_15834_));
 sky130_vsdinv _46391_ (.A(_15834_),
    .Y(_15835_));
 sky130_vsdinv _46392_ (.A(_15833_),
    .Y(_15836_));
 sky130_fd_sc_hd__nand3_4 _46393_ (.A(_15836_),
    .B(_15831_),
    .C(_15832_),
    .Y(_15837_));
 sky130_fd_sc_hd__nand2_4 _46394_ (.A(_08528_),
    .B(_12410_),
    .Y(_15838_));
 sky130_fd_sc_hd__nand2_4 _46395_ (.A(_11593_),
    .B(_12409_),
    .Y(_15839_));
 sky130_fd_sc_hd__nand2_4 _46396_ (.A(_15838_),
    .B(_15839_),
    .Y(_15840_));
 sky130_fd_sc_hd__nand4_4 _46397_ (.A(_13087_),
    .B(_13084_),
    .C(_15478_),
    .D(_03614_),
    .Y(_15841_));
 sky130_fd_sc_hd__nand2_4 _46398_ (.A(_10788_),
    .B(_03601_),
    .Y(_15842_));
 sky130_vsdinv _46399_ (.A(_15842_),
    .Y(_15843_));
 sky130_fd_sc_hd__a21o_4 _46400_ (.A1(_15840_),
    .A2(_15841_),
    .B1(_15843_),
    .X(_15844_));
 sky130_fd_sc_hd__nand3_4 _46401_ (.A(_15840_),
    .B(_15841_),
    .C(_15843_),
    .Y(_15845_));
 sky130_fd_sc_hd__and2_4 _46402_ (.A(_15844_),
    .B(_15845_),
    .X(_15846_));
 sky130_fd_sc_hd__buf_1 _46403_ (.A(_15846_),
    .X(_15847_));
 sky130_fd_sc_hd__a21o_4 _46404_ (.A1(_15835_),
    .A2(_15837_),
    .B1(_15847_),
    .X(_15848_));
 sky130_fd_sc_hd__nand3_4 _46405_ (.A(_15835_),
    .B(_15837_),
    .C(_15847_),
    .Y(_15849_));
 sky130_vsdinv _46406_ (.A(_15678_),
    .Y(_15850_));
 sky130_fd_sc_hd__o21a_4 _46407_ (.A1(_15666_),
    .A2(_15850_),
    .B1(_15669_),
    .X(_15851_));
 sky130_vsdinv _46408_ (.A(_15851_),
    .Y(_15852_));
 sky130_fd_sc_hd__a21oi_4 _46409_ (.A1(_15848_),
    .A2(_15849_),
    .B1(_15852_),
    .Y(_15853_));
 sky130_vsdinv _46410_ (.A(_15853_),
    .Y(_15854_));
 sky130_fd_sc_hd__nand3_4 _46411_ (.A(_15852_),
    .B(_15848_),
    .C(_15849_),
    .Y(_15855_));
 sky130_fd_sc_hd__a21boi_4 _46412_ (.A1(_15691_),
    .A2(_15694_),
    .B1_N(_15692_),
    .Y(_15856_));
 sky130_fd_sc_hd__a21boi_4 _46413_ (.A1(_15672_),
    .A2(_15675_),
    .B1_N(_15673_),
    .Y(_15857_));
 sky130_fd_sc_hd__buf_1 _46414_ (.A(_12719_),
    .X(_15858_));
 sky130_fd_sc_hd__nand2_4 _46415_ (.A(_12533_),
    .B(_15858_),
    .Y(_15859_));
 sky130_fd_sc_hd__buf_1 _46416_ (.A(_12114_),
    .X(_15860_));
 sky130_fd_sc_hd__nand2_4 _46417_ (.A(_12233_),
    .B(_15860_),
    .Y(_15861_));
 sky130_fd_sc_hd__nand2_4 _46418_ (.A(_15859_),
    .B(_15861_),
    .Y(_15862_));
 sky130_fd_sc_hd__buf_1 _46419_ (.A(_10789_),
    .X(_15863_));
 sky130_fd_sc_hd__buf_1 _46420_ (.A(_11893_),
    .X(_15864_));
 sky130_fd_sc_hd__buf_1 _46421_ (.A(_15494_),
    .X(_15865_));
 sky130_fd_sc_hd__nand4_4 _46422_ (.A(_15863_),
    .B(_15864_),
    .C(_03589_),
    .D(_15865_),
    .Y(_15866_));
 sky130_fd_sc_hd__nand2_4 _46423_ (.A(_13117_),
    .B(_03583_),
    .Y(_15867_));
 sky130_vsdinv _46424_ (.A(_15867_),
    .Y(_15868_));
 sky130_fd_sc_hd__a21o_4 _46425_ (.A1(_15862_),
    .A2(_15866_),
    .B1(_15868_),
    .X(_15869_));
 sky130_fd_sc_hd__nand3_4 _46426_ (.A(_15862_),
    .B(_15866_),
    .C(_15868_),
    .Y(_15870_));
 sky130_fd_sc_hd__nand2_4 _46427_ (.A(_15869_),
    .B(_15870_),
    .Y(_15871_));
 sky130_fd_sc_hd__xnor2_4 _46428_ (.A(_15857_),
    .B(_15871_),
    .Y(_15872_));
 sky130_fd_sc_hd__xor2_4 _46429_ (.A(_15856_),
    .B(_15872_),
    .X(_15873_));
 sky130_fd_sc_hd__a21o_4 _46430_ (.A1(_15854_),
    .A2(_15855_),
    .B1(_15873_),
    .X(_15874_));
 sky130_fd_sc_hd__nand3_4 _46431_ (.A(_15854_),
    .B(_15855_),
    .C(_15873_),
    .Y(_15875_));
 sky130_vsdinv _46432_ (.A(_15701_),
    .Y(_15876_));
 sky130_fd_sc_hd__o21a_4 _46433_ (.A1(_15682_),
    .A2(_15876_),
    .B1(_15685_),
    .X(_15877_));
 sky130_fd_sc_hd__a21boi_4 _46434_ (.A1(_15874_),
    .A2(_15875_),
    .B1_N(_15877_),
    .Y(_15878_));
 sky130_vsdinv _46435_ (.A(_15877_),
    .Y(_15879_));
 sky130_fd_sc_hd__nand3_4 _46436_ (.A(_15879_),
    .B(_15874_),
    .C(_15875_),
    .Y(_15880_));
 sky130_vsdinv _46437_ (.A(_15880_),
    .Y(_15881_));
 sky130_fd_sc_hd__maj3_4 _46438_ (.A(_15686_),
    .B(_15697_),
    .C(_15688_),
    .X(_15882_));
 sky130_fd_sc_hd__nand2_4 _46439_ (.A(_11957_),
    .B(_11172_),
    .Y(_15883_));
 sky130_fd_sc_hd__o21ai_4 _46440_ (.A1(_03384_),
    .A2(_03578_),
    .B1(_15883_),
    .Y(_15884_));
 sky130_fd_sc_hd__buf_1 _46441_ (.A(_12278_),
    .X(_15885_));
 sky130_fd_sc_hd__nand4_4 _46442_ (.A(_11955_),
    .B(_15885_),
    .C(_14869_),
    .D(_14867_),
    .Y(_15886_));
 sky130_fd_sc_hd__nand2_4 _46443_ (.A(_15132_),
    .B(_13872_),
    .Y(_15887_));
 sky130_vsdinv _46444_ (.A(_15887_),
    .Y(_15888_));
 sky130_fd_sc_hd__a21o_4 _46445_ (.A1(_15884_),
    .A2(_15886_),
    .B1(_15888_),
    .X(_15889_));
 sky130_fd_sc_hd__nand3_4 _46446_ (.A(_15884_),
    .B(_15886_),
    .C(_15888_),
    .Y(_15890_));
 sky130_fd_sc_hd__a21boi_4 _46447_ (.A1(_15709_),
    .A2(_15712_),
    .B1_N(_15710_),
    .Y(_15891_));
 sky130_vsdinv _46448_ (.A(_15891_),
    .Y(_15892_));
 sky130_fd_sc_hd__a21o_4 _46449_ (.A1(_15889_),
    .A2(_15890_),
    .B1(_15892_),
    .X(_15893_));
 sky130_fd_sc_hd__nand3_4 _46450_ (.A(_15892_),
    .B(_15889_),
    .C(_15890_),
    .Y(_15894_));
 sky130_fd_sc_hd__nand2_4 _46451_ (.A(_11692_),
    .B(_12456_),
    .Y(_15895_));
 sky130_fd_sc_hd__buf_1 _46452_ (.A(_15895_),
    .X(_15896_));
 sky130_fd_sc_hd__buf_1 _46453_ (.A(_13169_),
    .X(_15897_));
 sky130_fd_sc_hd__nand2_4 _46454_ (.A(_15897_),
    .B(_13885_),
    .Y(_15898_));
 sky130_fd_sc_hd__buf_1 _46455_ (.A(_12313_),
    .X(_15899_));
 sky130_fd_sc_hd__nand2_4 _46456_ (.A(_15899_),
    .B(_13884_),
    .Y(_15900_));
 sky130_fd_sc_hd__xnor2_4 _46457_ (.A(_15898_),
    .B(_15900_),
    .Y(_15901_));
 sky130_fd_sc_hd__xor2_4 _46458_ (.A(_15896_),
    .B(_15901_),
    .X(_15902_));
 sky130_fd_sc_hd__a21o_4 _46459_ (.A1(_15893_),
    .A2(_15894_),
    .B1(_15902_),
    .X(_15903_));
 sky130_fd_sc_hd__nand3_4 _46460_ (.A(_15902_),
    .B(_15893_),
    .C(_15894_),
    .Y(_15904_));
 sky130_fd_sc_hd__nand2_4 _46461_ (.A(_15903_),
    .B(_15904_),
    .Y(_15905_));
 sky130_fd_sc_hd__or2_4 _46462_ (.A(_15882_),
    .B(_15905_),
    .X(_15906_));
 sky130_fd_sc_hd__nand2_4 _46463_ (.A(_15905_),
    .B(_15882_),
    .Y(_15907_));
 sky130_fd_sc_hd__a21boi_4 _46464_ (.A1(_15724_),
    .A2(_15717_),
    .B1_N(_15718_),
    .Y(_15908_));
 sky130_vsdinv _46465_ (.A(_15908_),
    .Y(_15909_));
 sky130_fd_sc_hd__a21o_4 _46466_ (.A1(_15906_),
    .A2(_15907_),
    .B1(_15909_),
    .X(_15910_));
 sky130_fd_sc_hd__nand3_4 _46467_ (.A(_15906_),
    .B(_15909_),
    .C(_15907_),
    .Y(_15911_));
 sky130_fd_sc_hd__nand2_4 _46468_ (.A(_15910_),
    .B(_15911_),
    .Y(_15912_));
 sky130_fd_sc_hd__o21ai_4 _46469_ (.A1(_15878_),
    .A2(_15881_),
    .B1(_15912_),
    .Y(_15913_));
 sky130_vsdinv _46470_ (.A(_15878_),
    .Y(_15914_));
 sky130_fd_sc_hd__nand4_4 _46471_ (.A(_15914_),
    .B(_15880_),
    .C(_15911_),
    .D(_15910_),
    .Y(_15915_));
 sky130_fd_sc_hd__nand3_4 _46472_ (.A(_15825_),
    .B(_15913_),
    .C(_15915_),
    .Y(_15916_));
 sky130_fd_sc_hd__nand2_4 _46473_ (.A(_15913_),
    .B(_15915_),
    .Y(_15917_));
 sky130_fd_sc_hd__nand2_4 _46474_ (.A(_15917_),
    .B(_15824_),
    .Y(_15918_));
 sky130_fd_sc_hd__nand2_4 _46475_ (.A(_15916_),
    .B(_15918_),
    .Y(_15919_));
 sky130_fd_sc_hd__maj3_4 _46476_ (.A(_15721_),
    .B(_15722_),
    .C(_15719_),
    .X(_15920_));
 sky130_fd_sc_hd__and2_4 _46477_ (.A(_15748_),
    .B(_15747_),
    .X(_15921_));
 sky130_fd_sc_hd__buf_1 _46478_ (.A(_15921_),
    .X(_15922_));
 sky130_vsdinv _46479_ (.A(_15922_),
    .Y(_15923_));
 sky130_fd_sc_hd__or2_4 _46480_ (.A(_15920_),
    .B(_15923_),
    .X(_15924_));
 sky130_fd_sc_hd__buf_1 _46481_ (.A(_15747_),
    .X(_15925_));
 sky130_fd_sc_hd__a21bo_4 _46482_ (.A1(_15925_),
    .A2(_15748_),
    .B1_N(_15920_),
    .X(_15926_));
 sky130_fd_sc_hd__buf_1 _46483_ (.A(_15746_),
    .X(_15927_));
 sky130_fd_sc_hd__a21boi_4 _46484_ (.A1(_15745_),
    .A2(_15553_),
    .B1_N(_15927_),
    .Y(_15928_));
 sky130_vsdinv _46485_ (.A(_15928_),
    .Y(_15929_));
 sky130_fd_sc_hd__a21o_4 _46486_ (.A1(_15924_),
    .A2(_15926_),
    .B1(_15929_),
    .X(_15930_));
 sky130_fd_sc_hd__nand3_4 _46487_ (.A(_15924_),
    .B(_15926_),
    .C(_15929_),
    .Y(_15931_));
 sky130_fd_sc_hd__nand2_4 _46488_ (.A(_15930_),
    .B(_15931_),
    .Y(_15932_));
 sky130_fd_sc_hd__a21boi_4 _46489_ (.A1(_15751_),
    .A2(_15754_),
    .B1_N(_15752_),
    .Y(_15933_));
 sky130_fd_sc_hd__nand2_4 _46490_ (.A(_15932_),
    .B(_15933_),
    .Y(_15934_));
 sky130_vsdinv _46491_ (.A(_15933_),
    .Y(_15935_));
 sky130_fd_sc_hd__nand3_4 _46492_ (.A(_15930_),
    .B(_15931_),
    .C(_15935_),
    .Y(_15936_));
 sky130_fd_sc_hd__a21o_4 _46493_ (.A1(_15934_),
    .A2(_15936_),
    .B1(_15571_),
    .X(_15937_));
 sky130_fd_sc_hd__nand3_4 _46494_ (.A(_15934_),
    .B(_15767_),
    .C(_15936_),
    .Y(_15938_));
 sky130_fd_sc_hd__maj3_4 _46495_ (.A(_15731_),
    .B(_15727_),
    .C(_15707_),
    .X(_15939_));
 sky130_vsdinv _46496_ (.A(_15939_),
    .Y(_15940_));
 sky130_fd_sc_hd__a21o_4 _46497_ (.A1(_15937_),
    .A2(_15938_),
    .B1(_15940_),
    .X(_15941_));
 sky130_fd_sc_hd__nand3_4 _46498_ (.A(_15937_),
    .B(_15940_),
    .C(_15938_),
    .Y(_15942_));
 sky130_fd_sc_hd__buf_1 _46499_ (.A(_15762_),
    .X(_15943_));
 sky130_fd_sc_hd__a21boi_4 _46500_ (.A1(_15759_),
    .A2(_15943_),
    .B1_N(_15760_),
    .Y(_15944_));
 sky130_vsdinv _46501_ (.A(_15944_),
    .Y(_15945_));
 sky130_fd_sc_hd__a21oi_4 _46502_ (.A1(_15941_),
    .A2(_15942_),
    .B1(_15945_),
    .Y(_15946_));
 sky130_vsdinv _46503_ (.A(_15946_),
    .Y(_15947_));
 sky130_fd_sc_hd__nand3_4 _46504_ (.A(_15941_),
    .B(_15945_),
    .C(_15942_),
    .Y(_15948_));
 sky130_fd_sc_hd__nand2_4 _46505_ (.A(_15947_),
    .B(_15948_),
    .Y(_15949_));
 sky130_fd_sc_hd__nand2_4 _46506_ (.A(_15919_),
    .B(_15949_),
    .Y(_15950_));
 sky130_vsdinv _46507_ (.A(_15948_),
    .Y(_15951_));
 sky130_fd_sc_hd__nor2_4 _46508_ (.A(_15946_),
    .B(_15951_),
    .Y(_15952_));
 sky130_fd_sc_hd__nand3_4 _46509_ (.A(_15916_),
    .B(_15918_),
    .C(_15952_),
    .Y(_15953_));
 sky130_fd_sc_hd__nand2_4 _46510_ (.A(_15950_),
    .B(_15953_),
    .Y(_15954_));
 sky130_fd_sc_hd__a21boi_4 _46511_ (.A1(_15741_),
    .A2(_15772_),
    .B1_N(_15743_),
    .Y(_15955_));
 sky130_fd_sc_hd__nand2_4 _46512_ (.A(_15954_),
    .B(_15955_),
    .Y(_15956_));
 sky130_fd_sc_hd__nand2_4 _46513_ (.A(_15773_),
    .B(_15743_),
    .Y(_15957_));
 sky130_fd_sc_hd__nand3_4 _46514_ (.A(_15957_),
    .B(_15950_),
    .C(_15953_),
    .Y(_15958_));
 sky130_fd_sc_hd__nand2_4 _46515_ (.A(_15956_),
    .B(_15958_),
    .Y(_15959_));
 sky130_fd_sc_hd__a21o_4 _46516_ (.A1(_15771_),
    .A2(_15765_),
    .B1(_15787_),
    .X(_15960_));
 sky130_fd_sc_hd__buf_1 _46517_ (.A(_15786_),
    .X(_15961_));
 sky130_fd_sc_hd__buf_1 _46518_ (.A(_15961_),
    .X(_15962_));
 sky130_fd_sc_hd__nand3_4 _46519_ (.A(_15771_),
    .B(_15962_),
    .C(_15765_),
    .Y(_15963_));
 sky130_fd_sc_hd__a21boi_4 _46520_ (.A1(_14015_),
    .A2(_15783_),
    .B1_N(_15781_),
    .Y(_15964_));
 sky130_vsdinv _46521_ (.A(_15964_),
    .Y(_15965_));
 sky130_fd_sc_hd__buf_1 _46522_ (.A(_15965_),
    .X(_15966_));
 sky130_fd_sc_hd__a21o_4 _46523_ (.A1(_15960_),
    .A2(_15963_),
    .B1(_15966_),
    .X(_15967_));
 sky130_fd_sc_hd__nand3_4 _46524_ (.A(_15960_),
    .B(_15966_),
    .C(_15963_),
    .Y(_15968_));
 sky130_fd_sc_hd__and2_4 _46525_ (.A(_15967_),
    .B(_15968_),
    .X(_15969_));
 sky130_vsdinv _46526_ (.A(_15969_),
    .Y(_15970_));
 sky130_fd_sc_hd__nand2_4 _46527_ (.A(_15959_),
    .B(_15970_),
    .Y(_15971_));
 sky130_fd_sc_hd__nand3_4 _46528_ (.A(_15956_),
    .B(_15958_),
    .C(_15969_),
    .Y(_15972_));
 sky130_fd_sc_hd__nand2_4 _46529_ (.A(_15971_),
    .B(_15972_),
    .Y(_15973_));
 sky130_fd_sc_hd__a21boi_4 _46530_ (.A1(_15793_),
    .A2(_15779_),
    .B1_N(_15777_),
    .Y(_15974_));
 sky130_fd_sc_hd__nand2_4 _46531_ (.A(_15973_),
    .B(_15974_),
    .Y(_15975_));
 sky130_fd_sc_hd__a21boi_4 _46532_ (.A1(_15776_),
    .A2(_15773_),
    .B1_N(_15653_),
    .Y(_15976_));
 sky130_fd_sc_hd__o21ai_4 _46533_ (.A1(_15791_),
    .A2(_15976_),
    .B1(_15777_),
    .Y(_15977_));
 sky130_fd_sc_hd__nand3_4 _46534_ (.A(_15977_),
    .B(_15971_),
    .C(_15972_),
    .Y(_15978_));
 sky130_fd_sc_hd__nand2_4 _46535_ (.A(_15975_),
    .B(_15978_),
    .Y(_15979_));
 sky130_fd_sc_hd__a21bo_4 _46536_ (.A1(_15782_),
    .A2(_15789_),
    .B1_N(_15788_),
    .X(_15980_));
 sky130_fd_sc_hd__xor2_4 _46537_ (.A(_15801_),
    .B(_15980_),
    .X(_15981_));
 sky130_vsdinv _46538_ (.A(_15981_),
    .Y(_15982_));
 sky130_fd_sc_hd__nand2_4 _46539_ (.A(_15979_),
    .B(_15982_),
    .Y(_15983_));
 sky130_fd_sc_hd__nand3_4 _46540_ (.A(_15975_),
    .B(_15981_),
    .C(_15978_),
    .Y(_15984_));
 sky130_fd_sc_hd__nand2_4 _46541_ (.A(_15983_),
    .B(_15984_),
    .Y(_15985_));
 sky130_fd_sc_hd__a21boi_4 _46542_ (.A1(_15798_),
    .A2(_15805_),
    .B1_N(_15799_),
    .Y(_15986_));
 sky130_fd_sc_hd__nand2_4 _46543_ (.A(_15985_),
    .B(_15986_),
    .Y(_15987_));
 sky130_fd_sc_hd__nand2_4 _46544_ (.A(_15806_),
    .B(_15799_),
    .Y(_15988_));
 sky130_fd_sc_hd__nand3_4 _46545_ (.A(_15988_),
    .B(_15984_),
    .C(_15983_),
    .Y(_15989_));
 sky130_fd_sc_hd__nand2_4 _46546_ (.A(_15987_),
    .B(_15989_),
    .Y(_15990_));
 sky130_fd_sc_hd__a21oi_4 _46547_ (.A1(_15605_),
    .A2(_15601_),
    .B1(_15452_),
    .Y(_15991_));
 sky130_vsdinv _46548_ (.A(_15991_),
    .Y(_15992_));
 sky130_fd_sc_hd__nand2_4 _46549_ (.A(_15990_),
    .B(_15992_),
    .Y(_15993_));
 sky130_fd_sc_hd__nand3_4 _46550_ (.A(_15987_),
    .B(_15989_),
    .C(_15991_),
    .Y(_15994_));
 sky130_fd_sc_hd__nand2_4 _46551_ (.A(_15993_),
    .B(_15994_),
    .Y(_15995_));
 sky130_fd_sc_hd__a21boi_4 _46552_ (.A1(_15809_),
    .A2(_15813_),
    .B1_N(_15811_),
    .Y(_15996_));
 sky130_fd_sc_hd__nand2_4 _46553_ (.A(_15995_),
    .B(_15996_),
    .Y(_15997_));
 sky130_fd_sc_hd__nand2_4 _46554_ (.A(_15816_),
    .B(_15811_),
    .Y(_15998_));
 sky130_fd_sc_hd__nand3_4 _46555_ (.A(_15998_),
    .B(_15993_),
    .C(_15994_),
    .Y(_15999_));
 sky130_fd_sc_hd__and2_4 _46556_ (.A(_15997_),
    .B(_15999_),
    .X(_16000_));
 sky130_fd_sc_hd__buf_1 _46557_ (.A(_16000_),
    .X(_16001_));
 sky130_vsdinv _46558_ (.A(_16001_),
    .Y(_16002_));
 sky130_fd_sc_hd__nand2_4 _46559_ (.A(_15815_),
    .B(_15816_),
    .Y(_16003_));
 sky130_vsdinv _46560_ (.A(_15818_),
    .Y(_16004_));
 sky130_fd_sc_hd__nand2_4 _46561_ (.A(_16003_),
    .B(_16004_),
    .Y(_16005_));
 sky130_fd_sc_hd__nand2_4 _46562_ (.A(_15820_),
    .B(_15634_),
    .Y(_16006_));
 sky130_fd_sc_hd__a32oi_4 _46563_ (.A1(_15652_),
    .A2(_15636_),
    .A3(_15822_),
    .B1(_16005_),
    .B2(_16006_),
    .Y(_16007_));
 sky130_fd_sc_hd__xor2_4 _46564_ (.A(_16002_),
    .B(_16007_),
    .X(_01455_));
 sky130_fd_sc_hd__nand2_4 _46565_ (.A(_11904_),
    .B(_15033_),
    .Y(_16008_));
 sky130_fd_sc_hd__o21ai_4 _46566_ (.A1(_11022_),
    .A2(_03634_),
    .B1(_16008_),
    .Y(_16009_));
 sky130_fd_sc_hd__nand4_4 _46567_ (.A(_03343_),
    .B(_11243_),
    .C(_15659_),
    .D(_15253_),
    .Y(_16010_));
 sky130_fd_sc_hd__nand2_4 _46568_ (.A(_08754_),
    .B(_03621_),
    .Y(_16011_));
 sky130_vsdinv _46569_ (.A(_16011_),
    .Y(_16012_));
 sky130_fd_sc_hd__a21o_4 _46570_ (.A1(_16009_),
    .A2(_16010_),
    .B1(_16012_),
    .X(_16013_));
 sky130_fd_sc_hd__nand3_4 _46571_ (.A(_16009_),
    .B(_16010_),
    .C(_16012_),
    .Y(_16014_));
 sky130_fd_sc_hd__a21boi_4 _46572_ (.A1(_15827_),
    .A2(_15830_),
    .B1_N(_15828_),
    .Y(_16015_));
 sky130_vsdinv _46573_ (.A(_16015_),
    .Y(_16016_));
 sky130_fd_sc_hd__a21o_4 _46574_ (.A1(_16013_),
    .A2(_16014_),
    .B1(_16016_),
    .X(_16017_));
 sky130_fd_sc_hd__nand3_4 _46575_ (.A(_16016_),
    .B(_16013_),
    .C(_16014_),
    .Y(_16018_));
 sky130_fd_sc_hd__nand2_4 _46576_ (.A(_12530_),
    .B(_10509_),
    .Y(_16019_));
 sky130_fd_sc_hd__nand2_4 _46577_ (.A(_11912_),
    .B(_03614_),
    .Y(_16020_));
 sky130_fd_sc_hd__nand2_4 _46578_ (.A(_15496_),
    .B(_15478_),
    .Y(_16021_));
 sky130_fd_sc_hd__nand2_4 _46579_ (.A(_16020_),
    .B(_16021_),
    .Y(_16022_));
 sky130_fd_sc_hd__nand4_4 _46580_ (.A(_08756_),
    .B(_15496_),
    .C(_15478_),
    .D(_03614_),
    .Y(_16023_));
 sky130_fd_sc_hd__nand2_4 _46581_ (.A(_16022_),
    .B(_16023_),
    .Y(_16024_));
 sky130_fd_sc_hd__xor2_4 _46582_ (.A(_16019_),
    .B(_16024_),
    .X(_16025_));
 sky130_fd_sc_hd__a21o_4 _46583_ (.A1(_16017_),
    .A2(_16018_),
    .B1(_16025_),
    .X(_16026_));
 sky130_fd_sc_hd__nand3_4 _46584_ (.A(_16017_),
    .B(_16018_),
    .C(_16025_),
    .Y(_16027_));
 sky130_fd_sc_hd__a21boi_4 _46585_ (.A1(_15835_),
    .A2(_15847_),
    .B1_N(_15837_),
    .Y(_16028_));
 sky130_vsdinv _46586_ (.A(_16028_),
    .Y(_16029_));
 sky130_fd_sc_hd__a21o_4 _46587_ (.A1(_16026_),
    .A2(_16027_),
    .B1(_16029_),
    .X(_16030_));
 sky130_fd_sc_hd__nand3_4 _46588_ (.A(_16029_),
    .B(_16026_),
    .C(_16027_),
    .Y(_16031_));
 sky130_fd_sc_hd__a21boi_4 _46589_ (.A1(_15862_),
    .A2(_15868_),
    .B1_N(_15866_),
    .Y(_16032_));
 sky130_fd_sc_hd__a21boi_4 _46590_ (.A1(_15840_),
    .A2(_15843_),
    .B1_N(_15841_),
    .Y(_16033_));
 sky130_fd_sc_hd__nand2_4 _46591_ (.A(_12824_),
    .B(_15865_),
    .Y(_16034_));
 sky130_fd_sc_hd__nand2_4 _46592_ (.A(_13117_),
    .B(_15860_),
    .Y(_16035_));
 sky130_fd_sc_hd__nand2_4 _46593_ (.A(_16034_),
    .B(_16035_),
    .Y(_16036_));
 sky130_fd_sc_hd__buf_1 _46594_ (.A(_12821_),
    .X(_16037_));
 sky130_fd_sc_hd__buf_1 _46595_ (.A(_11949_),
    .X(_16038_));
 sky130_fd_sc_hd__nand4_4 _46596_ (.A(_16037_),
    .B(_16038_),
    .C(_15860_),
    .D(_15865_),
    .Y(_16039_));
 sky130_fd_sc_hd__buf_1 _46597_ (.A(_12273_),
    .X(_16040_));
 sky130_fd_sc_hd__nand2_4 _46598_ (.A(_16040_),
    .B(_03583_),
    .Y(_16041_));
 sky130_vsdinv _46599_ (.A(_16041_),
    .Y(_16042_));
 sky130_fd_sc_hd__a21o_4 _46600_ (.A1(_16036_),
    .A2(_16039_),
    .B1(_16042_),
    .X(_16043_));
 sky130_fd_sc_hd__nand3_4 _46601_ (.A(_16036_),
    .B(_16039_),
    .C(_16042_),
    .Y(_16044_));
 sky130_fd_sc_hd__nand2_4 _46602_ (.A(_16043_),
    .B(_16044_),
    .Y(_16045_));
 sky130_fd_sc_hd__xnor2_4 _46603_ (.A(_16033_),
    .B(_16045_),
    .Y(_16046_));
 sky130_fd_sc_hd__xor2_4 _46604_ (.A(_16032_),
    .B(_16046_),
    .X(_16047_));
 sky130_fd_sc_hd__a21o_4 _46605_ (.A1(_16030_),
    .A2(_16031_),
    .B1(_16047_),
    .X(_16048_));
 sky130_fd_sc_hd__nand3_4 _46606_ (.A(_16030_),
    .B(_16031_),
    .C(_16047_),
    .Y(_16049_));
 sky130_fd_sc_hd__a21boi_4 _46607_ (.A1(_15854_),
    .A2(_15873_),
    .B1_N(_15855_),
    .Y(_16050_));
 sky130_vsdinv _46608_ (.A(_16050_),
    .Y(_16051_));
 sky130_fd_sc_hd__a21o_4 _46609_ (.A1(_16048_),
    .A2(_16049_),
    .B1(_16051_),
    .X(_16052_));
 sky130_fd_sc_hd__nand3_4 _46610_ (.A(_16051_),
    .B(_16048_),
    .C(_16049_),
    .Y(_16053_));
 sky130_fd_sc_hd__nand2_4 _46611_ (.A(_16052_),
    .B(_16053_),
    .Y(_16054_));
 sky130_fd_sc_hd__maj3_4 _46612_ (.A(_15856_),
    .B(_15871_),
    .C(_15857_),
    .X(_16055_));
 sky130_fd_sc_hd__a21boi_4 _46613_ (.A1(_15884_),
    .A2(_15888_),
    .B1_N(_15886_),
    .Y(_16056_));
 sky130_fd_sc_hd__nand2_4 _46614_ (.A(_11319_),
    .B(_10885_),
    .Y(_16057_));
 sky130_fd_sc_hd__nand2_4 _46615_ (.A(_10715_),
    .B(_11829_),
    .Y(_16058_));
 sky130_fd_sc_hd__nand2_4 _46616_ (.A(_16057_),
    .B(_16058_),
    .Y(_16059_));
 sky130_fd_sc_hd__nand4_4 _46617_ (.A(_10827_),
    .B(_10843_),
    .C(_11502_),
    .D(_11167_),
    .Y(_16060_));
 sky130_fd_sc_hd__nand2_4 _46618_ (.A(_11334_),
    .B(_08635_),
    .Y(_16061_));
 sky130_vsdinv _46619_ (.A(_16061_),
    .Y(_16062_));
 sky130_fd_sc_hd__a21o_4 _46620_ (.A1(_16059_),
    .A2(_16060_),
    .B1(_16062_),
    .X(_16063_));
 sky130_fd_sc_hd__nand3_4 _46621_ (.A(_16059_),
    .B(_16060_),
    .C(_16062_),
    .Y(_16064_));
 sky130_fd_sc_hd__nand2_4 _46622_ (.A(_16063_),
    .B(_16064_),
    .Y(_16065_));
 sky130_fd_sc_hd__nor2_4 _46623_ (.A(_16056_),
    .B(_16065_),
    .Y(_16066_));
 sky130_vsdinv _46624_ (.A(_16066_),
    .Y(_16067_));
 sky130_fd_sc_hd__nand2_4 _46625_ (.A(_16065_),
    .B(_16056_),
    .Y(_16068_));
 sky130_fd_sc_hd__nand2_4 _46626_ (.A(_14204_),
    .B(_13055_),
    .Y(_16069_));
 sky130_fd_sc_hd__nand2_4 _46627_ (.A(_11691_),
    .B(_03552_),
    .Y(_16070_));
 sky130_fd_sc_hd__xnor2_4 _46628_ (.A(_16069_),
    .B(_16070_),
    .Y(_16071_));
 sky130_fd_sc_hd__xor2_4 _46629_ (.A(_15896_),
    .B(_16071_),
    .X(_16072_));
 sky130_fd_sc_hd__a21o_4 _46630_ (.A1(_16067_),
    .A2(_16068_),
    .B1(_16072_),
    .X(_16073_));
 sky130_fd_sc_hd__nand3_4 _46631_ (.A(_16072_),
    .B(_16068_),
    .C(_16067_),
    .Y(_16074_));
 sky130_fd_sc_hd__nand2_4 _46632_ (.A(_16073_),
    .B(_16074_),
    .Y(_16075_));
 sky130_fd_sc_hd__or2_4 _46633_ (.A(_16055_),
    .B(_16075_),
    .X(_16076_));
 sky130_fd_sc_hd__nand2_4 _46634_ (.A(_16075_),
    .B(_16055_),
    .Y(_16077_));
 sky130_fd_sc_hd__a21boi_4 _46635_ (.A1(_15902_),
    .A2(_15893_),
    .B1_N(_15894_),
    .Y(_16078_));
 sky130_vsdinv _46636_ (.A(_16078_),
    .Y(_16079_));
 sky130_fd_sc_hd__a21o_4 _46637_ (.A1(_16076_),
    .A2(_16077_),
    .B1(_16079_),
    .X(_16080_));
 sky130_fd_sc_hd__nand3_4 _46638_ (.A(_16076_),
    .B(_16079_),
    .C(_16077_),
    .Y(_16081_));
 sky130_fd_sc_hd__and2_4 _46639_ (.A(_16080_),
    .B(_16081_),
    .X(_16082_));
 sky130_vsdinv _46640_ (.A(_16082_),
    .Y(_16083_));
 sky130_fd_sc_hd__nand2_4 _46641_ (.A(_16054_),
    .B(_16083_),
    .Y(_16084_));
 sky130_fd_sc_hd__nand3_4 _46642_ (.A(_16052_),
    .B(_16082_),
    .C(_16053_),
    .Y(_16085_));
 sky130_fd_sc_hd__nand2_4 _46643_ (.A(_16084_),
    .B(_16085_),
    .Y(_16086_));
 sky130_fd_sc_hd__o21ai_4 _46644_ (.A1(_15912_),
    .A2(_15878_),
    .B1(_15880_),
    .Y(_16087_));
 sky130_vsdinv _46645_ (.A(_16087_),
    .Y(_16088_));
 sky130_fd_sc_hd__nand2_4 _46646_ (.A(_16086_),
    .B(_16088_),
    .Y(_16089_));
 sky130_fd_sc_hd__nand3_4 _46647_ (.A(_16084_),
    .B(_16087_),
    .C(_16085_),
    .Y(_16090_));
 sky130_fd_sc_hd__maj3_4 _46648_ (.A(_15898_),
    .B(_15900_),
    .C(_15896_),
    .X(_16091_));
 sky130_fd_sc_hd__xor2_4 _46649_ (.A(_16091_),
    .B(_15922_),
    .X(_16092_));
 sky130_fd_sc_hd__a21o_4 _46650_ (.A1(_15927_),
    .A2(_15925_),
    .B1(_16092_),
    .X(_16093_));
 sky130_fd_sc_hd__buf_1 _46651_ (.A(_15928_),
    .X(_16094_));
 sky130_fd_sc_hd__nand2_4 _46652_ (.A(_16092_),
    .B(_16094_),
    .Y(_16095_));
 sky130_fd_sc_hd__nand2_4 _46653_ (.A(_16093_),
    .B(_16095_),
    .Y(_16096_));
 sky130_fd_sc_hd__maj3_4 _46654_ (.A(_15920_),
    .B(_15923_),
    .C(_15928_),
    .X(_16097_));
 sky130_fd_sc_hd__nand2_4 _46655_ (.A(_16096_),
    .B(_16097_),
    .Y(_16098_));
 sky130_vsdinv _46656_ (.A(_16097_),
    .Y(_16099_));
 sky130_fd_sc_hd__nand3_4 _46657_ (.A(_16093_),
    .B(_16099_),
    .C(_16095_),
    .Y(_16100_));
 sky130_fd_sc_hd__a21o_4 _46658_ (.A1(_16098_),
    .A2(_16100_),
    .B1(_15571_),
    .X(_16101_));
 sky130_fd_sc_hd__nand3_4 _46659_ (.A(_16098_),
    .B(_16100_),
    .C(_15767_),
    .Y(_16102_));
 sky130_fd_sc_hd__maj3_4 _46660_ (.A(_15908_),
    .B(_15905_),
    .C(_15882_),
    .X(_16103_));
 sky130_vsdinv _46661_ (.A(_16103_),
    .Y(_16104_));
 sky130_fd_sc_hd__a21o_4 _46662_ (.A1(_16101_),
    .A2(_16102_),
    .B1(_16104_),
    .X(_16105_));
 sky130_fd_sc_hd__nand3_4 _46663_ (.A(_16101_),
    .B(_16104_),
    .C(_16102_),
    .Y(_16106_));
 sky130_fd_sc_hd__a21boi_4 _46664_ (.A1(_15934_),
    .A2(_15943_),
    .B1_N(_15936_),
    .Y(_16107_));
 sky130_vsdinv _46665_ (.A(_16107_),
    .Y(_16108_));
 sky130_fd_sc_hd__a21oi_4 _46666_ (.A1(_16105_),
    .A2(_16106_),
    .B1(_16108_),
    .Y(_16109_));
 sky130_fd_sc_hd__nand3_4 _46667_ (.A(_16105_),
    .B(_16108_),
    .C(_16106_),
    .Y(_16110_));
 sky130_vsdinv _46668_ (.A(_16110_),
    .Y(_16111_));
 sky130_fd_sc_hd__nor2_4 _46669_ (.A(_16109_),
    .B(_16111_),
    .Y(_16112_));
 sky130_fd_sc_hd__a21o_4 _46670_ (.A1(_16089_),
    .A2(_16090_),
    .B1(_16112_),
    .X(_16113_));
 sky130_fd_sc_hd__nand3_4 _46671_ (.A(_16112_),
    .B(_16089_),
    .C(_16090_),
    .Y(_16114_));
 sky130_fd_sc_hd__nand2_4 _46672_ (.A(_16113_),
    .B(_16114_),
    .Y(_16115_));
 sky130_fd_sc_hd__a21boi_4 _46673_ (.A1(_15918_),
    .A2(_15952_),
    .B1_N(_15916_),
    .Y(_16116_));
 sky130_fd_sc_hd__nand2_4 _46674_ (.A(_16115_),
    .B(_16116_),
    .Y(_16117_));
 sky130_fd_sc_hd__nand2_4 _46675_ (.A(_15953_),
    .B(_15916_),
    .Y(_16118_));
 sky130_fd_sc_hd__nand3_4 _46676_ (.A(_16118_),
    .B(_16114_),
    .C(_16113_),
    .Y(_16119_));
 sky130_fd_sc_hd__nand2_4 _46677_ (.A(_16117_),
    .B(_16119_),
    .Y(_16120_));
 sky130_fd_sc_hd__a21o_4 _46678_ (.A1(_15948_),
    .A2(_15942_),
    .B1(_15961_),
    .X(_16121_));
 sky130_fd_sc_hd__nand3_4 _46679_ (.A(_15948_),
    .B(_15961_),
    .C(_15942_),
    .Y(_16122_));
 sky130_fd_sc_hd__buf_1 _46680_ (.A(_15965_),
    .X(_16123_));
 sky130_fd_sc_hd__a21oi_4 _46681_ (.A1(_16121_),
    .A2(_16122_),
    .B1(_16123_),
    .Y(_16124_));
 sky130_fd_sc_hd__nand3_4 _46682_ (.A(_16121_),
    .B(_15966_),
    .C(_16122_),
    .Y(_16125_));
 sky130_vsdinv _46683_ (.A(_16125_),
    .Y(_16126_));
 sky130_fd_sc_hd__nor2_4 _46684_ (.A(_16124_),
    .B(_16126_),
    .Y(_16127_));
 sky130_vsdinv _46685_ (.A(_16127_),
    .Y(_16128_));
 sky130_fd_sc_hd__nand2_4 _46686_ (.A(_16120_),
    .B(_16128_),
    .Y(_16129_));
 sky130_fd_sc_hd__nand3_4 _46687_ (.A(_16117_),
    .B(_16119_),
    .C(_16127_),
    .Y(_16130_));
 sky130_fd_sc_hd__nand2_4 _46688_ (.A(_16129_),
    .B(_16130_),
    .Y(_16131_));
 sky130_fd_sc_hd__a21boi_4 _46689_ (.A1(_15956_),
    .A2(_15969_),
    .B1_N(_15958_),
    .Y(_16132_));
 sky130_fd_sc_hd__nand2_4 _46690_ (.A(_16131_),
    .B(_16132_),
    .Y(_16133_));
 sky130_fd_sc_hd__nand2_4 _46691_ (.A(_15972_),
    .B(_15958_),
    .Y(_16134_));
 sky130_fd_sc_hd__nand3_4 _46692_ (.A(_16134_),
    .B(_16130_),
    .C(_16129_),
    .Y(_16135_));
 sky130_fd_sc_hd__nand2_4 _46693_ (.A(_16133_),
    .B(_16135_),
    .Y(_16136_));
 sky130_fd_sc_hd__nand2_4 _46694_ (.A(_15968_),
    .B(_15960_),
    .Y(_16137_));
 sky130_fd_sc_hd__xor2_4 _46695_ (.A(_15801_),
    .B(_16137_),
    .X(_16138_));
 sky130_vsdinv _46696_ (.A(_16138_),
    .Y(_16139_));
 sky130_fd_sc_hd__nand2_4 _46697_ (.A(_16136_),
    .B(_16139_),
    .Y(_16140_));
 sky130_fd_sc_hd__nand3_4 _46698_ (.A(_16133_),
    .B(_16135_),
    .C(_16138_),
    .Y(_16141_));
 sky130_fd_sc_hd__nand2_4 _46699_ (.A(_16140_),
    .B(_16141_),
    .Y(_16142_));
 sky130_fd_sc_hd__a21boi_4 _46700_ (.A1(_15975_),
    .A2(_15981_),
    .B1_N(_15978_),
    .Y(_16143_));
 sky130_fd_sc_hd__nand2_4 _46701_ (.A(_16142_),
    .B(_16143_),
    .Y(_16144_));
 sky130_fd_sc_hd__nand2_4 _46702_ (.A(_15984_),
    .B(_15978_),
    .Y(_16145_));
 sky130_fd_sc_hd__nand3_4 _46703_ (.A(_16145_),
    .B(_16141_),
    .C(_16140_),
    .Y(_16146_));
 sky130_fd_sc_hd__nand2_4 _46704_ (.A(_16144_),
    .B(_16146_),
    .Y(_16147_));
 sky130_fd_sc_hd__buf_8 _46705_ (.A(_15440_),
    .X(_16148_));
 sky130_fd_sc_hd__buf_1 _46706_ (.A(_16148_),
    .X(_16149_));
 sky130_fd_sc_hd__buf_1 _46707_ (.A(_16149_),
    .X(_16150_));
 sky130_fd_sc_hd__and2_4 _46708_ (.A(_15980_),
    .B(_16150_),
    .X(_16151_));
 sky130_vsdinv _46709_ (.A(_16151_),
    .Y(_16152_));
 sky130_fd_sc_hd__nand2_4 _46710_ (.A(_16147_),
    .B(_16152_),
    .Y(_16153_));
 sky130_fd_sc_hd__nand3_4 _46711_ (.A(_16144_),
    .B(_16146_),
    .C(_16151_),
    .Y(_16154_));
 sky130_fd_sc_hd__nand2_4 _46712_ (.A(_16153_),
    .B(_16154_),
    .Y(_16155_));
 sky130_fd_sc_hd__a21boi_4 _46713_ (.A1(_15987_),
    .A2(_15991_),
    .B1_N(_15989_),
    .Y(_16156_));
 sky130_fd_sc_hd__nand2_4 _46714_ (.A(_16155_),
    .B(_16156_),
    .Y(_16157_));
 sky130_fd_sc_hd__nand2_4 _46715_ (.A(_15994_),
    .B(_15989_),
    .Y(_16158_));
 sky130_fd_sc_hd__nand3_4 _46716_ (.A(_16158_),
    .B(_16154_),
    .C(_16153_),
    .Y(_16159_));
 sky130_fd_sc_hd__and2_4 _46717_ (.A(_16157_),
    .B(_16159_),
    .X(_16160_));
 sky130_fd_sc_hd__buf_1 _46718_ (.A(_16160_),
    .X(_16161_));
 sky130_fd_sc_hd__o21ai_4 _46719_ (.A1(_16002_),
    .A2(_16007_),
    .B1(_15999_),
    .Y(_16162_));
 sky130_fd_sc_hd__xor2_4 _46720_ (.A(_16161_),
    .B(_16162_),
    .X(_01456_));
 sky130_fd_sc_hd__nand2_4 _46721_ (.A(_08754_),
    .B(_15250_),
    .Y(_16163_));
 sky130_fd_sc_hd__o21ai_4 _46722_ (.A1(_11910_),
    .A2(_15249_),
    .B1(_16163_),
    .Y(_16164_));
 sky130_fd_sc_hd__nand4_4 _46723_ (.A(_03348_),
    .B(_13610_),
    .C(_15659_),
    .D(_15253_),
    .Y(_16165_));
 sky130_fd_sc_hd__nand2_4 _46724_ (.A(_14140_),
    .B(_03621_),
    .Y(_16166_));
 sky130_vsdinv _46725_ (.A(_16166_),
    .Y(_16167_));
 sky130_fd_sc_hd__a21o_4 _46726_ (.A1(_16164_),
    .A2(_16165_),
    .B1(_16167_),
    .X(_16168_));
 sky130_fd_sc_hd__nand3_4 _46727_ (.A(_16164_),
    .B(_16165_),
    .C(_16167_),
    .Y(_16169_));
 sky130_fd_sc_hd__a21boi_4 _46728_ (.A1(_16009_),
    .A2(_16012_),
    .B1_N(_16010_),
    .Y(_16170_));
 sky130_fd_sc_hd__a21boi_4 _46729_ (.A1(_16168_),
    .A2(_16169_),
    .B1_N(_16170_),
    .Y(_16171_));
 sky130_vsdinv _46730_ (.A(_16171_),
    .Y(_16172_));
 sky130_vsdinv _46731_ (.A(_16170_),
    .Y(_16173_));
 sky130_fd_sc_hd__nand3_4 _46732_ (.A(_16173_),
    .B(_16168_),
    .C(_16169_),
    .Y(_16174_));
 sky130_fd_sc_hd__nand2_4 _46733_ (.A(_12233_),
    .B(_10513_),
    .Y(_16175_));
 sky130_fd_sc_hd__nand2_4 _46734_ (.A(_12226_),
    .B(_15268_),
    .Y(_16176_));
 sky130_fd_sc_hd__nand2_4 _46735_ (.A(_12231_),
    .B(_15267_),
    .Y(_16177_));
 sky130_fd_sc_hd__nand2_4 _46736_ (.A(_16176_),
    .B(_16177_),
    .Y(_16178_));
 sky130_fd_sc_hd__buf_1 _46737_ (.A(_15496_),
    .X(_16179_));
 sky130_fd_sc_hd__buf_1 _46738_ (.A(_12231_),
    .X(_16180_));
 sky130_fd_sc_hd__nand4_4 _46739_ (.A(_16179_),
    .B(_16180_),
    .C(_03608_),
    .D(_03615_),
    .Y(_16181_));
 sky130_fd_sc_hd__nand2_4 _46740_ (.A(_16178_),
    .B(_16181_),
    .Y(_16182_));
 sky130_fd_sc_hd__xor2_4 _46741_ (.A(_16175_),
    .B(_16182_),
    .X(_16183_));
 sky130_fd_sc_hd__a21o_4 _46742_ (.A1(_16172_),
    .A2(_16174_),
    .B1(_16183_),
    .X(_16184_));
 sky130_fd_sc_hd__nand3_4 _46743_ (.A(_16172_),
    .B(_16174_),
    .C(_16183_),
    .Y(_16185_));
 sky130_fd_sc_hd__a21boi_4 _46744_ (.A1(_16017_),
    .A2(_16025_),
    .B1_N(_16018_),
    .Y(_16186_));
 sky130_vsdinv _46745_ (.A(_16186_),
    .Y(_16187_));
 sky130_fd_sc_hd__a21oi_4 _46746_ (.A1(_16184_),
    .A2(_16185_),
    .B1(_16187_),
    .Y(_16188_));
 sky130_fd_sc_hd__nand3_4 _46747_ (.A(_16187_),
    .B(_16184_),
    .C(_16185_),
    .Y(_16189_));
 sky130_vsdinv _46748_ (.A(_16189_),
    .Y(_16190_));
 sky130_fd_sc_hd__nand2_4 _46749_ (.A(_13114_),
    .B(_15494_),
    .Y(_16191_));
 sky130_fd_sc_hd__nand2_4 _46750_ (.A(_13127_),
    .B(_03588_),
    .Y(_16192_));
 sky130_fd_sc_hd__nand2_4 _46751_ (.A(_16191_),
    .B(_16192_),
    .Y(_16193_));
 sky130_fd_sc_hd__nand4_4 _46752_ (.A(_14884_),
    .B(_14882_),
    .C(_13842_),
    .D(_03597_),
    .Y(_16194_));
 sky130_fd_sc_hd__buf_1 _46753_ (.A(_11473_),
    .X(_16195_));
 sky130_fd_sc_hd__nand2_4 _46754_ (.A(_12279_),
    .B(_16195_),
    .Y(_16196_));
 sky130_vsdinv _46755_ (.A(_16196_),
    .Y(_16197_));
 sky130_fd_sc_hd__a21o_4 _46756_ (.A1(_16193_),
    .A2(_16194_),
    .B1(_16197_),
    .X(_16198_));
 sky130_fd_sc_hd__nand3_4 _46757_ (.A(_16193_),
    .B(_16194_),
    .C(_16197_),
    .Y(_16199_));
 sky130_vsdinv _46758_ (.A(_16019_),
    .Y(_16200_));
 sky130_fd_sc_hd__a21boi_4 _46759_ (.A1(_16022_),
    .A2(_16200_),
    .B1_N(_16023_),
    .Y(_16201_));
 sky130_fd_sc_hd__a21boi_4 _46760_ (.A1(_16198_),
    .A2(_16199_),
    .B1_N(_16201_),
    .Y(_16202_));
 sky130_vsdinv _46761_ (.A(_16202_),
    .Y(_16203_));
 sky130_vsdinv _46762_ (.A(_16201_),
    .Y(_16204_));
 sky130_fd_sc_hd__nand3_4 _46763_ (.A(_16204_),
    .B(_16198_),
    .C(_16199_),
    .Y(_16205_));
 sky130_fd_sc_hd__a21boi_4 _46764_ (.A1(_16036_),
    .A2(_16042_),
    .B1_N(_16039_),
    .Y(_16206_));
 sky130_vsdinv _46765_ (.A(_16206_),
    .Y(_16207_));
 sky130_fd_sc_hd__a21oi_4 _46766_ (.A1(_16203_),
    .A2(_16205_),
    .B1(_16207_),
    .Y(_16208_));
 sky130_fd_sc_hd__nand3_4 _46767_ (.A(_16203_),
    .B(_16207_),
    .C(_16205_),
    .Y(_16209_));
 sky130_vsdinv _46768_ (.A(_16209_),
    .Y(_16210_));
 sky130_fd_sc_hd__nor2_4 _46769_ (.A(_16208_),
    .B(_16210_),
    .Y(_16211_));
 sky130_vsdinv _46770_ (.A(_16211_),
    .Y(_16212_));
 sky130_fd_sc_hd__o21ai_4 _46771_ (.A1(_16188_),
    .A2(_16190_),
    .B1(_16212_),
    .Y(_16213_));
 sky130_vsdinv _46772_ (.A(_16188_),
    .Y(_16214_));
 sky130_fd_sc_hd__nand3_4 _46773_ (.A(_16214_),
    .B(_16189_),
    .C(_16211_),
    .Y(_16215_));
 sky130_fd_sc_hd__a21boi_4 _46774_ (.A1(_16030_),
    .A2(_16047_),
    .B1_N(_16031_),
    .Y(_16216_));
 sky130_fd_sc_hd__a21boi_4 _46775_ (.A1(_16213_),
    .A2(_16215_),
    .B1_N(_16216_),
    .Y(_16217_));
 sky130_vsdinv _46776_ (.A(_16217_),
    .Y(_16218_));
 sky130_vsdinv _46777_ (.A(_16216_),
    .Y(_16219_));
 sky130_fd_sc_hd__nand3_4 _46778_ (.A(_16219_),
    .B(_16213_),
    .C(_16215_),
    .Y(_16220_));
 sky130_fd_sc_hd__a21oi_4 _46779_ (.A1(_16072_),
    .A2(_16068_),
    .B1(_16066_),
    .Y(_16221_));
 sky130_vsdinv _46780_ (.A(_16221_),
    .Y(_16222_));
 sky130_fd_sc_hd__maj3_4 _46781_ (.A(_16032_),
    .B(_16045_),
    .C(_16033_),
    .X(_16223_));
 sky130_fd_sc_hd__nand2_4 _46782_ (.A(_15136_),
    .B(_14867_),
    .Y(_16224_));
 sky130_fd_sc_hd__nand2_4 _46783_ (.A(_13410_),
    .B(_14869_),
    .Y(_16225_));
 sky130_fd_sc_hd__nand2_4 _46784_ (.A(_16224_),
    .B(_16225_),
    .Y(_16226_));
 sky130_fd_sc_hd__nand4_4 _46785_ (.A(_10840_),
    .B(_03397_),
    .C(_14869_),
    .D(_14867_),
    .Y(_16227_));
 sky130_fd_sc_hd__nand2_4 _46786_ (.A(_10837_),
    .B(_08636_),
    .Y(_16228_));
 sky130_vsdinv _46787_ (.A(_16228_),
    .Y(_16229_));
 sky130_fd_sc_hd__a21o_4 _46788_ (.A1(_16226_),
    .A2(_16227_),
    .B1(_16229_),
    .X(_16230_));
 sky130_fd_sc_hd__nand3_4 _46789_ (.A(_16226_),
    .B(_16227_),
    .C(_16229_),
    .Y(_16231_));
 sky130_fd_sc_hd__a21boi_4 _46790_ (.A1(_16059_),
    .A2(_16062_),
    .B1_N(_16060_),
    .Y(_16232_));
 sky130_vsdinv _46791_ (.A(_16232_),
    .Y(_16233_));
 sky130_fd_sc_hd__a21o_4 _46792_ (.A1(_16230_),
    .A2(_16231_),
    .B1(_16233_),
    .X(_16234_));
 sky130_fd_sc_hd__nand3_4 _46793_ (.A(_16233_),
    .B(_16230_),
    .C(_16231_),
    .Y(_16235_));
 sky130_vsdinv _46794_ (.A(_15895_),
    .Y(_16236_));
 sky130_fd_sc_hd__nand2_4 _46795_ (.A(_03406_),
    .B(_09486_),
    .Y(_16237_));
 sky130_fd_sc_hd__nand2_4 _46796_ (.A(_16070_),
    .B(_16237_),
    .Y(_16238_));
 sky130_fd_sc_hd__nand3_4 _46797_ (.A(_12909_),
    .B(_12762_),
    .C(_08198_),
    .Y(_16239_));
 sky130_fd_sc_hd__and2_4 _46798_ (.A(_16238_),
    .B(_16239_),
    .X(_16240_));
 sky130_fd_sc_hd__xor2_4 _46799_ (.A(_16236_),
    .B(_16240_),
    .X(_16241_));
 sky130_fd_sc_hd__buf_1 _46800_ (.A(_16241_),
    .X(_16242_));
 sky130_fd_sc_hd__a21o_4 _46801_ (.A1(_16234_),
    .A2(_16235_),
    .B1(_16242_),
    .X(_16243_));
 sky130_fd_sc_hd__buf_1 _46802_ (.A(_16242_),
    .X(_16244_));
 sky130_fd_sc_hd__nand3_4 _46803_ (.A(_16244_),
    .B(_16234_),
    .C(_16235_),
    .Y(_16245_));
 sky130_fd_sc_hd__nand2_4 _46804_ (.A(_16243_),
    .B(_16245_),
    .Y(_16246_));
 sky130_fd_sc_hd__xnor2_4 _46805_ (.A(_16223_),
    .B(_16246_),
    .Y(_16247_));
 sky130_fd_sc_hd__xor2_4 _46806_ (.A(_16222_),
    .B(_16247_),
    .X(_16248_));
 sky130_vsdinv _46807_ (.A(_16248_),
    .Y(_16249_));
 sky130_fd_sc_hd__a21o_4 _46808_ (.A1(_16218_),
    .A2(_16220_),
    .B1(_16249_),
    .X(_16250_));
 sky130_fd_sc_hd__nand3_4 _46809_ (.A(_16249_),
    .B(_16218_),
    .C(_16220_),
    .Y(_16251_));
 sky130_fd_sc_hd__a21boi_4 _46810_ (.A1(_16052_),
    .A2(_16082_),
    .B1_N(_16053_),
    .Y(_16252_));
 sky130_fd_sc_hd__a21boi_4 _46811_ (.A1(_16250_),
    .A2(_16251_),
    .B1_N(_16252_),
    .Y(_16253_));
 sky130_vsdinv _46812_ (.A(_16252_),
    .Y(_16254_));
 sky130_fd_sc_hd__nand3_4 _46813_ (.A(_16254_),
    .B(_16250_),
    .C(_16251_),
    .Y(_16255_));
 sky130_vsdinv _46814_ (.A(_16255_),
    .Y(_16256_));
 sky130_fd_sc_hd__maj3_4 _46815_ (.A(_15896_),
    .B(_16069_),
    .C(_16070_),
    .X(_16257_));
 sky130_fd_sc_hd__xor2_4 _46816_ (.A(_16257_),
    .B(_15922_),
    .X(_16258_));
 sky130_fd_sc_hd__a21o_4 _46817_ (.A1(_15927_),
    .A2(_15925_),
    .B1(_16258_),
    .X(_16259_));
 sky130_fd_sc_hd__nand2_4 _46818_ (.A(_16258_),
    .B(_16094_),
    .Y(_16260_));
 sky130_fd_sc_hd__maj3_4 _46819_ (.A(_16094_),
    .B(_15923_),
    .C(_16091_),
    .X(_16261_));
 sky130_vsdinv _46820_ (.A(_16261_),
    .Y(_16262_));
 sky130_fd_sc_hd__a21o_4 _46821_ (.A1(_16259_),
    .A2(_16260_),
    .B1(_16262_),
    .X(_16263_));
 sky130_fd_sc_hd__nand3_4 _46822_ (.A(_16259_),
    .B(_16262_),
    .C(_16260_),
    .Y(_16264_));
 sky130_fd_sc_hd__a21o_4 _46823_ (.A1(_16263_),
    .A2(_16264_),
    .B1(_15943_),
    .X(_16265_));
 sky130_fd_sc_hd__buf_1 _46824_ (.A(_15762_),
    .X(_16266_));
 sky130_fd_sc_hd__nand3_4 _46825_ (.A(_16263_),
    .B(_16266_),
    .C(_16264_),
    .Y(_16267_));
 sky130_fd_sc_hd__maj3_4 _46826_ (.A(_16078_),
    .B(_16075_),
    .C(_16055_),
    .X(_16268_));
 sky130_vsdinv _46827_ (.A(_16268_),
    .Y(_16269_));
 sky130_fd_sc_hd__a21o_4 _46828_ (.A1(_16265_),
    .A2(_16267_),
    .B1(_16269_),
    .X(_16270_));
 sky130_fd_sc_hd__nand3_4 _46829_ (.A(_16265_),
    .B(_16269_),
    .C(_16267_),
    .Y(_16271_));
 sky130_fd_sc_hd__a21boi_4 _46830_ (.A1(_16098_),
    .A2(_16266_),
    .B1_N(_16100_),
    .Y(_16272_));
 sky130_vsdinv _46831_ (.A(_16272_),
    .Y(_16273_));
 sky130_fd_sc_hd__a21oi_4 _46832_ (.A1(_16270_),
    .A2(_16271_),
    .B1(_16273_),
    .Y(_16274_));
 sky130_vsdinv _46833_ (.A(_16274_),
    .Y(_16275_));
 sky130_fd_sc_hd__nand3_4 _46834_ (.A(_16270_),
    .B(_16273_),
    .C(_16271_),
    .Y(_16276_));
 sky130_fd_sc_hd__nand2_4 _46835_ (.A(_16275_),
    .B(_16276_),
    .Y(_16277_));
 sky130_fd_sc_hd__o21ai_4 _46836_ (.A1(_16253_),
    .A2(_16256_),
    .B1(_16277_),
    .Y(_16278_));
 sky130_vsdinv _46837_ (.A(_16253_),
    .Y(_16279_));
 sky130_fd_sc_hd__nand4_4 _46838_ (.A(_16279_),
    .B(_16255_),
    .C(_16276_),
    .D(_16275_),
    .Y(_16280_));
 sky130_fd_sc_hd__nand2_4 _46839_ (.A(_16278_),
    .B(_16280_),
    .Y(_16281_));
 sky130_fd_sc_hd__a21boi_4 _46840_ (.A1(_16112_),
    .A2(_16089_),
    .B1_N(_16090_),
    .Y(_16282_));
 sky130_fd_sc_hd__nand2_4 _46841_ (.A(_16281_),
    .B(_16282_),
    .Y(_16283_));
 sky130_vsdinv _46842_ (.A(_16282_),
    .Y(_16284_));
 sky130_fd_sc_hd__nand3_4 _46843_ (.A(_16284_),
    .B(_16278_),
    .C(_16280_),
    .Y(_16285_));
 sky130_fd_sc_hd__nand2_4 _46844_ (.A(_16283_),
    .B(_16285_),
    .Y(_16286_));
 sky130_fd_sc_hd__a21o_4 _46845_ (.A1(_16110_),
    .A2(_16106_),
    .B1(_15962_),
    .X(_16287_));
 sky130_fd_sc_hd__buf_1 _46846_ (.A(_15961_),
    .X(_16288_));
 sky130_fd_sc_hd__nand3_4 _46847_ (.A(_16110_),
    .B(_16288_),
    .C(_16106_),
    .Y(_16289_));
 sky130_fd_sc_hd__buf_1 _46848_ (.A(_15966_),
    .X(_16290_));
 sky130_fd_sc_hd__a21o_4 _46849_ (.A1(_16287_),
    .A2(_16289_),
    .B1(_16290_),
    .X(_16291_));
 sky130_fd_sc_hd__nand3_4 _46850_ (.A(_16287_),
    .B(_16123_),
    .C(_16289_),
    .Y(_16292_));
 sky130_fd_sc_hd__nand2_4 _46851_ (.A(_16291_),
    .B(_16292_),
    .Y(_16293_));
 sky130_fd_sc_hd__nand2_4 _46852_ (.A(_16286_),
    .B(_16293_),
    .Y(_16294_));
 sky130_vsdinv _46853_ (.A(_16293_),
    .Y(_16295_));
 sky130_fd_sc_hd__nand3_4 _46854_ (.A(_16283_),
    .B(_16285_),
    .C(_16295_),
    .Y(_16296_));
 sky130_fd_sc_hd__nand2_4 _46855_ (.A(_16294_),
    .B(_16296_),
    .Y(_16297_));
 sky130_fd_sc_hd__a21boi_4 _46856_ (.A1(_16117_),
    .A2(_16127_),
    .B1_N(_16119_),
    .Y(_16298_));
 sky130_fd_sc_hd__nand2_4 _46857_ (.A(_16297_),
    .B(_16298_),
    .Y(_16299_));
 sky130_vsdinv _46858_ (.A(_16298_),
    .Y(_16300_));
 sky130_fd_sc_hd__nand3_4 _46859_ (.A(_16300_),
    .B(_16294_),
    .C(_16296_),
    .Y(_16301_));
 sky130_fd_sc_hd__nand2_4 _46860_ (.A(_16299_),
    .B(_16301_),
    .Y(_16302_));
 sky130_fd_sc_hd__nand2_4 _46861_ (.A(_16125_),
    .B(_16121_),
    .Y(_16303_));
 sky130_fd_sc_hd__xor2_4 _46862_ (.A(_15801_),
    .B(_16303_),
    .X(_16304_));
 sky130_vsdinv _46863_ (.A(_16304_),
    .Y(_16305_));
 sky130_fd_sc_hd__nand2_4 _46864_ (.A(_16302_),
    .B(_16305_),
    .Y(_16306_));
 sky130_fd_sc_hd__nand3_4 _46865_ (.A(_16299_),
    .B(_16301_),
    .C(_16304_),
    .Y(_16307_));
 sky130_fd_sc_hd__nand2_4 _46866_ (.A(_16306_),
    .B(_16307_),
    .Y(_16308_));
 sky130_fd_sc_hd__nand2_4 _46867_ (.A(_16141_),
    .B(_16135_),
    .Y(_16309_));
 sky130_vsdinv _46868_ (.A(_16309_),
    .Y(_16310_));
 sky130_fd_sc_hd__nand2_4 _46869_ (.A(_16308_),
    .B(_16310_),
    .Y(_16311_));
 sky130_fd_sc_hd__nand3_4 _46870_ (.A(_16306_),
    .B(_16309_),
    .C(_16307_),
    .Y(_16312_));
 sky130_fd_sc_hd__nand2_4 _46871_ (.A(_16311_),
    .B(_16312_),
    .Y(_16313_));
 sky130_fd_sc_hd__buf_1 _46872_ (.A(_15452_),
    .X(_16314_));
 sky130_fd_sc_hd__a21oi_4 _46873_ (.A1(_15968_),
    .A2(_15960_),
    .B1(_16314_),
    .Y(_16315_));
 sky130_vsdinv _46874_ (.A(_16315_),
    .Y(_16316_));
 sky130_fd_sc_hd__nand2_4 _46875_ (.A(_16313_),
    .B(_16316_),
    .Y(_16317_));
 sky130_fd_sc_hd__nand3_4 _46876_ (.A(_16311_),
    .B(_16315_),
    .C(_16312_),
    .Y(_16318_));
 sky130_fd_sc_hd__nand2_4 _46877_ (.A(_16317_),
    .B(_16318_),
    .Y(_16319_));
 sky130_fd_sc_hd__nand2_4 _46878_ (.A(_16154_),
    .B(_16146_),
    .Y(_16320_));
 sky130_vsdinv _46879_ (.A(_16320_),
    .Y(_16321_));
 sky130_fd_sc_hd__nand2_4 _46880_ (.A(_16319_),
    .B(_16321_),
    .Y(_16322_));
 sky130_fd_sc_hd__nand3_4 _46881_ (.A(_16317_),
    .B(_16320_),
    .C(_16318_),
    .Y(_16323_));
 sky130_fd_sc_hd__and2_4 _46882_ (.A(_16322_),
    .B(_16323_),
    .X(_16324_));
 sky130_fd_sc_hd__buf_1 _46883_ (.A(_16324_),
    .X(_16325_));
 sky130_vsdinv _46884_ (.A(_16325_),
    .Y(_16326_));
 sky130_fd_sc_hd__nand4_4 _46885_ (.A(_15636_),
    .B(_16001_),
    .C(_15822_),
    .D(_16161_),
    .Y(_16327_));
 sky130_vsdinv _46886_ (.A(_16327_),
    .Y(_16328_));
 sky130_fd_sc_hd__nand2_4 _46887_ (.A(_16006_),
    .B(_16005_),
    .Y(_16329_));
 sky130_fd_sc_hd__nand4_4 _46888_ (.A(_15999_),
    .B(_15997_),
    .C(_16157_),
    .D(_16159_),
    .Y(_16330_));
 sky130_vsdinv _46889_ (.A(_15999_),
    .Y(_16331_));
 sky130_fd_sc_hd__a21boi_4 _46890_ (.A1(_16331_),
    .A2(_16157_),
    .B1_N(_16159_),
    .Y(_16332_));
 sky130_fd_sc_hd__o21ai_4 _46891_ (.A1(_16329_),
    .A2(_16330_),
    .B1(_16332_),
    .Y(_16333_));
 sky130_fd_sc_hd__a21oi_4 _46892_ (.A1(_15652_),
    .A2(_16328_),
    .B1(_16333_),
    .Y(_16334_));
 sky130_fd_sc_hd__xor2_4 _46893_ (.A(_16326_),
    .B(_16334_),
    .X(_01457_));
 sky130_fd_sc_hd__buf_1 _46894_ (.A(_15033_),
    .X(_16335_));
 sky130_fd_sc_hd__nand2_4 _46895_ (.A(_14140_),
    .B(_16335_),
    .Y(_16336_));
 sky130_fd_sc_hd__o21ai_4 _46896_ (.A1(_13610_),
    .A2(_15249_),
    .B1(_16336_),
    .Y(_16337_));
 sky130_fd_sc_hd__buf_1 _46897_ (.A(_15250_),
    .X(_16338_));
 sky130_fd_sc_hd__nand4_4 _46898_ (.A(_03355_),
    .B(_11915_),
    .C(_16338_),
    .D(_11385_),
    .Y(_16339_));
 sky130_fd_sc_hd__nand2_4 _46899_ (.A(_12226_),
    .B(_03621_),
    .Y(_16340_));
 sky130_vsdinv _46900_ (.A(_16340_),
    .Y(_16341_));
 sky130_fd_sc_hd__a21o_4 _46901_ (.A1(_16337_),
    .A2(_16339_),
    .B1(_16341_),
    .X(_16342_));
 sky130_fd_sc_hd__nand3_4 _46902_ (.A(_16337_),
    .B(_16339_),
    .C(_16341_),
    .Y(_16343_));
 sky130_fd_sc_hd__a21boi_4 _46903_ (.A1(_16164_),
    .A2(_16167_),
    .B1_N(_16165_),
    .Y(_16344_));
 sky130_vsdinv _46904_ (.A(_16344_),
    .Y(_16345_));
 sky130_fd_sc_hd__a21o_4 _46905_ (.A1(_16342_),
    .A2(_16343_),
    .B1(_16345_),
    .X(_16346_));
 sky130_fd_sc_hd__nand3_4 _46906_ (.A(_16345_),
    .B(_16342_),
    .C(_16343_),
    .Y(_16347_));
 sky130_fd_sc_hd__nand2_4 _46907_ (.A(_16038_),
    .B(_03602_),
    .Y(_16348_));
 sky130_fd_sc_hd__nand2_4 _46908_ (.A(_15863_),
    .B(_15268_),
    .Y(_16349_));
 sky130_fd_sc_hd__nand2_4 _46909_ (.A(_12824_),
    .B(_15267_),
    .Y(_16350_));
 sky130_fd_sc_hd__nand2_4 _46910_ (.A(_16349_),
    .B(_16350_),
    .Y(_16351_));
 sky130_fd_sc_hd__nand4_4 _46911_ (.A(_16180_),
    .B(_16037_),
    .C(_03608_),
    .D(_03615_),
    .Y(_16352_));
 sky130_fd_sc_hd__nand2_4 _46912_ (.A(_16351_),
    .B(_16352_),
    .Y(_16353_));
 sky130_fd_sc_hd__xor2_4 _46913_ (.A(_16348_),
    .B(_16353_),
    .X(_16354_));
 sky130_fd_sc_hd__a21o_4 _46914_ (.A1(_16346_),
    .A2(_16347_),
    .B1(_16354_),
    .X(_16355_));
 sky130_fd_sc_hd__nand3_4 _46915_ (.A(_16346_),
    .B(_16354_),
    .C(_16347_),
    .Y(_16356_));
 sky130_fd_sc_hd__a21boi_4 _46916_ (.A1(_16172_),
    .A2(_16183_),
    .B1_N(_16174_),
    .Y(_16357_));
 sky130_vsdinv _46917_ (.A(_16357_),
    .Y(_16358_));
 sky130_fd_sc_hd__a21o_4 _46918_ (.A1(_16355_),
    .A2(_16356_),
    .B1(_16358_),
    .X(_16359_));
 sky130_fd_sc_hd__nand3_4 _46919_ (.A(_16358_),
    .B(_16355_),
    .C(_16356_),
    .Y(_16360_));
 sky130_fd_sc_hd__a21boi_4 _46920_ (.A1(_16193_),
    .A2(_16197_),
    .B1_N(_16194_),
    .Y(_16361_));
 sky130_fd_sc_hd__maj3_4 _46921_ (.A(_16176_),
    .B(_16177_),
    .C(_16175_),
    .X(_16362_));
 sky130_fd_sc_hd__nand2_4 _46922_ (.A(_13127_),
    .B(_15494_),
    .Y(_16363_));
 sky130_fd_sc_hd__nand2_4 _46923_ (.A(_14426_),
    .B(_12721_),
    .Y(_16364_));
 sky130_fd_sc_hd__nand2_4 _46924_ (.A(_16363_),
    .B(_16364_),
    .Y(_16365_));
 sky130_fd_sc_hd__nand4_4 _46925_ (.A(_11955_),
    .B(_15885_),
    .C(_13842_),
    .D(_03597_),
    .Y(_16366_));
 sky130_fd_sc_hd__nand2_4 _46926_ (.A(_15132_),
    .B(_16195_),
    .Y(_16367_));
 sky130_vsdinv _46927_ (.A(_16367_),
    .Y(_16368_));
 sky130_fd_sc_hd__a21o_4 _46928_ (.A1(_16365_),
    .A2(_16366_),
    .B1(_16368_),
    .X(_16369_));
 sky130_fd_sc_hd__nand3_4 _46929_ (.A(_16365_),
    .B(_16366_),
    .C(_16368_),
    .Y(_16370_));
 sky130_fd_sc_hd__nand2_4 _46930_ (.A(_16369_),
    .B(_16370_),
    .Y(_16371_));
 sky130_fd_sc_hd__or2_4 _46931_ (.A(_16362_),
    .B(_16371_),
    .X(_16372_));
 sky130_fd_sc_hd__buf_1 _46932_ (.A(_16372_),
    .X(_16373_));
 sky130_fd_sc_hd__nand2_4 _46933_ (.A(_16371_),
    .B(_16362_),
    .Y(_16374_));
 sky130_fd_sc_hd__nand2_4 _46934_ (.A(_16373_),
    .B(_16374_),
    .Y(_16375_));
 sky130_fd_sc_hd__xor2_4 _46935_ (.A(_16361_),
    .B(_16375_),
    .X(_16376_));
 sky130_fd_sc_hd__a21o_4 _46936_ (.A1(_16359_),
    .A2(_16360_),
    .B1(_16376_),
    .X(_16377_));
 sky130_fd_sc_hd__nand3_4 _46937_ (.A(_16359_),
    .B(_16376_),
    .C(_16360_),
    .Y(_16378_));
 sky130_fd_sc_hd__nand2_4 _46938_ (.A(_16377_),
    .B(_16378_),
    .Y(_16379_));
 sky130_fd_sc_hd__a21o_4 _46939_ (.A1(_16189_),
    .A2(_16215_),
    .B1(_16379_),
    .X(_16380_));
 sky130_fd_sc_hd__o21a_4 _46940_ (.A1(_16212_),
    .A2(_16188_),
    .B1(_16189_),
    .X(_16381_));
 sky130_fd_sc_hd__nand2_4 _46941_ (.A(_16379_),
    .B(_16381_),
    .Y(_16382_));
 sky130_fd_sc_hd__nand2_4 _46942_ (.A(_10847_),
    .B(_14873_),
    .Y(_16383_));
 sky130_fd_sc_hd__nand2_4 _46943_ (.A(_15899_),
    .B(_14872_),
    .Y(_16384_));
 sky130_fd_sc_hd__nand2_4 _46944_ (.A(_16383_),
    .B(_16384_),
    .Y(_16385_));
 sky130_fd_sc_hd__nand4_4 _46945_ (.A(_15897_),
    .B(_15899_),
    .C(_03571_),
    .D(_14873_),
    .Y(_16386_));
 sky130_fd_sc_hd__nand2_4 _46946_ (.A(_12907_),
    .B(_08636_),
    .Y(_16387_));
 sky130_vsdinv _46947_ (.A(_16387_),
    .Y(_16388_));
 sky130_fd_sc_hd__a21o_4 _46948_ (.A1(_16385_),
    .A2(_16386_),
    .B1(_16388_),
    .X(_16389_));
 sky130_fd_sc_hd__nand3_4 _46949_ (.A(_16385_),
    .B(_16386_),
    .C(_16388_),
    .Y(_16390_));
 sky130_fd_sc_hd__a21boi_4 _46950_ (.A1(_16226_),
    .A2(_16229_),
    .B1_N(_16227_),
    .Y(_16391_));
 sky130_vsdinv _46951_ (.A(_16391_),
    .Y(_16392_));
 sky130_fd_sc_hd__a21o_4 _46952_ (.A1(_16389_),
    .A2(_16390_),
    .B1(_16392_),
    .X(_16393_));
 sky130_fd_sc_hd__nand3_4 _46953_ (.A(_16392_),
    .B(_16389_),
    .C(_16390_),
    .Y(_16394_));
 sky130_fd_sc_hd__a21o_4 _46954_ (.A1(_16393_),
    .A2(_16394_),
    .B1(_16242_),
    .X(_16395_));
 sky130_fd_sc_hd__nand3_4 _46955_ (.A(_16242_),
    .B(_16393_),
    .C(_16394_),
    .Y(_16396_));
 sky130_fd_sc_hd__nand2_4 _46956_ (.A(_16395_),
    .B(_16396_),
    .Y(_16397_));
 sky130_fd_sc_hd__a21o_4 _46957_ (.A1(_16205_),
    .A2(_16209_),
    .B1(_16397_),
    .X(_16398_));
 sky130_fd_sc_hd__nand3_4 _46958_ (.A(_16397_),
    .B(_16205_),
    .C(_16209_),
    .Y(_16399_));
 sky130_fd_sc_hd__nand2_4 _46959_ (.A(_16398_),
    .B(_16399_),
    .Y(_16400_));
 sky130_fd_sc_hd__a21o_4 _46960_ (.A1(_16235_),
    .A2(_16245_),
    .B1(_16400_),
    .X(_16401_));
 sky130_fd_sc_hd__nand3_4 _46961_ (.A(_16400_),
    .B(_16235_),
    .C(_16245_),
    .Y(_16402_));
 sky130_fd_sc_hd__nand2_4 _46962_ (.A(_16401_),
    .B(_16402_),
    .Y(_16403_));
 sky130_vsdinv _46963_ (.A(_16403_),
    .Y(_16404_));
 sky130_fd_sc_hd__a21o_4 _46964_ (.A1(_16380_),
    .A2(_16382_),
    .B1(_16404_),
    .X(_16405_));
 sky130_fd_sc_hd__nand3_4 _46965_ (.A(_16380_),
    .B(_16382_),
    .C(_16404_),
    .Y(_16406_));
 sky130_fd_sc_hd__nand2_4 _46966_ (.A(_16405_),
    .B(_16406_),
    .Y(_16407_));
 sky130_fd_sc_hd__o21a_4 _46967_ (.A1(_16217_),
    .A2(_16248_),
    .B1(_16220_),
    .X(_16408_));
 sky130_fd_sc_hd__nand2_4 _46968_ (.A(_16407_),
    .B(_16408_),
    .Y(_16409_));
 sky130_vsdinv _46969_ (.A(_16408_),
    .Y(_16410_));
 sky130_fd_sc_hd__nand3_4 _46970_ (.A(_16405_),
    .B(_16410_),
    .C(_16406_),
    .Y(_16411_));
 sky130_fd_sc_hd__nand2_4 _46971_ (.A(_16409_),
    .B(_16411_),
    .Y(_16412_));
 sky130_fd_sc_hd__a21boi_4 _46972_ (.A1(_16238_),
    .A2(_16236_),
    .B1_N(_16239_),
    .Y(_16413_));
 sky130_fd_sc_hd__xor2_4 _46973_ (.A(_16413_),
    .B(_15922_),
    .X(_16414_));
 sky130_fd_sc_hd__a21o_4 _46974_ (.A1(_15927_),
    .A2(_15925_),
    .B1(_16414_),
    .X(_16415_));
 sky130_fd_sc_hd__nand2_4 _46975_ (.A(_16414_),
    .B(_16094_),
    .Y(_16416_));
 sky130_fd_sc_hd__maj3_4 _46976_ (.A(_15928_),
    .B(_15923_),
    .C(_16257_),
    .X(_16417_));
 sky130_vsdinv _46977_ (.A(_16417_),
    .Y(_16418_));
 sky130_fd_sc_hd__a21o_4 _46978_ (.A1(_16415_),
    .A2(_16416_),
    .B1(_16418_),
    .X(_16419_));
 sky130_fd_sc_hd__nand3_4 _46979_ (.A(_16415_),
    .B(_16418_),
    .C(_16416_),
    .Y(_16420_));
 sky130_fd_sc_hd__a21o_4 _46980_ (.A1(_16419_),
    .A2(_16420_),
    .B1(_15571_),
    .X(_16421_));
 sky130_fd_sc_hd__nand3_4 _46981_ (.A(_16419_),
    .B(_15767_),
    .C(_16420_),
    .Y(_16422_));
 sky130_fd_sc_hd__maj3_4 _46982_ (.A(_16221_),
    .B(_16246_),
    .C(_16223_),
    .X(_16423_));
 sky130_vsdinv _46983_ (.A(_16423_),
    .Y(_16424_));
 sky130_fd_sc_hd__a21o_4 _46984_ (.A1(_16421_),
    .A2(_16422_),
    .B1(_16424_),
    .X(_16425_));
 sky130_fd_sc_hd__nand3_4 _46985_ (.A(_16421_),
    .B(_16424_),
    .C(_16422_),
    .Y(_16426_));
 sky130_fd_sc_hd__a21boi_4 _46986_ (.A1(_16263_),
    .A2(_15943_),
    .B1_N(_16264_),
    .Y(_16427_));
 sky130_vsdinv _46987_ (.A(_16427_),
    .Y(_16428_));
 sky130_fd_sc_hd__a21oi_4 _46988_ (.A1(_16425_),
    .A2(_16426_),
    .B1(_16428_),
    .Y(_16429_));
 sky130_fd_sc_hd__nand3_4 _46989_ (.A(_16425_),
    .B(_16428_),
    .C(_16426_),
    .Y(_16430_));
 sky130_vsdinv _46990_ (.A(_16430_),
    .Y(_16431_));
 sky130_fd_sc_hd__nor2_4 _46991_ (.A(_16429_),
    .B(_16431_),
    .Y(_16432_));
 sky130_vsdinv _46992_ (.A(_16432_),
    .Y(_16433_));
 sky130_fd_sc_hd__nand2_4 _46993_ (.A(_16412_),
    .B(_16433_),
    .Y(_16434_));
 sky130_fd_sc_hd__nand3_4 _46994_ (.A(_16409_),
    .B(_16432_),
    .C(_16411_),
    .Y(_16435_));
 sky130_fd_sc_hd__nand2_4 _46995_ (.A(_16434_),
    .B(_16435_),
    .Y(_16436_));
 sky130_fd_sc_hd__o21ai_4 _46996_ (.A1(_16253_),
    .A2(_16277_),
    .B1(_16255_),
    .Y(_16437_));
 sky130_vsdinv _46997_ (.A(_16437_),
    .Y(_16438_));
 sky130_fd_sc_hd__nand2_4 _46998_ (.A(_16436_),
    .B(_16438_),
    .Y(_16439_));
 sky130_fd_sc_hd__nand3_4 _46999_ (.A(_16437_),
    .B(_16434_),
    .C(_16435_),
    .Y(_16440_));
 sky130_fd_sc_hd__nand2_4 _47000_ (.A(_16439_),
    .B(_16440_),
    .Y(_16441_));
 sky130_fd_sc_hd__a21o_4 _47001_ (.A1(_16276_),
    .A2(_16271_),
    .B1(_15787_),
    .X(_16442_));
 sky130_fd_sc_hd__nand3_4 _47002_ (.A(_16276_),
    .B(_15962_),
    .C(_16271_),
    .Y(_16443_));
 sky130_fd_sc_hd__buf_1 _47003_ (.A(_16123_),
    .X(_16444_));
 sky130_fd_sc_hd__a21oi_4 _47004_ (.A1(_16442_),
    .A2(_16443_),
    .B1(_16444_),
    .Y(_16445_));
 sky130_fd_sc_hd__nand3_4 _47005_ (.A(_16442_),
    .B(_16443_),
    .C(_16123_),
    .Y(_16446_));
 sky130_vsdinv _47006_ (.A(_16446_),
    .Y(_16447_));
 sky130_fd_sc_hd__nor2_4 _47007_ (.A(_16445_),
    .B(_16447_),
    .Y(_16448_));
 sky130_vsdinv _47008_ (.A(_16448_),
    .Y(_16449_));
 sky130_fd_sc_hd__nand2_4 _47009_ (.A(_16441_),
    .B(_16449_),
    .Y(_16450_));
 sky130_fd_sc_hd__nand3_4 _47010_ (.A(_16439_),
    .B(_16440_),
    .C(_16448_),
    .Y(_16451_));
 sky130_fd_sc_hd__nand2_4 _47011_ (.A(_16450_),
    .B(_16451_),
    .Y(_16452_));
 sky130_vsdinv _47012_ (.A(_16285_),
    .Y(_16453_));
 sky130_fd_sc_hd__a21oi_4 _47013_ (.A1(_16283_),
    .A2(_16295_),
    .B1(_16453_),
    .Y(_16454_));
 sky130_fd_sc_hd__nand2_4 _47014_ (.A(_16452_),
    .B(_16454_),
    .Y(_16455_));
 sky130_fd_sc_hd__a21o_4 _47015_ (.A1(_16283_),
    .A2(_16295_),
    .B1(_16453_),
    .X(_16456_));
 sky130_fd_sc_hd__nand3_4 _47016_ (.A(_16456_),
    .B(_16450_),
    .C(_16451_),
    .Y(_16457_));
 sky130_fd_sc_hd__nand2_4 _47017_ (.A(_16455_),
    .B(_16457_),
    .Y(_16458_));
 sky130_fd_sc_hd__nand2_4 _47018_ (.A(_16292_),
    .B(_16287_),
    .Y(_16459_));
 sky130_fd_sc_hd__xor2_4 _47019_ (.A(_16148_),
    .B(_16459_),
    .X(_16460_));
 sky130_vsdinv _47020_ (.A(_16460_),
    .Y(_16461_));
 sky130_fd_sc_hd__nand2_4 _47021_ (.A(_16458_),
    .B(_16461_),
    .Y(_16462_));
 sky130_fd_sc_hd__nand3_4 _47022_ (.A(_16455_),
    .B(_16457_),
    .C(_16460_),
    .Y(_16463_));
 sky130_fd_sc_hd__nand2_4 _47023_ (.A(_16462_),
    .B(_16463_),
    .Y(_16464_));
 sky130_fd_sc_hd__a21boi_4 _47024_ (.A1(_16299_),
    .A2(_16304_),
    .B1_N(_16301_),
    .Y(_16465_));
 sky130_fd_sc_hd__nand2_4 _47025_ (.A(_16464_),
    .B(_16465_),
    .Y(_16466_));
 sky130_fd_sc_hd__nand2_4 _47026_ (.A(_16307_),
    .B(_16301_),
    .Y(_16467_));
 sky130_fd_sc_hd__nand3_4 _47027_ (.A(_16467_),
    .B(_16462_),
    .C(_16463_),
    .Y(_16468_));
 sky130_fd_sc_hd__nand2_4 _47028_ (.A(_16466_),
    .B(_16468_),
    .Y(_16469_));
 sky130_fd_sc_hd__a21oi_4 _47029_ (.A1(_16125_),
    .A2(_16121_),
    .B1(_15627_),
    .Y(_16470_));
 sky130_vsdinv _47030_ (.A(_16470_),
    .Y(_16471_));
 sky130_fd_sc_hd__nand2_4 _47031_ (.A(_16469_),
    .B(_16471_),
    .Y(_16472_));
 sky130_fd_sc_hd__nand3_4 _47032_ (.A(_16466_),
    .B(_16468_),
    .C(_16470_),
    .Y(_16473_));
 sky130_fd_sc_hd__nand2_4 _47033_ (.A(_16472_),
    .B(_16473_),
    .Y(_16474_));
 sky130_fd_sc_hd__a21boi_4 _47034_ (.A1(_16311_),
    .A2(_16315_),
    .B1_N(_16312_),
    .Y(_16475_));
 sky130_fd_sc_hd__nand2_4 _47035_ (.A(_16474_),
    .B(_16475_),
    .Y(_16476_));
 sky130_fd_sc_hd__nand2_4 _47036_ (.A(_16318_),
    .B(_16312_),
    .Y(_16477_));
 sky130_fd_sc_hd__nand3_4 _47037_ (.A(_16477_),
    .B(_16473_),
    .C(_16472_),
    .Y(_16478_));
 sky130_fd_sc_hd__and2_4 _47038_ (.A(_16476_),
    .B(_16478_),
    .X(_16479_));
 sky130_fd_sc_hd__buf_1 _47039_ (.A(_16479_),
    .X(_16480_));
 sky130_fd_sc_hd__o21a_4 _47040_ (.A1(_16326_),
    .A2(_16334_),
    .B1(_16323_),
    .X(_16481_));
 sky130_fd_sc_hd__xnor2_4 _47041_ (.A(_16480_),
    .B(_16481_),
    .Y(_01458_));
 sky130_fd_sc_hd__maj3_4 _47042_ (.A(_16379_),
    .B(_16403_),
    .C(_16381_),
    .X(_16482_));
 sky130_vsdinv _47043_ (.A(_16482_),
    .Y(_16483_));
 sky130_fd_sc_hd__nand2_4 _47044_ (.A(_16179_),
    .B(_16335_),
    .Y(_16484_));
 sky130_fd_sc_hd__o21ai_4 _47045_ (.A1(_11915_),
    .A2(_03635_),
    .B1(_16484_),
    .Y(_16485_));
 sky130_fd_sc_hd__nand4_4 _47046_ (.A(_03359_),
    .B(_16179_),
    .C(_16338_),
    .D(_11385_),
    .Y(_16486_));
 sky130_fd_sc_hd__nand2_4 _47047_ (.A(_15863_),
    .B(_03622_),
    .Y(_16487_));
 sky130_vsdinv _47048_ (.A(_16487_),
    .Y(_16488_));
 sky130_fd_sc_hd__a21o_4 _47049_ (.A1(_16485_),
    .A2(_16486_),
    .B1(_16488_),
    .X(_16489_));
 sky130_fd_sc_hd__nand3_4 _47050_ (.A(_16485_),
    .B(_16486_),
    .C(_16488_),
    .Y(_16490_));
 sky130_fd_sc_hd__a21boi_4 _47051_ (.A1(_16337_),
    .A2(_16341_),
    .B1_N(_16339_),
    .Y(_16491_));
 sky130_fd_sc_hd__a21boi_4 _47052_ (.A1(_16489_),
    .A2(_16490_),
    .B1_N(_16491_),
    .Y(_16492_));
 sky130_vsdinv _47053_ (.A(_16492_),
    .Y(_16493_));
 sky130_vsdinv _47054_ (.A(_16491_),
    .Y(_16494_));
 sky130_fd_sc_hd__nand3_4 _47055_ (.A(_16494_),
    .B(_16489_),
    .C(_16490_),
    .Y(_16495_));
 sky130_fd_sc_hd__nand2_4 _47056_ (.A(_12277_),
    .B(_03602_),
    .Y(_16496_));
 sky130_fd_sc_hd__nand2_4 _47057_ (.A(_15864_),
    .B(_15268_),
    .Y(_16497_));
 sky130_fd_sc_hd__nand2_4 _47058_ (.A(_16038_),
    .B(_15267_),
    .Y(_16498_));
 sky130_fd_sc_hd__xnor2_4 _47059_ (.A(_16497_),
    .B(_16498_),
    .Y(_16499_));
 sky130_fd_sc_hd__xor2_4 _47060_ (.A(_16496_),
    .B(_16499_),
    .X(_16500_));
 sky130_fd_sc_hd__a21o_4 _47061_ (.A1(_16493_),
    .A2(_16495_),
    .B1(_16500_),
    .X(_16501_));
 sky130_fd_sc_hd__nand3_4 _47062_ (.A(_16500_),
    .B(_16493_),
    .C(_16495_),
    .Y(_16502_));
 sky130_fd_sc_hd__a21boi_4 _47063_ (.A1(_16346_),
    .A2(_16354_),
    .B1_N(_16347_),
    .Y(_16503_));
 sky130_vsdinv _47064_ (.A(_16503_),
    .Y(_16504_));
 sky130_fd_sc_hd__a21oi_4 _47065_ (.A1(_16501_),
    .A2(_16502_),
    .B1(_16504_),
    .Y(_16505_));
 sky130_fd_sc_hd__nand3_4 _47066_ (.A(_16504_),
    .B(_16501_),
    .C(_16502_),
    .Y(_16506_));
 sky130_vsdinv _47067_ (.A(_16506_),
    .Y(_16507_));
 sky130_fd_sc_hd__a21boi_4 _47068_ (.A1(_16365_),
    .A2(_16368_),
    .B1_N(_16366_),
    .Y(_16508_));
 sky130_vsdinv _47069_ (.A(_16348_),
    .Y(_16509_));
 sky130_fd_sc_hd__nand3_4 _47070_ (.A(_16351_),
    .B(_16352_),
    .C(_16509_),
    .Y(_16510_));
 sky130_fd_sc_hd__nand2_4 _47071_ (.A(_13412_),
    .B(_15499_),
    .Y(_16511_));
 sky130_fd_sc_hd__buf_1 _47072_ (.A(_12114_),
    .X(_16512_));
 sky130_fd_sc_hd__nand2_4 _47073_ (.A(_15136_),
    .B(_16512_),
    .Y(_16513_));
 sky130_fd_sc_hd__nand2_4 _47074_ (.A(_16511_),
    .B(_16513_),
    .Y(_16514_));
 sky130_fd_sc_hd__nand4_4 _47075_ (.A(_13412_),
    .B(_15720_),
    .C(_16512_),
    .D(_15858_),
    .Y(_16515_));
 sky130_fd_sc_hd__nand2_4 _47076_ (.A(_16514_),
    .B(_16515_),
    .Y(_16516_));
 sky130_fd_sc_hd__buf_4 _47077_ (.A(_10847_),
    .X(_16517_));
 sky130_fd_sc_hd__nand2_4 _47078_ (.A(_16517_),
    .B(_03584_),
    .Y(_16518_));
 sky130_fd_sc_hd__nand2_4 _47079_ (.A(_16516_),
    .B(_16518_),
    .Y(_16519_));
 sky130_fd_sc_hd__nand4_4 _47080_ (.A(_16517_),
    .B(_16514_),
    .C(_16515_),
    .D(_03584_),
    .Y(_16520_));
 sky130_fd_sc_hd__nand2_4 _47081_ (.A(_16519_),
    .B(_16520_),
    .Y(_16521_));
 sky130_fd_sc_hd__a21o_4 _47082_ (.A1(_16352_),
    .A2(_16510_),
    .B1(_16521_),
    .X(_16522_));
 sky130_fd_sc_hd__a21boi_4 _47083_ (.A1(_16351_),
    .A2(_16509_),
    .B1_N(_16352_),
    .Y(_16523_));
 sky130_fd_sc_hd__nand2_4 _47084_ (.A(_16521_),
    .B(_16523_),
    .Y(_16524_));
 sky130_fd_sc_hd__nand2_4 _47085_ (.A(_16522_),
    .B(_16524_),
    .Y(_16525_));
 sky130_fd_sc_hd__xor2_4 _47086_ (.A(_16508_),
    .B(_16525_),
    .X(_16526_));
 sky130_vsdinv _47087_ (.A(_16526_),
    .Y(_16527_));
 sky130_fd_sc_hd__o21ai_4 _47088_ (.A1(_16505_),
    .A2(_16507_),
    .B1(_16527_),
    .Y(_16528_));
 sky130_vsdinv _47089_ (.A(_16505_),
    .Y(_16529_));
 sky130_fd_sc_hd__nand3_4 _47090_ (.A(_16529_),
    .B(_16506_),
    .C(_16526_),
    .Y(_16530_));
 sky130_fd_sc_hd__a21boi_4 _47091_ (.A1(_16359_),
    .A2(_16376_),
    .B1_N(_16360_),
    .Y(_16531_));
 sky130_fd_sc_hd__a21boi_4 _47092_ (.A1(_16528_),
    .A2(_16530_),
    .B1_N(_16531_),
    .Y(_16532_));
 sky130_vsdinv _47093_ (.A(_16532_),
    .Y(_16533_));
 sky130_vsdinv _47094_ (.A(_16531_),
    .Y(_16534_));
 sky130_fd_sc_hd__nand3_4 _47095_ (.A(_16534_),
    .B(_16528_),
    .C(_16530_),
    .Y(_16535_));
 sky130_fd_sc_hd__buf_1 _47096_ (.A(_16244_),
    .X(_16536_));
 sky130_fd_sc_hd__a21boi_4 _47097_ (.A1(_16536_),
    .A2(_16393_),
    .B1_N(_16394_),
    .Y(_16537_));
 sky130_vsdinv _47098_ (.A(_16361_),
    .Y(_16538_));
 sky130_fd_sc_hd__nand3_4 _47099_ (.A(_16373_),
    .B(_16538_),
    .C(_16374_),
    .Y(_16539_));
 sky130_fd_sc_hd__buf_1 _47100_ (.A(_12910_),
    .X(_16540_));
 sky130_fd_sc_hd__nand2_4 _47101_ (.A(_16540_),
    .B(_03572_),
    .Y(_16541_));
 sky130_fd_sc_hd__o21ai_4 _47102_ (.A1(_03401_),
    .A2(_03578_),
    .B1(_16541_),
    .Y(_16542_));
 sky130_fd_sc_hd__buf_1 _47103_ (.A(_15899_),
    .X(_16543_));
 sky130_fd_sc_hd__buf_1 _47104_ (.A(_14377_),
    .X(_16544_));
 sky130_fd_sc_hd__nand4_4 _47105_ (.A(_16543_),
    .B(_16540_),
    .C(_03572_),
    .D(_16544_),
    .Y(_16545_));
 sky130_fd_sc_hd__buf_1 _47106_ (.A(_16388_),
    .X(_16546_));
 sky130_fd_sc_hd__a21o_4 _47107_ (.A1(_16542_),
    .A2(_16545_),
    .B1(_16546_),
    .X(_16547_));
 sky130_fd_sc_hd__nand3_4 _47108_ (.A(_16542_),
    .B(_16545_),
    .C(_16546_),
    .Y(_16548_));
 sky130_fd_sc_hd__a21boi_4 _47109_ (.A1(_16385_),
    .A2(_16546_),
    .B1_N(_16386_),
    .Y(_16549_));
 sky130_vsdinv _47110_ (.A(_16549_),
    .Y(_16550_));
 sky130_fd_sc_hd__a21o_4 _47111_ (.A1(_16547_),
    .A2(_16548_),
    .B1(_16550_),
    .X(_16551_));
 sky130_fd_sc_hd__nand3_4 _47112_ (.A(_16547_),
    .B(_16550_),
    .C(_16548_),
    .Y(_16552_));
 sky130_fd_sc_hd__a21o_4 _47113_ (.A1(_16551_),
    .A2(_16552_),
    .B1(_16244_),
    .X(_16553_));
 sky130_fd_sc_hd__nand3_4 _47114_ (.A(_16551_),
    .B(_16536_),
    .C(_16552_),
    .Y(_16554_));
 sky130_fd_sc_hd__nand2_4 _47115_ (.A(_16553_),
    .B(_16554_),
    .Y(_16555_));
 sky130_fd_sc_hd__a21o_4 _47116_ (.A1(_16373_),
    .A2(_16539_),
    .B1(_16555_),
    .X(_16556_));
 sky130_fd_sc_hd__nand3_4 _47117_ (.A(_16555_),
    .B(_16373_),
    .C(_16539_),
    .Y(_16557_));
 sky130_fd_sc_hd__nand2_4 _47118_ (.A(_16556_),
    .B(_16557_),
    .Y(_16558_));
 sky130_fd_sc_hd__xor2_4 _47119_ (.A(_16537_),
    .B(_16558_),
    .X(_16559_));
 sky130_fd_sc_hd__a21o_4 _47120_ (.A1(_16533_),
    .A2(_16535_),
    .B1(_16559_),
    .X(_16560_));
 sky130_fd_sc_hd__nand3_4 _47121_ (.A(_16533_),
    .B(_16535_),
    .C(_16559_),
    .Y(_16561_));
 sky130_fd_sc_hd__nand3_4 _47122_ (.A(_16483_),
    .B(_16560_),
    .C(_16561_),
    .Y(_16562_));
 sky130_fd_sc_hd__nand2_4 _47123_ (.A(_16560_),
    .B(_16561_),
    .Y(_16563_));
 sky130_fd_sc_hd__nand2_4 _47124_ (.A(_16563_),
    .B(_16482_),
    .Y(_16564_));
 sky130_fd_sc_hd__or4_4 _47125_ (.A(_15358_),
    .B(_15549_),
    .C(_15744_),
    .D(_16413_),
    .X(_16565_));
 sky130_fd_sc_hd__buf_1 _47126_ (.A(_16565_),
    .X(_16566_));
 sky130_fd_sc_hd__nand4_4 _47127_ (.A(_15358_),
    .B(_16413_),
    .C(_15549_),
    .D(_15744_),
    .Y(_16567_));
 sky130_fd_sc_hd__nand2_4 _47128_ (.A(_16566_),
    .B(_16567_),
    .Y(_16568_));
 sky130_fd_sc_hd__xor2_4 _47129_ (.A(_16568_),
    .B(_15762_),
    .X(_16569_));
 sky130_fd_sc_hd__buf_1 _47130_ (.A(_16569_),
    .X(_16570_));
 sky130_fd_sc_hd__a21o_4 _47131_ (.A1(_16401_),
    .A2(_16398_),
    .B1(_16570_),
    .X(_16571_));
 sky130_fd_sc_hd__nand3_4 _47132_ (.A(_16401_),
    .B(_16398_),
    .C(_16570_),
    .Y(_16572_));
 sky130_fd_sc_hd__nand2_4 _47133_ (.A(_16422_),
    .B(_16566_),
    .Y(_16573_));
 sky130_fd_sc_hd__a21o_4 _47134_ (.A1(_16571_),
    .A2(_16572_),
    .B1(_16573_),
    .X(_16574_));
 sky130_fd_sc_hd__nand3_4 _47135_ (.A(_16571_),
    .B(_16572_),
    .C(_16573_),
    .Y(_16575_));
 sky130_fd_sc_hd__and2_4 _47136_ (.A(_16574_),
    .B(_16575_),
    .X(_16576_));
 sky130_fd_sc_hd__a21o_4 _47137_ (.A1(_16562_),
    .A2(_16564_),
    .B1(_16576_),
    .X(_16577_));
 sky130_fd_sc_hd__nand3_4 _47138_ (.A(_16562_),
    .B(_16564_),
    .C(_16576_),
    .Y(_16578_));
 sky130_fd_sc_hd__nand2_4 _47139_ (.A(_16577_),
    .B(_16578_),
    .Y(_16579_));
 sky130_vsdinv _47140_ (.A(_16411_),
    .Y(_16580_));
 sky130_fd_sc_hd__a21oi_4 _47141_ (.A1(_16409_),
    .A2(_16432_),
    .B1(_16580_),
    .Y(_16581_));
 sky130_fd_sc_hd__nand2_4 _47142_ (.A(_16579_),
    .B(_16581_),
    .Y(_16582_));
 sky130_vsdinv _47143_ (.A(_16581_),
    .Y(_16583_));
 sky130_fd_sc_hd__nand3_4 _47144_ (.A(_16583_),
    .B(_16577_),
    .C(_16578_),
    .Y(_16584_));
 sky130_fd_sc_hd__nand2_4 _47145_ (.A(_16582_),
    .B(_16584_),
    .Y(_16585_));
 sky130_fd_sc_hd__a21o_4 _47146_ (.A1(_16430_),
    .A2(_16426_),
    .B1(_16288_),
    .X(_16586_));
 sky130_fd_sc_hd__buf_1 _47147_ (.A(_16288_),
    .X(_16587_));
 sky130_fd_sc_hd__nand3_4 _47148_ (.A(_16430_),
    .B(_16587_),
    .C(_16426_),
    .Y(_16588_));
 sky130_fd_sc_hd__a21o_4 _47149_ (.A1(_16586_),
    .A2(_16588_),
    .B1(_16444_),
    .X(_16589_));
 sky130_fd_sc_hd__nand3_4 _47150_ (.A(_16586_),
    .B(_16444_),
    .C(_16588_),
    .Y(_16590_));
 sky130_fd_sc_hd__nand2_4 _47151_ (.A(_16589_),
    .B(_16590_),
    .Y(_16591_));
 sky130_fd_sc_hd__nand2_4 _47152_ (.A(_16585_),
    .B(_16591_),
    .Y(_16592_));
 sky130_fd_sc_hd__nand4_4 _47153_ (.A(_16584_),
    .B(_16582_),
    .C(_16590_),
    .D(_16589_),
    .Y(_16593_));
 sky130_fd_sc_hd__nand2_4 _47154_ (.A(_16592_),
    .B(_16593_),
    .Y(_16594_));
 sky130_fd_sc_hd__a21boi_4 _47155_ (.A1(_16439_),
    .A2(_16448_),
    .B1_N(_16440_),
    .Y(_16595_));
 sky130_fd_sc_hd__nand2_4 _47156_ (.A(_16594_),
    .B(_16595_),
    .Y(_16596_));
 sky130_vsdinv _47157_ (.A(_16595_),
    .Y(_16597_));
 sky130_fd_sc_hd__nand3_4 _47158_ (.A(_16597_),
    .B(_16592_),
    .C(_16593_),
    .Y(_16598_));
 sky130_fd_sc_hd__nand2_4 _47159_ (.A(_16596_),
    .B(_16598_),
    .Y(_16599_));
 sky130_fd_sc_hd__nand2_4 _47160_ (.A(_16446_),
    .B(_16442_),
    .Y(_16600_));
 sky130_fd_sc_hd__xor2_4 _47161_ (.A(_16148_),
    .B(_16600_),
    .X(_16601_));
 sky130_vsdinv _47162_ (.A(_16601_),
    .Y(_16602_));
 sky130_fd_sc_hd__nand2_4 _47163_ (.A(_16599_),
    .B(_16602_),
    .Y(_16603_));
 sky130_fd_sc_hd__nand3_4 _47164_ (.A(_16596_),
    .B(_16598_),
    .C(_16601_),
    .Y(_16604_));
 sky130_fd_sc_hd__nand2_4 _47165_ (.A(_16603_),
    .B(_16604_),
    .Y(_16605_));
 sky130_fd_sc_hd__nand2_4 _47166_ (.A(_16463_),
    .B(_16457_),
    .Y(_16606_));
 sky130_vsdinv _47167_ (.A(_16606_),
    .Y(_16607_));
 sky130_fd_sc_hd__nand2_4 _47168_ (.A(_16605_),
    .B(_16607_),
    .Y(_16608_));
 sky130_fd_sc_hd__nand3_4 _47169_ (.A(_16606_),
    .B(_16603_),
    .C(_16604_),
    .Y(_16609_));
 sky130_fd_sc_hd__nand2_4 _47170_ (.A(_16608_),
    .B(_16609_),
    .Y(_16610_));
 sky130_fd_sc_hd__a21oi_4 _47171_ (.A1(_16292_),
    .A2(_16287_),
    .B1(_15627_),
    .Y(_16611_));
 sky130_vsdinv _47172_ (.A(_16611_),
    .Y(_16612_));
 sky130_fd_sc_hd__nand2_4 _47173_ (.A(_16610_),
    .B(_16612_),
    .Y(_16613_));
 sky130_fd_sc_hd__nand3_4 _47174_ (.A(_16608_),
    .B(_16611_),
    .C(_16609_),
    .Y(_16614_));
 sky130_fd_sc_hd__nand2_4 _47175_ (.A(_16473_),
    .B(_16468_),
    .Y(_16615_));
 sky130_fd_sc_hd__a21oi_4 _47176_ (.A1(_16613_),
    .A2(_16614_),
    .B1(_16615_),
    .Y(_16616_));
 sky130_fd_sc_hd__nand3_4 _47177_ (.A(_16615_),
    .B(_16613_),
    .C(_16614_),
    .Y(_16617_));
 sky130_vsdinv _47178_ (.A(_16617_),
    .Y(_16618_));
 sky130_fd_sc_hd__nor2_4 _47179_ (.A(_16616_),
    .B(_16618_),
    .Y(_16619_));
 sky130_fd_sc_hd__nand4_4 _47180_ (.A(_16323_),
    .B(_16322_),
    .C(_16476_),
    .D(_16478_),
    .Y(_16620_));
 sky130_fd_sc_hd__nand2_4 _47181_ (.A(_16478_),
    .B(_16323_),
    .Y(_16621_));
 sky130_fd_sc_hd__nand2_4 _47182_ (.A(_16621_),
    .B(_16476_),
    .Y(_16622_));
 sky130_fd_sc_hd__o21ai_4 _47183_ (.A1(_16620_),
    .A2(_16334_),
    .B1(_16622_),
    .Y(_16623_));
 sky130_fd_sc_hd__xor2_4 _47184_ (.A(_16619_),
    .B(_16623_),
    .X(_01459_));
 sky130_fd_sc_hd__buf_4 _47185_ (.A(_15659_),
    .X(_16624_));
 sky130_fd_sc_hd__nand2_4 _47186_ (.A(_16180_),
    .B(_16624_),
    .Y(_16625_));
 sky130_fd_sc_hd__o21ai_4 _47187_ (.A1(_16179_),
    .A2(_03635_),
    .B1(_16625_),
    .Y(_16626_));
 sky130_fd_sc_hd__nand4_4 _47188_ (.A(_03362_),
    .B(_16180_),
    .C(_16624_),
    .D(_11386_),
    .Y(_16627_));
 sky130_fd_sc_hd__nand2_4 _47189_ (.A(_16037_),
    .B(_03622_),
    .Y(_16628_));
 sky130_vsdinv _47190_ (.A(_16628_),
    .Y(_16629_));
 sky130_fd_sc_hd__a21o_4 _47191_ (.A1(_16626_),
    .A2(_16627_),
    .B1(_16629_),
    .X(_16630_));
 sky130_fd_sc_hd__nand3_4 _47192_ (.A(_16626_),
    .B(_16627_),
    .C(_16629_),
    .Y(_16631_));
 sky130_fd_sc_hd__a21boi_4 _47193_ (.A1(_16485_),
    .A2(_16488_),
    .B1_N(_16486_),
    .Y(_16632_));
 sky130_vsdinv _47194_ (.A(_16632_),
    .Y(_16633_));
 sky130_fd_sc_hd__a21o_4 _47195_ (.A1(_16630_),
    .A2(_16631_),
    .B1(_16633_),
    .X(_16634_));
 sky130_fd_sc_hd__nand3_4 _47196_ (.A(_16633_),
    .B(_16630_),
    .C(_16631_),
    .Y(_16635_));
 sky130_fd_sc_hd__nand2_4 _47197_ (.A(_15885_),
    .B(_03601_),
    .Y(_16636_));
 sky130_fd_sc_hd__nand2_4 _47198_ (.A(_11954_),
    .B(_15263_),
    .Y(_16637_));
 sky130_fd_sc_hd__nand2_4 _47199_ (.A(_11955_),
    .B(_03607_),
    .Y(_16638_));
 sky130_fd_sc_hd__xnor2_4 _47200_ (.A(_16637_),
    .B(_16638_),
    .Y(_16639_));
 sky130_fd_sc_hd__xor2_4 _47201_ (.A(_16636_),
    .B(_16639_),
    .X(_16640_));
 sky130_fd_sc_hd__a21o_4 _47202_ (.A1(_16634_),
    .A2(_16635_),
    .B1(_16640_),
    .X(_16641_));
 sky130_fd_sc_hd__nand3_4 _47203_ (.A(_16640_),
    .B(_16634_),
    .C(_16635_),
    .Y(_16642_));
 sky130_vsdinv _47204_ (.A(_16495_),
    .Y(_16643_));
 sky130_fd_sc_hd__a21oi_4 _47205_ (.A1(_16500_),
    .A2(_16493_),
    .B1(_16643_),
    .Y(_16644_));
 sky130_vsdinv _47206_ (.A(_16644_),
    .Y(_16645_));
 sky130_fd_sc_hd__a21o_4 _47207_ (.A1(_16641_),
    .A2(_16642_),
    .B1(_16645_),
    .X(_16646_));
 sky130_fd_sc_hd__nand3_4 _47208_ (.A(_16645_),
    .B(_16641_),
    .C(_16642_),
    .Y(_16647_));
 sky130_fd_sc_hd__maj3_4 _47209_ (.A(_16497_),
    .B(_16498_),
    .C(_16496_),
    .X(_16648_));
 sky130_vsdinv _47210_ (.A(_12721_),
    .Y(_16649_));
 sky130_fd_sc_hd__a2bb2o_4 _47211_ (.A1_N(_03398_),
    .A2_N(_16649_),
    .B1(_15720_),
    .B2(_15858_),
    .X(_16650_));
 sky130_fd_sc_hd__nand4_4 _47212_ (.A(_15720_),
    .B(_13410_),
    .C(_16512_),
    .D(_15499_),
    .Y(_16651_));
 sky130_fd_sc_hd__nand2_4 _47213_ (.A(_14204_),
    .B(_16195_),
    .Y(_16652_));
 sky130_vsdinv _47214_ (.A(_16652_),
    .Y(_16653_));
 sky130_fd_sc_hd__a21o_4 _47215_ (.A1(_16650_),
    .A2(_16651_),
    .B1(_16653_),
    .X(_16654_));
 sky130_fd_sc_hd__nand3_4 _47216_ (.A(_16650_),
    .B(_16651_),
    .C(_16653_),
    .Y(_16655_));
 sky130_fd_sc_hd__nand2_4 _47217_ (.A(_16654_),
    .B(_16655_),
    .Y(_16656_));
 sky130_fd_sc_hd__or2_4 _47218_ (.A(_16648_),
    .B(_16656_),
    .X(_16657_));
 sky130_fd_sc_hd__buf_1 _47219_ (.A(_16657_),
    .X(_16658_));
 sky130_fd_sc_hd__nand2_4 _47220_ (.A(_16656_),
    .B(_16648_),
    .Y(_16659_));
 sky130_fd_sc_hd__nand2_4 _47221_ (.A(_16520_),
    .B(_16515_),
    .Y(_16660_));
 sky130_fd_sc_hd__a21oi_4 _47222_ (.A1(_16658_),
    .A2(_16659_),
    .B1(_16660_),
    .Y(_16661_));
 sky130_fd_sc_hd__nand3_4 _47223_ (.A(_16658_),
    .B(_16660_),
    .C(_16659_),
    .Y(_16662_));
 sky130_vsdinv _47224_ (.A(_16662_),
    .Y(_16663_));
 sky130_fd_sc_hd__nor2_4 _47225_ (.A(_16661_),
    .B(_16663_),
    .Y(_16664_));
 sky130_fd_sc_hd__a21o_4 _47226_ (.A1(_16646_),
    .A2(_16647_),
    .B1(_16664_),
    .X(_16665_));
 sky130_fd_sc_hd__nand3_4 _47227_ (.A(_16664_),
    .B(_16646_),
    .C(_16647_),
    .Y(_16666_));
 sky130_fd_sc_hd__o21a_4 _47228_ (.A1(_16505_),
    .A2(_16527_),
    .B1(_16506_),
    .X(_16667_));
 sky130_vsdinv _47229_ (.A(_16667_),
    .Y(_16668_));
 sky130_fd_sc_hd__a21o_4 _47230_ (.A1(_16665_),
    .A2(_16666_),
    .B1(_16668_),
    .X(_16669_));
 sky130_fd_sc_hd__nand3_4 _47231_ (.A(_16668_),
    .B(_16665_),
    .C(_16666_),
    .Y(_16670_));
 sky130_fd_sc_hd__a21boi_4 _47232_ (.A1(_16551_),
    .A2(_16536_),
    .B1_N(_16552_),
    .Y(_16671_));
 sky130_fd_sc_hd__o21a_4 _47233_ (.A1(_03571_),
    .A2(_16544_),
    .B1(_03408_),
    .X(_16672_));
 sky130_fd_sc_hd__nand3_4 _47234_ (.A(_03409_),
    .B(_03572_),
    .C(_16544_),
    .Y(_16673_));
 sky130_fd_sc_hd__a21o_4 _47235_ (.A1(_16672_),
    .A2(_16673_),
    .B1(_16387_),
    .X(_16674_));
 sky130_fd_sc_hd__nand3_4 _47236_ (.A(_16672_),
    .B(_16387_),
    .C(_16673_),
    .Y(_16675_));
 sky130_fd_sc_hd__a21boi_4 _47237_ (.A1(_16542_),
    .A2(_16546_),
    .B1_N(_16545_),
    .Y(_16676_));
 sky130_vsdinv _47238_ (.A(_16676_),
    .Y(_16677_));
 sky130_fd_sc_hd__a21o_4 _47239_ (.A1(_16674_),
    .A2(_16675_),
    .B1(_16677_),
    .X(_16678_));
 sky130_fd_sc_hd__nand3_4 _47240_ (.A(_16677_),
    .B(_16674_),
    .C(_16675_),
    .Y(_16679_));
 sky130_vsdinv _47241_ (.A(_16244_),
    .Y(_16680_));
 sky130_fd_sc_hd__a21o_4 _47242_ (.A1(_16678_),
    .A2(_16679_),
    .B1(_16680_),
    .X(_16681_));
 sky130_fd_sc_hd__nand3_4 _47243_ (.A(_16680_),
    .B(_16678_),
    .C(_16679_),
    .Y(_16682_));
 sky130_fd_sc_hd__maj3_4 _47244_ (.A(_16508_),
    .B(_16521_),
    .C(_16523_),
    .X(_16683_));
 sky130_vsdinv _47245_ (.A(_16683_),
    .Y(_16684_));
 sky130_fd_sc_hd__a21o_4 _47246_ (.A1(_16681_),
    .A2(_16682_),
    .B1(_16684_),
    .X(_16685_));
 sky130_fd_sc_hd__nand3_4 _47247_ (.A(_16681_),
    .B(_16684_),
    .C(_16682_),
    .Y(_16686_));
 sky130_fd_sc_hd__nand2_4 _47248_ (.A(_16685_),
    .B(_16686_),
    .Y(_16687_));
 sky130_fd_sc_hd__xor2_4 _47249_ (.A(_16671_),
    .B(_16687_),
    .X(_16688_));
 sky130_fd_sc_hd__a21o_4 _47250_ (.A1(_16669_),
    .A2(_16670_),
    .B1(_16688_),
    .X(_16689_));
 sky130_fd_sc_hd__nand3_4 _47251_ (.A(_16669_),
    .B(_16670_),
    .C(_16688_),
    .Y(_16690_));
 sky130_fd_sc_hd__nand2_4 _47252_ (.A(_16689_),
    .B(_16690_),
    .Y(_16691_));
 sky130_fd_sc_hd__a21boi_4 _47253_ (.A1(_16533_),
    .A2(_16559_),
    .B1_N(_16535_),
    .Y(_16692_));
 sky130_fd_sc_hd__nand2_4 _47254_ (.A(_16691_),
    .B(_16692_),
    .Y(_16693_));
 sky130_vsdinv _47255_ (.A(_16692_),
    .Y(_16694_));
 sky130_fd_sc_hd__nand3_4 _47256_ (.A(_16694_),
    .B(_16689_),
    .C(_16690_),
    .Y(_16695_));
 sky130_fd_sc_hd__a21boi_4 _47257_ (.A1(_16266_),
    .A2(_16567_),
    .B1_N(_16566_),
    .Y(_16696_));
 sky130_fd_sc_hd__buf_8 _47258_ (.A(_16696_),
    .X(_16697_));
 sky130_fd_sc_hd__maj3_4 _47259_ (.A(_16361_),
    .B(_16371_),
    .C(_16362_),
    .X(_16698_));
 sky130_fd_sc_hd__maj3_4 _47260_ (.A(_16537_),
    .B(_16555_),
    .C(_16698_),
    .X(_16699_));
 sky130_fd_sc_hd__or2_4 _47261_ (.A(_16570_),
    .B(_16699_),
    .X(_16700_));
 sky130_fd_sc_hd__buf_1 _47262_ (.A(_16569_),
    .X(_16701_));
 sky130_fd_sc_hd__nand2_4 _47263_ (.A(_16699_),
    .B(_16701_),
    .Y(_16702_));
 sky130_fd_sc_hd__nand2_4 _47264_ (.A(_16700_),
    .B(_16702_),
    .Y(_16703_));
 sky130_fd_sc_hd__xor2_4 _47265_ (.A(_16697_),
    .B(_16703_),
    .X(_16704_));
 sky130_fd_sc_hd__a21o_4 _47266_ (.A1(_16693_),
    .A2(_16695_),
    .B1(_16704_),
    .X(_16705_));
 sky130_fd_sc_hd__nand3_4 _47267_ (.A(_16693_),
    .B(_16695_),
    .C(_16704_),
    .Y(_16706_));
 sky130_fd_sc_hd__nand2_4 _47268_ (.A(_16578_),
    .B(_16562_),
    .Y(_16707_));
 sky130_fd_sc_hd__a21oi_4 _47269_ (.A1(_16705_),
    .A2(_16706_),
    .B1(_16707_),
    .Y(_16708_));
 sky130_fd_sc_hd__nand3_4 _47270_ (.A(_16707_),
    .B(_16705_),
    .C(_16706_),
    .Y(_16709_));
 sky130_vsdinv _47271_ (.A(_16709_),
    .Y(_16710_));
 sky130_fd_sc_hd__a21o_4 _47272_ (.A1(_16575_),
    .A2(_16571_),
    .B1(_15962_),
    .X(_16711_));
 sky130_fd_sc_hd__nand3_4 _47273_ (.A(_16575_),
    .B(_16288_),
    .C(_16571_),
    .Y(_16712_));
 sky130_fd_sc_hd__a21o_4 _47274_ (.A1(_16711_),
    .A2(_16712_),
    .B1(_16290_),
    .X(_16713_));
 sky130_fd_sc_hd__nand3_4 _47275_ (.A(_16711_),
    .B(_16290_),
    .C(_16712_),
    .Y(_16714_));
 sky130_fd_sc_hd__and2_4 _47276_ (.A(_16713_),
    .B(_16714_),
    .X(_16715_));
 sky130_vsdinv _47277_ (.A(_16715_),
    .Y(_16716_));
 sky130_fd_sc_hd__o21ai_4 _47278_ (.A1(_16708_),
    .A2(_16710_),
    .B1(_16716_),
    .Y(_16717_));
 sky130_vsdinv _47279_ (.A(_16708_),
    .Y(_16718_));
 sky130_fd_sc_hd__nand3_4 _47280_ (.A(_16718_),
    .B(_16709_),
    .C(_16715_),
    .Y(_16719_));
 sky130_fd_sc_hd__nand2_4 _47281_ (.A(_16717_),
    .B(_16719_),
    .Y(_16720_));
 sky130_fd_sc_hd__a21boi_4 _47282_ (.A1(_16577_),
    .A2(_16578_),
    .B1_N(_16581_),
    .Y(_16721_));
 sky130_fd_sc_hd__o21ai_4 _47283_ (.A1(_16591_),
    .A2(_16721_),
    .B1(_16584_),
    .Y(_16722_));
 sky130_vsdinv _47284_ (.A(_16722_),
    .Y(_16723_));
 sky130_fd_sc_hd__nand2_4 _47285_ (.A(_16720_),
    .B(_16723_),
    .Y(_16724_));
 sky130_fd_sc_hd__nand3_4 _47286_ (.A(_16722_),
    .B(_16717_),
    .C(_16719_),
    .Y(_16725_));
 sky130_fd_sc_hd__nand2_4 _47287_ (.A(_16724_),
    .B(_16725_),
    .Y(_16726_));
 sky130_fd_sc_hd__nand2_4 _47288_ (.A(_16590_),
    .B(_16586_),
    .Y(_16727_));
 sky130_fd_sc_hd__xor2_4 _47289_ (.A(_16148_),
    .B(_16727_),
    .X(_16728_));
 sky130_vsdinv _47290_ (.A(_16728_),
    .Y(_16729_));
 sky130_fd_sc_hd__nand2_4 _47291_ (.A(_16726_),
    .B(_16729_),
    .Y(_16730_));
 sky130_fd_sc_hd__nand3_4 _47292_ (.A(_16724_),
    .B(_16725_),
    .C(_16728_),
    .Y(_16731_));
 sky130_fd_sc_hd__nand2_4 _47293_ (.A(_16730_),
    .B(_16731_),
    .Y(_16732_));
 sky130_fd_sc_hd__a21boi_4 _47294_ (.A1(_16596_),
    .A2(_16601_),
    .B1_N(_16598_),
    .Y(_16733_));
 sky130_fd_sc_hd__nand2_4 _47295_ (.A(_16732_),
    .B(_16733_),
    .Y(_16734_));
 sky130_fd_sc_hd__nand2_4 _47296_ (.A(_16604_),
    .B(_16598_),
    .Y(_16735_));
 sky130_fd_sc_hd__nand3_4 _47297_ (.A(_16735_),
    .B(_16731_),
    .C(_16730_),
    .Y(_16736_));
 sky130_fd_sc_hd__nand2_4 _47298_ (.A(_16734_),
    .B(_16736_),
    .Y(_16737_));
 sky130_fd_sc_hd__a21oi_4 _47299_ (.A1(_16446_),
    .A2(_16442_),
    .B1(_16314_),
    .Y(_16738_));
 sky130_vsdinv _47300_ (.A(_16738_),
    .Y(_16739_));
 sky130_fd_sc_hd__nand2_4 _47301_ (.A(_16737_),
    .B(_16739_),
    .Y(_16740_));
 sky130_fd_sc_hd__nand3_4 _47302_ (.A(_16734_),
    .B(_16738_),
    .C(_16736_),
    .Y(_16741_));
 sky130_fd_sc_hd__a21oi_4 _47303_ (.A1(_16603_),
    .A2(_16604_),
    .B1(_16606_),
    .Y(_16742_));
 sky130_fd_sc_hd__o21ai_4 _47304_ (.A1(_16612_),
    .A2(_16742_),
    .B1(_16609_),
    .Y(_16743_));
 sky130_fd_sc_hd__a21oi_4 _47305_ (.A1(_16740_),
    .A2(_16741_),
    .B1(_16743_),
    .Y(_16744_));
 sky130_fd_sc_hd__nand3_4 _47306_ (.A(_16740_),
    .B(_16743_),
    .C(_16741_),
    .Y(_16745_));
 sky130_vsdinv _47307_ (.A(_16745_),
    .Y(_16746_));
 sky130_fd_sc_hd__nor2_4 _47308_ (.A(_16744_),
    .B(_16746_),
    .Y(_16747_));
 sky130_fd_sc_hd__nand2_4 _47309_ (.A(_16613_),
    .B(_16614_),
    .Y(_16748_));
 sky130_vsdinv _47310_ (.A(_16615_),
    .Y(_16749_));
 sky130_fd_sc_hd__nand2_4 _47311_ (.A(_16748_),
    .B(_16749_),
    .Y(_16750_));
 sky130_fd_sc_hd__a21oi_4 _47312_ (.A1(_16623_),
    .A2(_16750_),
    .B1(_16618_),
    .Y(_16751_));
 sky130_fd_sc_hd__xnor2_4 _47313_ (.A(_16747_),
    .B(_16751_),
    .Y(_01460_));
 sky130_fd_sc_hd__buf_1 _47314_ (.A(_14884_),
    .X(_16752_));
 sky130_fd_sc_hd__nand2_4 _47315_ (.A(_16752_),
    .B(_03622_),
    .Y(_16753_));
 sky130_fd_sc_hd__a2bb2o_4 _47316_ (.A1_N(_15863_),
    .A2_N(_15249_),
    .B1(_15864_),
    .B2(_16335_),
    .X(_16754_));
 sky130_fd_sc_hd__nand4_4 _47317_ (.A(_03366_),
    .B(_15864_),
    .C(_16335_),
    .D(_11385_),
    .Y(_16755_));
 sky130_fd_sc_hd__and2_4 _47318_ (.A(_16754_),
    .B(_16755_),
    .X(_16756_));
 sky130_fd_sc_hd__xor2_4 _47319_ (.A(_16753_),
    .B(_16756_),
    .X(_16757_));
 sky130_fd_sc_hd__a21o_4 _47320_ (.A1(_16627_),
    .A2(_16631_),
    .B1(_16757_),
    .X(_16758_));
 sky130_fd_sc_hd__nand3_4 _47321_ (.A(_16757_),
    .B(_16627_),
    .C(_16631_),
    .Y(_16759_));
 sky130_fd_sc_hd__nand2_4 _47322_ (.A(_10844_),
    .B(_03602_),
    .Y(_16760_));
 sky130_fd_sc_hd__nand2_4 _47323_ (.A(_16040_),
    .B(_03615_),
    .Y(_16761_));
 sky130_fd_sc_hd__buf_1 _47324_ (.A(_15885_),
    .X(_16762_));
 sky130_fd_sc_hd__nand2_4 _47325_ (.A(_16762_),
    .B(_03608_),
    .Y(_16763_));
 sky130_fd_sc_hd__xnor2_4 _47326_ (.A(_16761_),
    .B(_16763_),
    .Y(_16764_));
 sky130_fd_sc_hd__xor2_4 _47327_ (.A(_16760_),
    .B(_16764_),
    .X(_16765_));
 sky130_fd_sc_hd__a21o_4 _47328_ (.A1(_16758_),
    .A2(_16759_),
    .B1(_16765_),
    .X(_16766_));
 sky130_fd_sc_hd__nand3_4 _47329_ (.A(_16758_),
    .B(_16759_),
    .C(_16765_),
    .Y(_16767_));
 sky130_fd_sc_hd__a21boi_4 _47330_ (.A1(_16640_),
    .A2(_16634_),
    .B1_N(_16635_),
    .Y(_16768_));
 sky130_vsdinv _47331_ (.A(_16768_),
    .Y(_16769_));
 sky130_fd_sc_hd__a21oi_4 _47332_ (.A1(_16766_),
    .A2(_16767_),
    .B1(_16769_),
    .Y(_16770_));
 sky130_fd_sc_hd__nand3_4 _47333_ (.A(_16766_),
    .B(_16767_),
    .C(_16769_),
    .Y(_16771_));
 sky130_vsdinv _47334_ (.A(_16771_),
    .Y(_16772_));
 sky130_fd_sc_hd__a2bb2o_4 _47335_ (.A1_N(_03401_),
    .A2_N(_16649_),
    .B1(_15897_),
    .B2(_03598_),
    .X(_16773_));
 sky130_fd_sc_hd__nand4_4 _47336_ (.A(_15897_),
    .B(_10838_),
    .C(_03589_),
    .D(_15865_),
    .Y(_16774_));
 sky130_fd_sc_hd__nand2_4 _47337_ (.A(_03407_),
    .B(_16195_),
    .Y(_16775_));
 sky130_vsdinv _47338_ (.A(_16775_),
    .Y(_16776_));
 sky130_fd_sc_hd__buf_1 _47339_ (.A(_16776_),
    .X(_16777_));
 sky130_fd_sc_hd__a21o_4 _47340_ (.A1(_16773_),
    .A2(_16774_),
    .B1(_16777_),
    .X(_16778_));
 sky130_fd_sc_hd__nand3_4 _47341_ (.A(_16773_),
    .B(_16774_),
    .C(_16776_),
    .Y(_16779_));
 sky130_fd_sc_hd__maj3_4 _47342_ (.A(_16637_),
    .B(_16638_),
    .C(_16636_),
    .X(_16780_));
 sky130_vsdinv _47343_ (.A(_16780_),
    .Y(_16781_));
 sky130_fd_sc_hd__a21o_4 _47344_ (.A1(_16778_),
    .A2(_16779_),
    .B1(_16781_),
    .X(_16782_));
 sky130_fd_sc_hd__nand3_4 _47345_ (.A(_16778_),
    .B(_16781_),
    .C(_16779_),
    .Y(_16783_));
 sky130_fd_sc_hd__nand2_4 _47346_ (.A(_16782_),
    .B(_16783_),
    .Y(_16784_));
 sky130_fd_sc_hd__a21o_4 _47347_ (.A1(_16651_),
    .A2(_16655_),
    .B1(_16784_),
    .X(_16785_));
 sky130_fd_sc_hd__nand3_4 _47348_ (.A(_16784_),
    .B(_16651_),
    .C(_16655_),
    .Y(_16786_));
 sky130_fd_sc_hd__and2_4 _47349_ (.A(_16785_),
    .B(_16786_),
    .X(_16787_));
 sky130_vsdinv _47350_ (.A(_16787_),
    .Y(_16788_));
 sky130_fd_sc_hd__o21ai_4 _47351_ (.A1(_16770_),
    .A2(_16772_),
    .B1(_16788_),
    .Y(_16789_));
 sky130_vsdinv _47352_ (.A(_16770_),
    .Y(_16790_));
 sky130_fd_sc_hd__nand3_4 _47353_ (.A(_16790_),
    .B(_16771_),
    .C(_16787_),
    .Y(_16791_));
 sky130_fd_sc_hd__a21boi_4 _47354_ (.A1(_16664_),
    .A2(_16646_),
    .B1_N(_16647_),
    .Y(_16792_));
 sky130_vsdinv _47355_ (.A(_16792_),
    .Y(_16793_));
 sky130_fd_sc_hd__a21o_4 _47356_ (.A1(_16789_),
    .A2(_16791_),
    .B1(_16793_),
    .X(_16794_));
 sky130_fd_sc_hd__nand3_4 _47357_ (.A(_16789_),
    .B(_16791_),
    .C(_16793_),
    .Y(_16795_));
 sky130_fd_sc_hd__nand4_4 _47358_ (.A(_16540_),
    .B(_03565_),
    .C(_03571_),
    .D(_16544_),
    .Y(_16796_));
 sky130_fd_sc_hd__nand2_4 _47359_ (.A(_16681_),
    .B(_16796_),
    .Y(_16797_));
 sky130_fd_sc_hd__o21a_4 _47360_ (.A1(_16388_),
    .A2(_16672_),
    .B1(_16796_),
    .X(_16798_));
 sky130_fd_sc_hd__xor2_4 _47361_ (.A(_16798_),
    .B(_16241_),
    .X(_16799_));
 sky130_vsdinv _47362_ (.A(_16799_),
    .Y(_16800_));
 sky130_fd_sc_hd__a21o_4 _47363_ (.A1(_16658_),
    .A2(_16662_),
    .B1(_16800_),
    .X(_16801_));
 sky130_fd_sc_hd__buf_4 _47364_ (.A(_16800_),
    .X(_16802_));
 sky130_fd_sc_hd__nand3_4 _47365_ (.A(_16802_),
    .B(_16662_),
    .C(_16658_),
    .Y(_16803_));
 sky130_fd_sc_hd__nand2_4 _47366_ (.A(_16801_),
    .B(_16803_),
    .Y(_16804_));
 sky130_fd_sc_hd__xnor2_4 _47367_ (.A(_16797_),
    .B(_16804_),
    .Y(_16805_));
 sky130_fd_sc_hd__a21o_4 _47368_ (.A1(_16794_),
    .A2(_16795_),
    .B1(_16805_),
    .X(_16806_));
 sky130_fd_sc_hd__nand3_4 _47369_ (.A(_16794_),
    .B(_16795_),
    .C(_16805_),
    .Y(_16807_));
 sky130_fd_sc_hd__a21boi_4 _47370_ (.A1(_16669_),
    .A2(_16688_),
    .B1_N(_16670_),
    .Y(_16808_));
 sky130_vsdinv _47371_ (.A(_16808_),
    .Y(_16809_));
 sky130_fd_sc_hd__a21oi_4 _47372_ (.A1(_16806_),
    .A2(_16807_),
    .B1(_16809_),
    .Y(_16810_));
 sky130_vsdinv _47373_ (.A(_16810_),
    .Y(_16811_));
 sky130_fd_sc_hd__nand3_4 _47374_ (.A(_16806_),
    .B(_16807_),
    .C(_16809_),
    .Y(_16812_));
 sky130_vsdinv _47375_ (.A(_16671_),
    .Y(_16813_));
 sky130_fd_sc_hd__nand3_4 _47376_ (.A(_16685_),
    .B(_16813_),
    .C(_16686_),
    .Y(_16814_));
 sky130_fd_sc_hd__a21o_4 _47377_ (.A1(_16814_),
    .A2(_16686_),
    .B1(_16701_),
    .X(_16815_));
 sky130_fd_sc_hd__nand3_4 _47378_ (.A(_16814_),
    .B(_16701_),
    .C(_16686_),
    .Y(_16816_));
 sky130_fd_sc_hd__nand2_4 _47379_ (.A(_16815_),
    .B(_16816_),
    .Y(_16817_));
 sky130_fd_sc_hd__xor2_4 _47380_ (.A(_16697_),
    .B(_16817_),
    .X(_16818_));
 sky130_fd_sc_hd__a21o_4 _47381_ (.A1(_16811_),
    .A2(_16812_),
    .B1(_16818_),
    .X(_16819_));
 sky130_fd_sc_hd__nand3_4 _47382_ (.A(_16811_),
    .B(_16812_),
    .C(_16818_),
    .Y(_16820_));
 sky130_fd_sc_hd__nand2_4 _47383_ (.A(_16819_),
    .B(_16820_),
    .Y(_16821_));
 sky130_fd_sc_hd__a21boi_4 _47384_ (.A1(_16693_),
    .A2(_16704_),
    .B1_N(_16695_),
    .Y(_16822_));
 sky130_fd_sc_hd__nand2_4 _47385_ (.A(_16821_),
    .B(_16822_),
    .Y(_16823_));
 sky130_vsdinv _47386_ (.A(_16822_),
    .Y(_16824_));
 sky130_fd_sc_hd__nand3_4 _47387_ (.A(_16819_),
    .B(_16820_),
    .C(_16824_),
    .Y(_16825_));
 sky130_fd_sc_hd__nand2_4 _47388_ (.A(_16823_),
    .B(_16825_),
    .Y(_16826_));
 sky130_fd_sc_hd__buf_1 _47389_ (.A(_15964_),
    .X(_16827_));
 sky130_vsdinv _47390_ (.A(_16696_),
    .Y(_16828_));
 sky130_fd_sc_hd__buf_1 _47391_ (.A(_16828_),
    .X(_16829_));
 sky130_fd_sc_hd__a21bo_4 _47392_ (.A1(_16829_),
    .A2(_16702_),
    .B1_N(_16700_),
    .X(_16830_));
 sky130_fd_sc_hd__xor2_4 _47393_ (.A(_16587_),
    .B(_16830_),
    .X(_16831_));
 sky130_fd_sc_hd__xor2_4 _47394_ (.A(_16827_),
    .B(_16831_),
    .X(_16832_));
 sky130_vsdinv _47395_ (.A(_16832_),
    .Y(_16833_));
 sky130_fd_sc_hd__nand2_4 _47396_ (.A(_16826_),
    .B(_16833_),
    .Y(_16834_));
 sky130_fd_sc_hd__nand3_4 _47397_ (.A(_16823_),
    .B(_16825_),
    .C(_16832_),
    .Y(_16835_));
 sky130_fd_sc_hd__nand2_4 _47398_ (.A(_16834_),
    .B(_16835_),
    .Y(_16836_));
 sky130_fd_sc_hd__o21a_4 _47399_ (.A1(_16708_),
    .A2(_16716_),
    .B1(_16709_),
    .X(_16837_));
 sky130_fd_sc_hd__nand2_4 _47400_ (.A(_16836_),
    .B(_16837_),
    .Y(_16838_));
 sky130_vsdinv _47401_ (.A(_16837_),
    .Y(_16839_));
 sky130_fd_sc_hd__nand3_4 _47402_ (.A(_16834_),
    .B(_16835_),
    .C(_16839_),
    .Y(_16840_));
 sky130_fd_sc_hd__nand2_4 _47403_ (.A(_16838_),
    .B(_16840_),
    .Y(_16841_));
 sky130_fd_sc_hd__nand2_4 _47404_ (.A(_16714_),
    .B(_16711_),
    .Y(_16842_));
 sky130_fd_sc_hd__xor2_4 _47405_ (.A(_16149_),
    .B(_16842_),
    .X(_16843_));
 sky130_vsdinv _47406_ (.A(_16843_),
    .Y(_16844_));
 sky130_fd_sc_hd__nand2_4 _47407_ (.A(_16841_),
    .B(_16844_),
    .Y(_16845_));
 sky130_fd_sc_hd__nand3_4 _47408_ (.A(_16838_),
    .B(_16840_),
    .C(_16843_),
    .Y(_16846_));
 sky130_fd_sc_hd__nand2_4 _47409_ (.A(_16845_),
    .B(_16846_),
    .Y(_16847_));
 sky130_fd_sc_hd__a21boi_4 _47410_ (.A1(_16724_),
    .A2(_16728_),
    .B1_N(_16725_),
    .Y(_16848_));
 sky130_fd_sc_hd__nand2_4 _47411_ (.A(_16847_),
    .B(_16848_),
    .Y(_16849_));
 sky130_vsdinv _47412_ (.A(_16848_),
    .Y(_16850_));
 sky130_fd_sc_hd__nand3_4 _47413_ (.A(_16845_),
    .B(_16846_),
    .C(_16850_),
    .Y(_16851_));
 sky130_fd_sc_hd__buf_1 _47414_ (.A(_16314_),
    .X(_16852_));
 sky130_fd_sc_hd__a21oi_4 _47415_ (.A1(_16590_),
    .A2(_16586_),
    .B1(_16852_),
    .Y(_16853_));
 sky130_fd_sc_hd__a21o_4 _47416_ (.A1(_16849_),
    .A2(_16851_),
    .B1(_16853_),
    .X(_16854_));
 sky130_fd_sc_hd__nand3_4 _47417_ (.A(_16849_),
    .B(_16853_),
    .C(_16851_),
    .Y(_16855_));
 sky130_fd_sc_hd__nand2_4 _47418_ (.A(_16741_),
    .B(_16736_),
    .Y(_16856_));
 sky130_fd_sc_hd__a21oi_4 _47419_ (.A1(_16854_),
    .A2(_16855_),
    .B1(_16856_),
    .Y(_16857_));
 sky130_fd_sc_hd__nand3_4 _47420_ (.A(_16854_),
    .B(_16855_),
    .C(_16856_),
    .Y(_16858_));
 sky130_vsdinv _47421_ (.A(_16858_),
    .Y(_16859_));
 sky130_fd_sc_hd__nor2_4 _47422_ (.A(_16857_),
    .B(_16859_),
    .Y(_16860_));
 sky130_fd_sc_hd__nand4_4 _47423_ (.A(_16325_),
    .B(_16619_),
    .C(_16747_),
    .D(_16480_),
    .Y(_16861_));
 sky130_fd_sc_hd__nor2_4 _47424_ (.A(_16327_),
    .B(_16861_),
    .Y(_16862_));
 sky130_fd_sc_hd__nand2_4 _47425_ (.A(_16740_),
    .B(_16741_),
    .Y(_16863_));
 sky130_vsdinv _47426_ (.A(_16743_),
    .Y(_16864_));
 sky130_fd_sc_hd__nand2_4 _47427_ (.A(_16863_),
    .B(_16864_),
    .Y(_16865_));
 sky130_fd_sc_hd__nand4_4 _47428_ (.A(_16617_),
    .B(_16750_),
    .C(_16865_),
    .D(_16745_),
    .Y(_16866_));
 sky130_fd_sc_hd__nor2_4 _47429_ (.A(_16620_),
    .B(_16866_),
    .Y(_16867_));
 sky130_fd_sc_hd__nand2_4 _47430_ (.A(_16333_),
    .B(_16867_),
    .Y(_16868_));
 sky130_fd_sc_hd__a21oi_4 _47431_ (.A1(_16618_),
    .A2(_16865_),
    .B1(_16746_),
    .Y(_16869_));
 sky130_fd_sc_hd__o21a_4 _47432_ (.A1(_16622_),
    .A2(_16866_),
    .B1(_16869_),
    .X(_16870_));
 sky130_fd_sc_hd__nand2_4 _47433_ (.A(_16868_),
    .B(_16870_),
    .Y(_16871_));
 sky130_fd_sc_hd__a21oi_4 _47434_ (.A1(_15651_),
    .A2(_16862_),
    .B1(_16871_),
    .Y(_16872_));
 sky130_fd_sc_hd__xnor2_4 _47435_ (.A(_16860_),
    .B(_16872_),
    .Y(_01461_));
 sky130_fd_sc_hd__a21boi_4 _47436_ (.A1(_16823_),
    .A2(_16832_),
    .B1_N(_16825_),
    .Y(_16873_));
 sky130_vsdinv _47437_ (.A(_16873_),
    .Y(_16874_));
 sky130_fd_sc_hd__nand4_4 _47438_ (.A(_16752_),
    .B(_16754_),
    .C(_03624_),
    .D(_16755_),
    .Y(_16875_));
 sky130_fd_sc_hd__buf_1 _47439_ (.A(_16040_),
    .X(_16876_));
 sky130_fd_sc_hd__nand2_4 _47440_ (.A(_16876_),
    .B(_03623_),
    .Y(_16877_));
 sky130_fd_sc_hd__a2bb2o_4 _47441_ (.A1_N(_16037_),
    .A2_N(_03635_),
    .B1(_16752_),
    .B2(_16624_),
    .X(_16878_));
 sky130_fd_sc_hd__nand4_4 _47442_ (.A(_03377_),
    .B(_16038_),
    .C(_16338_),
    .D(_11386_),
    .Y(_16879_));
 sky130_fd_sc_hd__and2_4 _47443_ (.A(_16878_),
    .B(_16879_),
    .X(_16880_));
 sky130_fd_sc_hd__xor2_4 _47444_ (.A(_16877_),
    .B(_16880_),
    .X(_16881_));
 sky130_fd_sc_hd__a21o_4 _47445_ (.A1(_16755_),
    .A2(_16875_),
    .B1(_16881_),
    .X(_16882_));
 sky130_fd_sc_hd__nand3_4 _47446_ (.A(_16881_),
    .B(_16755_),
    .C(_16875_),
    .Y(_16883_));
 sky130_fd_sc_hd__nand2_4 _47447_ (.A(_16517_),
    .B(_03603_),
    .Y(_16884_));
 sky130_fd_sc_hd__nand2_4 _47448_ (.A(_16762_),
    .B(_03616_),
    .Y(_16885_));
 sky130_fd_sc_hd__buf_1 _47449_ (.A(_10844_),
    .X(_16886_));
 sky130_fd_sc_hd__nand2_4 _47450_ (.A(_16886_),
    .B(_03609_),
    .Y(_16887_));
 sky130_fd_sc_hd__xnor2_4 _47451_ (.A(_16885_),
    .B(_16887_),
    .Y(_16888_));
 sky130_fd_sc_hd__xor2_4 _47452_ (.A(_16884_),
    .B(_16888_),
    .X(_16889_));
 sky130_fd_sc_hd__a21o_4 _47453_ (.A1(_16882_),
    .A2(_16883_),
    .B1(_16889_),
    .X(_16890_));
 sky130_fd_sc_hd__nand3_4 _47454_ (.A(_16882_),
    .B(_16883_),
    .C(_16889_),
    .Y(_16891_));
 sky130_fd_sc_hd__a21boi_4 _47455_ (.A1(_16759_),
    .A2(_16765_),
    .B1_N(_16758_),
    .Y(_16892_));
 sky130_fd_sc_hd__a21boi_4 _47456_ (.A1(_16890_),
    .A2(_16891_),
    .B1_N(_16892_),
    .Y(_16893_));
 sky130_vsdinv _47457_ (.A(_16892_),
    .Y(_16894_));
 sky130_fd_sc_hd__nand3_4 _47458_ (.A(_16894_),
    .B(_16890_),
    .C(_16891_),
    .Y(_16895_));
 sky130_vsdinv _47459_ (.A(_16895_),
    .Y(_16896_));
 sky130_vsdinv _47460_ (.A(_16540_),
    .Y(_16897_));
 sky130_fd_sc_hd__a2bb2o_4 _47461_ (.A1_N(_16897_),
    .A2_N(_16649_),
    .B1(_10838_),
    .B2(_03598_),
    .X(_16898_));
 sky130_fd_sc_hd__nand4_4 _47462_ (.A(_16543_),
    .B(_03409_),
    .C(_03589_),
    .D(_03598_),
    .Y(_16899_));
 sky130_fd_sc_hd__a21o_4 _47463_ (.A1(_16898_),
    .A2(_16899_),
    .B1(_16777_),
    .X(_16900_));
 sky130_fd_sc_hd__nand3_4 _47464_ (.A(_16898_),
    .B(_16899_),
    .C(_16777_),
    .Y(_16901_));
 sky130_fd_sc_hd__maj3_4 _47465_ (.A(_16761_),
    .B(_16763_),
    .C(_16760_),
    .X(_16902_));
 sky130_vsdinv _47466_ (.A(_16902_),
    .Y(_16903_));
 sky130_fd_sc_hd__a21o_4 _47467_ (.A1(_16900_),
    .A2(_16901_),
    .B1(_16903_),
    .X(_16904_));
 sky130_fd_sc_hd__nand3_4 _47468_ (.A(_16900_),
    .B(_16903_),
    .C(_16901_),
    .Y(_16905_));
 sky130_fd_sc_hd__nand2_4 _47469_ (.A(_16904_),
    .B(_16905_),
    .Y(_16906_));
 sky130_fd_sc_hd__a21o_4 _47470_ (.A1(_16774_),
    .A2(_16779_),
    .B1(_16906_),
    .X(_16907_));
 sky130_fd_sc_hd__nand3_4 _47471_ (.A(_16906_),
    .B(_16774_),
    .C(_16779_),
    .Y(_16908_));
 sky130_fd_sc_hd__and2_4 _47472_ (.A(_16907_),
    .B(_16908_),
    .X(_16909_));
 sky130_vsdinv _47473_ (.A(_16909_),
    .Y(_16910_));
 sky130_fd_sc_hd__o21ai_4 _47474_ (.A1(_16893_),
    .A2(_16896_),
    .B1(_16910_),
    .Y(_16911_));
 sky130_vsdinv _47475_ (.A(_16893_),
    .Y(_16912_));
 sky130_fd_sc_hd__nand3_4 _47476_ (.A(_16912_),
    .B(_16895_),
    .C(_16909_),
    .Y(_16913_));
 sky130_fd_sc_hd__o21a_4 _47477_ (.A1(_16788_),
    .A2(_16770_),
    .B1(_16771_),
    .X(_16914_));
 sky130_fd_sc_hd__a21boi_4 _47478_ (.A1(_16911_),
    .A2(_16913_),
    .B1_N(_16914_),
    .Y(_16915_));
 sky130_vsdinv _47479_ (.A(_16914_),
    .Y(_16916_));
 sky130_fd_sc_hd__nand3_4 _47480_ (.A(_16916_),
    .B(_16911_),
    .C(_16913_),
    .Y(_16917_));
 sky130_vsdinv _47481_ (.A(_16917_),
    .Y(_16918_));
 sky130_fd_sc_hd__a21o_4 _47482_ (.A1(_16785_),
    .A2(_16783_),
    .B1(_16802_),
    .X(_16919_));
 sky130_fd_sc_hd__nand3_4 _47483_ (.A(_16785_),
    .B(_16783_),
    .C(_16802_),
    .Y(_16920_));
 sky130_fd_sc_hd__buf_1 _47484_ (.A(_03409_),
    .X(_16921_));
 sky130_fd_sc_hd__a21o_4 _47485_ (.A1(_16921_),
    .A2(_03566_),
    .B1(_16672_),
    .X(_16922_));
 sky130_vsdinv _47486_ (.A(_16796_),
    .Y(_16923_));
 sky130_fd_sc_hd__a21oi_4 _47487_ (.A1(_16536_),
    .A2(_16922_),
    .B1(_16923_),
    .Y(_16924_));
 sky130_vsdinv _47488_ (.A(_16924_),
    .Y(_16925_));
 sky130_fd_sc_hd__a21o_4 _47489_ (.A1(_16919_),
    .A2(_16920_),
    .B1(_16925_),
    .X(_16926_));
 sky130_fd_sc_hd__buf_1 _47490_ (.A(_16925_),
    .X(_16927_));
 sky130_fd_sc_hd__nand3_4 _47491_ (.A(_16919_),
    .B(_16927_),
    .C(_16920_),
    .Y(_16928_));
 sky130_fd_sc_hd__and2_4 _47492_ (.A(_16926_),
    .B(_16928_),
    .X(_16929_));
 sky130_vsdinv _47493_ (.A(_16929_),
    .Y(_16930_));
 sky130_fd_sc_hd__o21ai_4 _47494_ (.A1(_16915_),
    .A2(_16918_),
    .B1(_16930_),
    .Y(_16931_));
 sky130_vsdinv _47495_ (.A(_16915_),
    .Y(_16932_));
 sky130_fd_sc_hd__nand3_4 _47496_ (.A(_16932_),
    .B(_16917_),
    .C(_16929_),
    .Y(_16933_));
 sky130_fd_sc_hd__a21boi_4 _47497_ (.A1(_16794_),
    .A2(_16805_),
    .B1_N(_16795_),
    .Y(_16934_));
 sky130_vsdinv _47498_ (.A(_16934_),
    .Y(_16935_));
 sky130_fd_sc_hd__a21oi_4 _47499_ (.A1(_16931_),
    .A2(_16933_),
    .B1(_16935_),
    .Y(_16936_));
 sky130_fd_sc_hd__nand3_4 _47500_ (.A(_16935_),
    .B(_16931_),
    .C(_16933_),
    .Y(_16937_));
 sky130_vsdinv _47501_ (.A(_16937_),
    .Y(_16938_));
 sky130_fd_sc_hd__a21boi_4 _47502_ (.A1(_16803_),
    .A2(_16797_),
    .B1_N(_16801_),
    .Y(_16939_));
 sky130_fd_sc_hd__or2_4 _47503_ (.A(_16569_),
    .B(_16939_),
    .X(_16940_));
 sky130_fd_sc_hd__buf_1 _47504_ (.A(_16940_),
    .X(_16941_));
 sky130_fd_sc_hd__nand2_4 _47505_ (.A(_16939_),
    .B(_16701_),
    .Y(_16942_));
 sky130_fd_sc_hd__a21o_4 _47506_ (.A1(_16941_),
    .A2(_16942_),
    .B1(_16828_),
    .X(_16943_));
 sky130_fd_sc_hd__nand3_4 _47507_ (.A(_16941_),
    .B(_16828_),
    .C(_16942_),
    .Y(_16944_));
 sky130_fd_sc_hd__and2_4 _47508_ (.A(_16943_),
    .B(_16944_),
    .X(_16945_));
 sky130_vsdinv _47509_ (.A(_16945_),
    .Y(_16946_));
 sky130_fd_sc_hd__o21ai_4 _47510_ (.A1(_16936_),
    .A2(_16938_),
    .B1(_16946_),
    .Y(_16947_));
 sky130_vsdinv _47511_ (.A(_16936_),
    .Y(_16948_));
 sky130_fd_sc_hd__nand3_4 _47512_ (.A(_16948_),
    .B(_16937_),
    .C(_16945_),
    .Y(_16949_));
 sky130_vsdinv _47513_ (.A(_16818_),
    .Y(_16950_));
 sky130_fd_sc_hd__o21a_4 _47514_ (.A1(_16950_),
    .A2(_16810_),
    .B1(_16812_),
    .X(_16951_));
 sky130_fd_sc_hd__a21boi_4 _47515_ (.A1(_16947_),
    .A2(_16949_),
    .B1_N(_16951_),
    .Y(_16952_));
 sky130_vsdinv _47516_ (.A(_16951_),
    .Y(_16953_));
 sky130_fd_sc_hd__nand3_4 _47517_ (.A(_16953_),
    .B(_16947_),
    .C(_16949_),
    .Y(_16954_));
 sky130_vsdinv _47518_ (.A(_16954_),
    .Y(_16955_));
 sky130_fd_sc_hd__a21bo_4 _47519_ (.A1(_16828_),
    .A2(_16816_),
    .B1_N(_16815_),
    .X(_16956_));
 sky130_fd_sc_hd__or2_4 _47520_ (.A(_15785_),
    .B(_16956_),
    .X(_16957_));
 sky130_fd_sc_hd__nand2_4 _47521_ (.A(_16956_),
    .B(_15785_),
    .Y(_16958_));
 sky130_fd_sc_hd__a21o_4 _47522_ (.A1(_16957_),
    .A2(_16958_),
    .B1(_16444_),
    .X(_16959_));
 sky130_fd_sc_hd__buf_1 _47523_ (.A(_16290_),
    .X(_16960_));
 sky130_fd_sc_hd__nand3_4 _47524_ (.A(_16957_),
    .B(_16960_),
    .C(_16958_),
    .Y(_16961_));
 sky130_fd_sc_hd__and2_4 _47525_ (.A(_16959_),
    .B(_16961_),
    .X(_16962_));
 sky130_vsdinv _47526_ (.A(_16962_),
    .Y(_16963_));
 sky130_fd_sc_hd__o21ai_4 _47527_ (.A1(_16952_),
    .A2(_16955_),
    .B1(_16963_),
    .Y(_16964_));
 sky130_vsdinv _47528_ (.A(_16952_),
    .Y(_16965_));
 sky130_fd_sc_hd__nand3_4 _47529_ (.A(_16965_),
    .B(_16954_),
    .C(_16962_),
    .Y(_16966_));
 sky130_fd_sc_hd__nand3_4 _47530_ (.A(_16874_),
    .B(_16964_),
    .C(_16966_),
    .Y(_16967_));
 sky130_fd_sc_hd__nand2_4 _47531_ (.A(_16964_),
    .B(_16966_),
    .Y(_16968_));
 sky130_fd_sc_hd__nand2_4 _47532_ (.A(_16968_),
    .B(_16873_),
    .Y(_16969_));
 sky130_fd_sc_hd__nand2_4 _47533_ (.A(_16967_),
    .B(_16969_),
    .Y(_16970_));
 sky130_fd_sc_hd__buf_1 _47534_ (.A(_15785_),
    .X(_16971_));
 sky130_fd_sc_hd__buf_1 _47535_ (.A(_16971_),
    .X(_16972_));
 sky130_fd_sc_hd__maj3_4 _47536_ (.A(_16972_),
    .B(_16830_),
    .C(_16960_),
    .X(_16973_));
 sky130_fd_sc_hd__xor2_4 _47537_ (.A(_16149_),
    .B(_16973_),
    .X(_16974_));
 sky130_vsdinv _47538_ (.A(_16974_),
    .Y(_16975_));
 sky130_fd_sc_hd__nand2_4 _47539_ (.A(_16970_),
    .B(_16975_),
    .Y(_16976_));
 sky130_fd_sc_hd__nand3_4 _47540_ (.A(_16967_),
    .B(_16969_),
    .C(_16974_),
    .Y(_16977_));
 sky130_fd_sc_hd__nand2_4 _47541_ (.A(_16976_),
    .B(_16977_),
    .Y(_16978_));
 sky130_fd_sc_hd__a21boi_4 _47542_ (.A1(_16838_),
    .A2(_16843_),
    .B1_N(_16840_),
    .Y(_16979_));
 sky130_fd_sc_hd__nand2_4 _47543_ (.A(_16978_),
    .B(_16979_),
    .Y(_16980_));
 sky130_vsdinv _47544_ (.A(_16979_),
    .Y(_16981_));
 sky130_fd_sc_hd__nand3_4 _47545_ (.A(_16981_),
    .B(_16976_),
    .C(_16977_),
    .Y(_16982_));
 sky130_fd_sc_hd__nand2_4 _47546_ (.A(_16980_),
    .B(_16982_),
    .Y(_16983_));
 sky130_fd_sc_hd__a21oi_4 _47547_ (.A1(_16714_),
    .A2(_16711_),
    .B1(_16852_),
    .Y(_16984_));
 sky130_vsdinv _47548_ (.A(_16984_),
    .Y(_16985_));
 sky130_fd_sc_hd__nand2_4 _47549_ (.A(_16983_),
    .B(_16985_),
    .Y(_16986_));
 sky130_fd_sc_hd__nand3_4 _47550_ (.A(_16980_),
    .B(_16982_),
    .C(_16984_),
    .Y(_16987_));
 sky130_fd_sc_hd__nand2_4 _47551_ (.A(_16986_),
    .B(_16987_),
    .Y(_16988_));
 sky130_fd_sc_hd__a21boi_4 _47552_ (.A1(_16849_),
    .A2(_16853_),
    .B1_N(_16851_),
    .Y(_16989_));
 sky130_fd_sc_hd__nand2_4 _47553_ (.A(_16988_),
    .B(_16989_),
    .Y(_16990_));
 sky130_vsdinv _47554_ (.A(_16989_),
    .Y(_16991_));
 sky130_fd_sc_hd__nand3_4 _47555_ (.A(_16991_),
    .B(_16986_),
    .C(_16987_),
    .Y(_16992_));
 sky130_fd_sc_hd__and2_4 _47556_ (.A(_16990_),
    .B(_16992_),
    .X(_16993_));
 sky130_fd_sc_hd__buf_1 _47557_ (.A(_16993_),
    .X(_16994_));
 sky130_fd_sc_hd__o21ai_4 _47558_ (.A1(_16857_),
    .A2(_16872_),
    .B1(_16858_),
    .Y(_16995_));
 sky130_fd_sc_hd__xor2_4 _47559_ (.A(_16994_),
    .B(_16995_),
    .X(_01462_));
 sky130_fd_sc_hd__buf_1 _47560_ (.A(_03623_),
    .X(_16996_));
 sky130_fd_sc_hd__nand4_4 _47561_ (.A(_16876_),
    .B(_16878_),
    .C(_16996_),
    .D(_16879_),
    .Y(_16997_));
 sky130_fd_sc_hd__buf_1 _47562_ (.A(_16762_),
    .X(_16998_));
 sky130_fd_sc_hd__nand2_4 _47563_ (.A(_16998_),
    .B(_03624_),
    .Y(_16999_));
 sky130_fd_sc_hd__buf_1 _47564_ (.A(_16338_),
    .X(_17000_));
 sky130_fd_sc_hd__a2bb2o_4 _47565_ (.A1_N(_16752_),
    .A2_N(_03636_),
    .B1(_16876_),
    .B2(_17000_),
    .X(_17001_));
 sky130_fd_sc_hd__nand4_4 _47566_ (.A(_03380_),
    .B(_16040_),
    .C(_17000_),
    .D(_11386_),
    .Y(_17002_));
 sky130_fd_sc_hd__and2_4 _47567_ (.A(_17001_),
    .B(_17002_),
    .X(_17003_));
 sky130_fd_sc_hd__xor2_4 _47568_ (.A(_16999_),
    .B(_17003_),
    .X(_17004_));
 sky130_fd_sc_hd__a21o_4 _47569_ (.A1(_16879_),
    .A2(_16997_),
    .B1(_17004_),
    .X(_17005_));
 sky130_fd_sc_hd__nand3_4 _47570_ (.A(_17004_),
    .B(_16879_),
    .C(_16997_),
    .Y(_17006_));
 sky130_fd_sc_hd__buf_1 _47571_ (.A(_16543_),
    .X(_17007_));
 sky130_fd_sc_hd__nand2_4 _47572_ (.A(_17007_),
    .B(_03603_),
    .Y(_17008_));
 sky130_fd_sc_hd__buf_1 _47573_ (.A(_16886_),
    .X(_17009_));
 sky130_fd_sc_hd__nand2_4 _47574_ (.A(_17009_),
    .B(_03616_),
    .Y(_17010_));
 sky130_fd_sc_hd__buf_4 _47575_ (.A(_16517_),
    .X(_17011_));
 sky130_fd_sc_hd__nand2_4 _47576_ (.A(_17011_),
    .B(_03609_),
    .Y(_17012_));
 sky130_fd_sc_hd__xnor2_4 _47577_ (.A(_17010_),
    .B(_17012_),
    .Y(_17013_));
 sky130_fd_sc_hd__xor2_4 _47578_ (.A(_17008_),
    .B(_17013_),
    .X(_17014_));
 sky130_fd_sc_hd__a21o_4 _47579_ (.A1(_17005_),
    .A2(_17006_),
    .B1(_17014_),
    .X(_17015_));
 sky130_fd_sc_hd__nand3_4 _47580_ (.A(_17005_),
    .B(_17006_),
    .C(_17014_),
    .Y(_17016_));
 sky130_fd_sc_hd__a21boi_4 _47581_ (.A1(_16883_),
    .A2(_16889_),
    .B1_N(_16882_),
    .Y(_17017_));
 sky130_fd_sc_hd__a21boi_4 _47582_ (.A1(_17015_),
    .A2(_17016_),
    .B1_N(_17017_),
    .Y(_17018_));
 sky130_vsdinv _47583_ (.A(_17017_),
    .Y(_17019_));
 sky130_fd_sc_hd__nand3_4 _47584_ (.A(_17019_),
    .B(_17015_),
    .C(_17016_),
    .Y(_17020_));
 sky130_vsdinv _47585_ (.A(_17020_),
    .Y(_17021_));
 sky130_fd_sc_hd__maj3_4 _47586_ (.A(_16885_),
    .B(_16887_),
    .C(_16884_),
    .X(_17022_));
 sky130_fd_sc_hd__o21a_4 _47587_ (.A1(_16512_),
    .A2(_15499_),
    .B1(_12910_),
    .X(_17023_));
 sky130_fd_sc_hd__nand3_4 _47588_ (.A(_03408_),
    .B(_15860_),
    .C(_15858_),
    .Y(_17024_));
 sky130_fd_sc_hd__a21o_4 _47589_ (.A1(_17023_),
    .A2(_17024_),
    .B1(_16776_),
    .X(_17025_));
 sky130_fd_sc_hd__nand3_4 _47590_ (.A(_17023_),
    .B(_16776_),
    .C(_17024_),
    .Y(_17026_));
 sky130_fd_sc_hd__and2_4 _47591_ (.A(_17025_),
    .B(_17026_),
    .X(_17027_));
 sky130_fd_sc_hd__buf_1 _47592_ (.A(_17027_),
    .X(_17028_));
 sky130_fd_sc_hd__xor2_4 _47593_ (.A(_17022_),
    .B(_17028_),
    .X(_17029_));
 sky130_fd_sc_hd__a21o_4 _47594_ (.A1(_16899_),
    .A2(_16901_),
    .B1(_17029_),
    .X(_17030_));
 sky130_fd_sc_hd__nand3_4 _47595_ (.A(_17029_),
    .B(_16899_),
    .C(_16901_),
    .Y(_17031_));
 sky130_fd_sc_hd__and2_4 _47596_ (.A(_17030_),
    .B(_17031_),
    .X(_17032_));
 sky130_vsdinv _47597_ (.A(_17032_),
    .Y(_17033_));
 sky130_fd_sc_hd__o21ai_4 _47598_ (.A1(_17018_),
    .A2(_17021_),
    .B1(_17033_),
    .Y(_17034_));
 sky130_vsdinv _47599_ (.A(_17018_),
    .Y(_17035_));
 sky130_fd_sc_hd__nand3_4 _47600_ (.A(_17035_),
    .B(_17020_),
    .C(_17032_),
    .Y(_17036_));
 sky130_fd_sc_hd__o21a_4 _47601_ (.A1(_16910_),
    .A2(_16893_),
    .B1(_16895_),
    .X(_17037_));
 sky130_fd_sc_hd__a21boi_4 _47602_ (.A1(_17034_),
    .A2(_17036_),
    .B1_N(_17037_),
    .Y(_17038_));
 sky130_vsdinv _47603_ (.A(_17037_),
    .Y(_17039_));
 sky130_fd_sc_hd__nand3_4 _47604_ (.A(_17039_),
    .B(_17034_),
    .C(_17036_),
    .Y(_17040_));
 sky130_vsdinv _47605_ (.A(_17040_),
    .Y(_17041_));
 sky130_fd_sc_hd__buf_4 _47606_ (.A(_16802_),
    .X(_17042_));
 sky130_fd_sc_hd__a21o_4 _47607_ (.A1(_16907_),
    .A2(_16905_),
    .B1(_17042_),
    .X(_17043_));
 sky130_fd_sc_hd__nand3_4 _47608_ (.A(_16907_),
    .B(_17042_),
    .C(_16905_),
    .Y(_17044_));
 sky130_fd_sc_hd__a21o_4 _47609_ (.A1(_17043_),
    .A2(_17044_),
    .B1(_16927_),
    .X(_17045_));
 sky130_fd_sc_hd__nand3_4 _47610_ (.A(_17043_),
    .B(_16927_),
    .C(_17044_),
    .Y(_17046_));
 sky130_fd_sc_hd__and2_4 _47611_ (.A(_17045_),
    .B(_17046_),
    .X(_17047_));
 sky130_vsdinv _47612_ (.A(_17047_),
    .Y(_17048_));
 sky130_fd_sc_hd__o21ai_4 _47613_ (.A1(_17038_),
    .A2(_17041_),
    .B1(_17048_),
    .Y(_17049_));
 sky130_vsdinv _47614_ (.A(_17038_),
    .Y(_17050_));
 sky130_fd_sc_hd__nand3_4 _47615_ (.A(_17050_),
    .B(_17040_),
    .C(_17047_),
    .Y(_17051_));
 sky130_fd_sc_hd__o21a_4 _47616_ (.A1(_16930_),
    .A2(_16915_),
    .B1(_16917_),
    .X(_17052_));
 sky130_fd_sc_hd__a21boi_4 _47617_ (.A1(_17049_),
    .A2(_17051_),
    .B1_N(_17052_),
    .Y(_17053_));
 sky130_vsdinv _47618_ (.A(_17052_),
    .Y(_17054_));
 sky130_fd_sc_hd__nand3_4 _47619_ (.A(_17054_),
    .B(_17049_),
    .C(_17051_),
    .Y(_17055_));
 sky130_vsdinv _47620_ (.A(_17055_),
    .Y(_17056_));
 sky130_fd_sc_hd__buf_1 _47621_ (.A(_16570_),
    .X(_17057_));
 sky130_fd_sc_hd__a21o_4 _47622_ (.A1(_16928_),
    .A2(_16919_),
    .B1(_17057_),
    .X(_17058_));
 sky130_fd_sc_hd__nand3_4 _47623_ (.A(_16928_),
    .B(_17057_),
    .C(_16919_),
    .Y(_17059_));
 sky130_fd_sc_hd__nand2_4 _47624_ (.A(_17058_),
    .B(_17059_),
    .Y(_17060_));
 sky130_fd_sc_hd__xor2_4 _47625_ (.A(_16697_),
    .B(_17060_),
    .X(_17061_));
 sky130_vsdinv _47626_ (.A(_17061_),
    .Y(_17062_));
 sky130_fd_sc_hd__o21ai_4 _47627_ (.A1(_17053_),
    .A2(_17056_),
    .B1(_17062_),
    .Y(_17063_));
 sky130_vsdinv _47628_ (.A(_17053_),
    .Y(_17064_));
 sky130_fd_sc_hd__nand3_4 _47629_ (.A(_17064_),
    .B(_17055_),
    .C(_17061_),
    .Y(_17065_));
 sky130_fd_sc_hd__o21a_4 _47630_ (.A1(_16946_),
    .A2(_16936_),
    .B1(_16937_),
    .X(_17066_));
 sky130_vsdinv _47631_ (.A(_17066_),
    .Y(_17067_));
 sky130_fd_sc_hd__a21o_4 _47632_ (.A1(_17063_),
    .A2(_17065_),
    .B1(_17067_),
    .X(_17068_));
 sky130_fd_sc_hd__nand3_4 _47633_ (.A(_17067_),
    .B(_17063_),
    .C(_17065_),
    .Y(_17069_));
 sky130_fd_sc_hd__a21o_4 _47634_ (.A1(_16944_),
    .A2(_16941_),
    .B1(_16587_),
    .X(_17070_));
 sky130_fd_sc_hd__buf_1 _47635_ (.A(_16587_),
    .X(_17071_));
 sky130_fd_sc_hd__nand3_4 _47636_ (.A(_16944_),
    .B(_17071_),
    .C(_16941_),
    .Y(_17072_));
 sky130_fd_sc_hd__and2_4 _47637_ (.A(_17070_),
    .B(_17072_),
    .X(_17073_));
 sky130_fd_sc_hd__xor2_4 _47638_ (.A(_16960_),
    .B(_17073_),
    .X(_17074_));
 sky130_fd_sc_hd__a21o_4 _47639_ (.A1(_17068_),
    .A2(_17069_),
    .B1(_17074_),
    .X(_17075_));
 sky130_fd_sc_hd__nand3_4 _47640_ (.A(_17068_),
    .B(_17074_),
    .C(_17069_),
    .Y(_17076_));
 sky130_fd_sc_hd__nand2_4 _47641_ (.A(_17075_),
    .B(_17076_),
    .Y(_17077_));
 sky130_fd_sc_hd__o21a_4 _47642_ (.A1(_16963_),
    .A2(_16952_),
    .B1(_16954_),
    .X(_17078_));
 sky130_fd_sc_hd__nand2_4 _47643_ (.A(_17077_),
    .B(_17078_),
    .Y(_17079_));
 sky130_vsdinv _47644_ (.A(_17078_),
    .Y(_17080_));
 sky130_fd_sc_hd__nand3_4 _47645_ (.A(_17080_),
    .B(_17075_),
    .C(_17076_),
    .Y(_17081_));
 sky130_fd_sc_hd__nand2_4 _47646_ (.A(_17079_),
    .B(_17081_),
    .Y(_17082_));
 sky130_fd_sc_hd__buf_1 _47647_ (.A(_16960_),
    .X(_17083_));
 sky130_fd_sc_hd__maj3_4 _47648_ (.A(_16972_),
    .B(_16956_),
    .C(_17083_),
    .X(_17084_));
 sky130_fd_sc_hd__xor2_4 _47649_ (.A(_16149_),
    .B(_17084_),
    .X(_17085_));
 sky130_vsdinv _47650_ (.A(_17085_),
    .Y(_17086_));
 sky130_fd_sc_hd__nand2_4 _47651_ (.A(_17082_),
    .B(_17086_),
    .Y(_17087_));
 sky130_fd_sc_hd__nand3_4 _47652_ (.A(_17079_),
    .B(_17081_),
    .C(_17085_),
    .Y(_17088_));
 sky130_fd_sc_hd__nand2_4 _47653_ (.A(_17087_),
    .B(_17088_),
    .Y(_17089_));
 sky130_fd_sc_hd__nand2_4 _47654_ (.A(_16977_),
    .B(_16967_),
    .Y(_17090_));
 sky130_vsdinv _47655_ (.A(_17090_),
    .Y(_17091_));
 sky130_fd_sc_hd__nand2_4 _47656_ (.A(_17089_),
    .B(_17091_),
    .Y(_17092_));
 sky130_fd_sc_hd__nand3_4 _47657_ (.A(_17087_),
    .B(_17090_),
    .C(_17088_),
    .Y(_17093_));
 sky130_fd_sc_hd__nand2_4 _47658_ (.A(_17092_),
    .B(_17093_),
    .Y(_17094_));
 sky130_fd_sc_hd__buf_1 _47659_ (.A(_16150_),
    .X(_17095_));
 sky130_fd_sc_hd__and2_4 _47660_ (.A(_16973_),
    .B(_17095_),
    .X(_17096_));
 sky130_vsdinv _47661_ (.A(_17096_),
    .Y(_17097_));
 sky130_fd_sc_hd__nand2_4 _47662_ (.A(_17094_),
    .B(_17097_),
    .Y(_17098_));
 sky130_fd_sc_hd__nand3_4 _47663_ (.A(_17092_),
    .B(_17096_),
    .C(_17093_),
    .Y(_17099_));
 sky130_fd_sc_hd__a21boi_4 _47664_ (.A1(_16976_),
    .A2(_16977_),
    .B1_N(_16979_),
    .Y(_17100_));
 sky130_fd_sc_hd__o21ai_4 _47665_ (.A1(_16985_),
    .A2(_17100_),
    .B1(_16982_),
    .Y(_17101_));
 sky130_fd_sc_hd__a21oi_4 _47666_ (.A1(_17098_),
    .A2(_17099_),
    .B1(_17101_),
    .Y(_17102_));
 sky130_fd_sc_hd__nand3_4 _47667_ (.A(_17098_),
    .B(_17101_),
    .C(_17099_),
    .Y(_17103_));
 sky130_vsdinv _47668_ (.A(_17103_),
    .Y(_17104_));
 sky130_fd_sc_hd__nor2_4 _47669_ (.A(_17102_),
    .B(_17104_),
    .Y(_17105_));
 sky130_vsdinv _47670_ (.A(_16872_),
    .Y(_17106_));
 sky130_fd_sc_hd__and2_4 _47671_ (.A(_16994_),
    .B(_16860_),
    .X(_17107_));
 sky130_fd_sc_hd__nand2_4 _47672_ (.A(_16992_),
    .B(_16858_),
    .Y(_17108_));
 sky130_fd_sc_hd__nand2_4 _47673_ (.A(_17108_),
    .B(_16990_),
    .Y(_17109_));
 sky130_fd_sc_hd__a21bo_4 _47674_ (.A1(_17106_),
    .A2(_17107_),
    .B1_N(_17109_),
    .X(_17110_));
 sky130_fd_sc_hd__xor2_4 _47675_ (.A(_17105_),
    .B(_17110_),
    .X(_01463_));
 sky130_fd_sc_hd__nand4_4 _47676_ (.A(_16998_),
    .B(_17001_),
    .C(_03625_),
    .D(_17002_),
    .Y(_17111_));
 sky130_fd_sc_hd__nand2_4 _47677_ (.A(_17009_),
    .B(_16996_),
    .Y(_17112_));
 sky130_fd_sc_hd__buf_4 _47678_ (.A(_16624_),
    .X(_17113_));
 sky130_fd_sc_hd__a2bb2o_4 _47679_ (.A1_N(_16876_),
    .A2_N(_03636_),
    .B1(_16998_),
    .B2(_17113_),
    .X(_17114_));
 sky130_fd_sc_hd__nand4_4 _47680_ (.A(_03384_),
    .B(_16998_),
    .C(_17113_),
    .D(_11387_),
    .Y(_17115_));
 sky130_fd_sc_hd__and2_4 _47681_ (.A(_17114_),
    .B(_17115_),
    .X(_17116_));
 sky130_fd_sc_hd__xor2_4 _47682_ (.A(_17112_),
    .B(_17116_),
    .X(_17117_));
 sky130_fd_sc_hd__a21o_4 _47683_ (.A1(_17002_),
    .A2(_17111_),
    .B1(_17117_),
    .X(_17118_));
 sky130_fd_sc_hd__nand3_4 _47684_ (.A(_17117_),
    .B(_17002_),
    .C(_17111_),
    .Y(_17119_));
 sky130_fd_sc_hd__nand2_4 _47685_ (.A(_16921_),
    .B(_03603_),
    .Y(_17120_));
 sky130_fd_sc_hd__buf_1 _47686_ (.A(_17120_),
    .X(_17121_));
 sky130_fd_sc_hd__buf_4 _47687_ (.A(_17011_),
    .X(_17122_));
 sky130_fd_sc_hd__nand2_4 _47688_ (.A(_17122_),
    .B(_03616_),
    .Y(_17123_));
 sky130_fd_sc_hd__nand2_4 _47689_ (.A(_17007_),
    .B(_03610_),
    .Y(_17124_));
 sky130_fd_sc_hd__xnor2_4 _47690_ (.A(_17123_),
    .B(_17124_),
    .Y(_17125_));
 sky130_fd_sc_hd__xor2_4 _47691_ (.A(_17121_),
    .B(_17125_),
    .X(_17126_));
 sky130_fd_sc_hd__a21o_4 _47692_ (.A1(_17118_),
    .A2(_17119_),
    .B1(_17126_),
    .X(_17127_));
 sky130_fd_sc_hd__nand3_4 _47693_ (.A(_17118_),
    .B(_17119_),
    .C(_17126_),
    .Y(_17128_));
 sky130_fd_sc_hd__a21boi_4 _47694_ (.A1(_17006_),
    .A2(_17014_),
    .B1_N(_17005_),
    .Y(_17129_));
 sky130_vsdinv _47695_ (.A(_17129_),
    .Y(_17130_));
 sky130_fd_sc_hd__a21o_4 _47696_ (.A1(_17127_),
    .A2(_17128_),
    .B1(_17130_),
    .X(_17131_));
 sky130_fd_sc_hd__nand3_4 _47697_ (.A(_17130_),
    .B(_17127_),
    .C(_17128_),
    .Y(_17132_));
 sky130_fd_sc_hd__a21boi_4 _47698_ (.A1(_17023_),
    .A2(_16777_),
    .B1_N(_17024_),
    .Y(_17133_));
 sky130_fd_sc_hd__maj3_4 _47699_ (.A(_17010_),
    .B(_17012_),
    .C(_17008_),
    .X(_17134_));
 sky130_vsdinv _47700_ (.A(_17134_),
    .Y(_17135_));
 sky130_fd_sc_hd__a21o_4 _47701_ (.A1(_17026_),
    .A2(_17025_),
    .B1(_17135_),
    .X(_17136_));
 sky130_fd_sc_hd__buf_1 _47702_ (.A(_17026_),
    .X(_17137_));
 sky130_fd_sc_hd__buf_1 _47703_ (.A(_17025_),
    .X(_17138_));
 sky130_fd_sc_hd__nand3_4 _47704_ (.A(_17135_),
    .B(_17137_),
    .C(_17138_),
    .Y(_17139_));
 sky130_fd_sc_hd__nand2_4 _47705_ (.A(_17136_),
    .B(_17139_),
    .Y(_17140_));
 sky130_fd_sc_hd__xor2_4 _47706_ (.A(_17133_),
    .B(_17140_),
    .X(_17141_));
 sky130_fd_sc_hd__a21o_4 _47707_ (.A1(_17131_),
    .A2(_17132_),
    .B1(_17141_),
    .X(_17142_));
 sky130_fd_sc_hd__nand3_4 _47708_ (.A(_17131_),
    .B(_17132_),
    .C(_17141_),
    .Y(_17143_));
 sky130_fd_sc_hd__o21a_4 _47709_ (.A1(_17033_),
    .A2(_17018_),
    .B1(_17020_),
    .X(_17144_));
 sky130_vsdinv _47710_ (.A(_17144_),
    .Y(_17145_));
 sky130_fd_sc_hd__a21o_4 _47711_ (.A1(_17142_),
    .A2(_17143_),
    .B1(_17145_),
    .X(_17146_));
 sky130_fd_sc_hd__nand3_4 _47712_ (.A(_17145_),
    .B(_17142_),
    .C(_17143_),
    .Y(_17147_));
 sky130_fd_sc_hd__buf_1 _47713_ (.A(_16924_),
    .X(_17148_));
 sky130_vsdinv _47714_ (.A(_17022_),
    .Y(_17149_));
 sky130_fd_sc_hd__nand3_4 _47715_ (.A(_17149_),
    .B(_17137_),
    .C(_17138_),
    .Y(_17150_));
 sky130_fd_sc_hd__a21o_4 _47716_ (.A1(_17150_),
    .A2(_17030_),
    .B1(_17042_),
    .X(_17151_));
 sky130_fd_sc_hd__nand3_4 _47717_ (.A(_17030_),
    .B(_17042_),
    .C(_17150_),
    .Y(_17152_));
 sky130_fd_sc_hd__nand2_4 _47718_ (.A(_17151_),
    .B(_17152_),
    .Y(_17153_));
 sky130_fd_sc_hd__xor2_4 _47719_ (.A(_17148_),
    .B(_17153_),
    .X(_17154_));
 sky130_fd_sc_hd__a21o_4 _47720_ (.A1(_17146_),
    .A2(_17147_),
    .B1(_17154_),
    .X(_17155_));
 sky130_fd_sc_hd__nand3_4 _47721_ (.A(_17146_),
    .B(_17147_),
    .C(_17154_),
    .Y(_17156_));
 sky130_fd_sc_hd__nand2_4 _47722_ (.A(_17155_),
    .B(_17156_),
    .Y(_17157_));
 sky130_fd_sc_hd__o21a_4 _47723_ (.A1(_17048_),
    .A2(_17038_),
    .B1(_17040_),
    .X(_17158_));
 sky130_fd_sc_hd__nand2_4 _47724_ (.A(_17157_),
    .B(_17158_),
    .Y(_17159_));
 sky130_vsdinv _47725_ (.A(_17158_),
    .Y(_17160_));
 sky130_fd_sc_hd__nand3_4 _47726_ (.A(_17160_),
    .B(_17155_),
    .C(_17156_),
    .Y(_17161_));
 sky130_fd_sc_hd__buf_8 _47727_ (.A(_16697_),
    .X(_17162_));
 sky130_fd_sc_hd__buf_1 _47728_ (.A(_17057_),
    .X(_17163_));
 sky130_fd_sc_hd__a21o_4 _47729_ (.A1(_17046_),
    .A2(_17043_),
    .B1(_17163_),
    .X(_17164_));
 sky130_fd_sc_hd__nand3_4 _47730_ (.A(_17046_),
    .B(_17163_),
    .C(_17043_),
    .Y(_17165_));
 sky130_fd_sc_hd__nand2_4 _47731_ (.A(_17164_),
    .B(_17165_),
    .Y(_17166_));
 sky130_fd_sc_hd__xor2_4 _47732_ (.A(_17162_),
    .B(_17166_),
    .X(_17167_));
 sky130_fd_sc_hd__a21o_4 _47733_ (.A1(_17159_),
    .A2(_17161_),
    .B1(_17167_),
    .X(_17168_));
 sky130_fd_sc_hd__nand3_4 _47734_ (.A(_17159_),
    .B(_17161_),
    .C(_17167_),
    .Y(_17169_));
 sky130_fd_sc_hd__nand2_4 _47735_ (.A(_17168_),
    .B(_17169_),
    .Y(_17170_));
 sky130_fd_sc_hd__o21a_4 _47736_ (.A1(_17062_),
    .A2(_17053_),
    .B1(_17055_),
    .X(_17171_));
 sky130_fd_sc_hd__nand2_4 _47737_ (.A(_17170_),
    .B(_17171_),
    .Y(_17172_));
 sky130_vsdinv _47738_ (.A(_17171_),
    .Y(_17173_));
 sky130_fd_sc_hd__nand3_4 _47739_ (.A(_17173_),
    .B(_17168_),
    .C(_17169_),
    .Y(_17174_));
 sky130_fd_sc_hd__a21boi_4 _47740_ (.A1(_16829_),
    .A2(_17059_),
    .B1_N(_17058_),
    .Y(_17175_));
 sky130_fd_sc_hd__xor2_4 _47741_ (.A(_16971_),
    .B(_17175_),
    .X(_17176_));
 sky130_fd_sc_hd__xor2_4 _47742_ (.A(_16827_),
    .B(_17176_),
    .X(_17177_));
 sky130_fd_sc_hd__a21oi_4 _47743_ (.A1(_17172_),
    .A2(_17174_),
    .B1(_17177_),
    .Y(_17178_));
 sky130_fd_sc_hd__nand3_4 _47744_ (.A(_17172_),
    .B(_17174_),
    .C(_17177_),
    .Y(_17179_));
 sky130_vsdinv _47745_ (.A(_17179_),
    .Y(_17180_));
 sky130_vsdinv _47746_ (.A(_17069_),
    .Y(_17181_));
 sky130_fd_sc_hd__a21oi_4 _47747_ (.A1(_17068_),
    .A2(_17074_),
    .B1(_17181_),
    .Y(_17182_));
 sky130_fd_sc_hd__o21ai_4 _47748_ (.A1(_17178_),
    .A2(_17180_),
    .B1(_17182_),
    .Y(_17183_));
 sky130_vsdinv _47749_ (.A(_17182_),
    .Y(_17184_));
 sky130_vsdinv _47750_ (.A(_17178_),
    .Y(_17185_));
 sky130_fd_sc_hd__nand3_4 _47751_ (.A(_17184_),
    .B(_17185_),
    .C(_17179_),
    .Y(_17186_));
 sky130_fd_sc_hd__nand2_4 _47752_ (.A(_17183_),
    .B(_17186_),
    .Y(_17187_));
 sky130_fd_sc_hd__a21boi_4 _47753_ (.A1(_17083_),
    .A2(_17072_),
    .B1_N(_17070_),
    .Y(_17188_));
 sky130_fd_sc_hd__xor2_4 _47754_ (.A(_15452_),
    .B(_17188_),
    .X(_17189_));
 sky130_vsdinv _47755_ (.A(_17189_),
    .Y(_17190_));
 sky130_fd_sc_hd__nand2_4 _47756_ (.A(_17187_),
    .B(_17190_),
    .Y(_17191_));
 sky130_fd_sc_hd__nand3_4 _47757_ (.A(_17183_),
    .B(_17186_),
    .C(_17189_),
    .Y(_17192_));
 sky130_fd_sc_hd__nand2_4 _47758_ (.A(_17191_),
    .B(_17192_),
    .Y(_17193_));
 sky130_fd_sc_hd__a21boi_4 _47759_ (.A1(_17079_),
    .A2(_17085_),
    .B1_N(_17081_),
    .Y(_17194_));
 sky130_fd_sc_hd__nand2_4 _47760_ (.A(_17193_),
    .B(_17194_),
    .Y(_17195_));
 sky130_fd_sc_hd__nand2_4 _47761_ (.A(_17088_),
    .B(_17081_),
    .Y(_17196_));
 sky130_fd_sc_hd__nand3_4 _47762_ (.A(_17196_),
    .B(_17191_),
    .C(_17192_),
    .Y(_17197_));
 sky130_fd_sc_hd__nand2_4 _47763_ (.A(_17195_),
    .B(_17197_),
    .Y(_17198_));
 sky130_fd_sc_hd__and2_4 _47764_ (.A(_17084_),
    .B(_17095_),
    .X(_17199_));
 sky130_vsdinv _47765_ (.A(_17199_),
    .Y(_17200_));
 sky130_fd_sc_hd__nand2_4 _47766_ (.A(_17198_),
    .B(_17200_),
    .Y(_17201_));
 sky130_fd_sc_hd__nand3_4 _47767_ (.A(_17195_),
    .B(_17197_),
    .C(_17199_),
    .Y(_17202_));
 sky130_fd_sc_hd__a21oi_4 _47768_ (.A1(_17087_),
    .A2(_17088_),
    .B1(_17090_),
    .Y(_17203_));
 sky130_fd_sc_hd__o21ai_4 _47769_ (.A1(_17097_),
    .A2(_17203_),
    .B1(_17093_),
    .Y(_17204_));
 sky130_fd_sc_hd__a21oi_4 _47770_ (.A1(_17201_),
    .A2(_17202_),
    .B1(_17204_),
    .Y(_17205_));
 sky130_fd_sc_hd__nand3_4 _47771_ (.A(_17204_),
    .B(_17201_),
    .C(_17202_),
    .Y(_17206_));
 sky130_vsdinv _47772_ (.A(_17206_),
    .Y(_17207_));
 sky130_fd_sc_hd__nor2_4 _47773_ (.A(_17205_),
    .B(_17207_),
    .Y(_17208_));
 sky130_fd_sc_hd__a21o_4 _47774_ (.A1(_17098_),
    .A2(_17099_),
    .B1(_17101_),
    .X(_17209_));
 sky130_fd_sc_hd__a21oi_4 _47775_ (.A1(_17110_),
    .A2(_17209_),
    .B1(_17104_),
    .Y(_17210_));
 sky130_fd_sc_hd__xnor2_4 _47776_ (.A(_17208_),
    .B(_17210_),
    .Y(_01464_));
 sky130_fd_sc_hd__maj3_4 _47777_ (.A(_17123_),
    .B(_17124_),
    .C(_17121_),
    .X(_17211_));
 sky130_fd_sc_hd__buf_1 _47778_ (.A(_17028_),
    .X(_17212_));
 sky130_fd_sc_hd__xor2_4 _47779_ (.A(_17211_),
    .B(_17212_),
    .X(_17213_));
 sky130_fd_sc_hd__xor2_4 _47780_ (.A(_17133_),
    .B(_17213_),
    .X(_17214_));
 sky130_fd_sc_hd__a21boi_4 _47781_ (.A1(_17119_),
    .A2(_17126_),
    .B1_N(_17118_),
    .Y(_17215_));
 sky130_vsdinv _47782_ (.A(_17215_),
    .Y(_17216_));
 sky130_vsdinv _47783_ (.A(_17120_),
    .Y(_17217_));
 sky130_fd_sc_hd__nand2_4 _47784_ (.A(_17007_),
    .B(_03617_),
    .Y(_17218_));
 sky130_fd_sc_hd__nand2_4 _47785_ (.A(_16921_),
    .B(_03609_),
    .Y(_17219_));
 sky130_fd_sc_hd__xnor2_4 _47786_ (.A(_17218_),
    .B(_17219_),
    .Y(_17220_));
 sky130_fd_sc_hd__xor2_4 _47787_ (.A(_17217_),
    .B(_17220_),
    .X(_17221_));
 sky130_fd_sc_hd__nand4_4 _47788_ (.A(_17009_),
    .B(_17114_),
    .C(_16996_),
    .D(_17115_),
    .Y(_17222_));
 sky130_fd_sc_hd__and2_4 _47789_ (.A(_17222_),
    .B(_17115_),
    .X(_17223_));
 sky130_fd_sc_hd__a2bb2o_4 _47790_ (.A1_N(_16762_),
    .A2_N(_03636_),
    .B1(_16886_),
    .B2(_17000_),
    .X(_17224_));
 sky130_fd_sc_hd__nand4_4 _47791_ (.A(_03388_),
    .B(_16886_),
    .C(_17000_),
    .D(_11387_),
    .Y(_17225_));
 sky130_fd_sc_hd__nand2_4 _47792_ (.A(_17011_),
    .B(_03623_),
    .Y(_17226_));
 sky130_fd_sc_hd__a21bo_4 _47793_ (.A1(_17224_),
    .A2(_17225_),
    .B1_N(_17226_),
    .X(_17227_));
 sky130_fd_sc_hd__nand4_4 _47794_ (.A(_17122_),
    .B(_17224_),
    .C(_03624_),
    .D(_17225_),
    .Y(_17228_));
 sky130_fd_sc_hd__and2_4 _47795_ (.A(_17227_),
    .B(_17228_),
    .X(_17229_));
 sky130_fd_sc_hd__buf_1 _47796_ (.A(_17229_),
    .X(_17230_));
 sky130_fd_sc_hd__xor2_4 _47797_ (.A(_17223_),
    .B(_17230_),
    .X(_17231_));
 sky130_fd_sc_hd__xor2_4 _47798_ (.A(_17221_),
    .B(_17231_),
    .X(_17232_));
 sky130_fd_sc_hd__xor2_4 _47799_ (.A(_17216_),
    .B(_17232_),
    .X(_17233_));
 sky130_fd_sc_hd__or2_4 _47800_ (.A(_17214_),
    .B(_17233_),
    .X(_17234_));
 sky130_fd_sc_hd__nand2_4 _47801_ (.A(_17233_),
    .B(_17214_),
    .Y(_17235_));
 sky130_fd_sc_hd__a21boi_4 _47802_ (.A1(_17131_),
    .A2(_17141_),
    .B1_N(_17132_),
    .Y(_17236_));
 sky130_vsdinv _47803_ (.A(_17236_),
    .Y(_17237_));
 sky130_fd_sc_hd__a21o_4 _47804_ (.A1(_17234_),
    .A2(_17235_),
    .B1(_17237_),
    .X(_17238_));
 sky130_fd_sc_hd__nand3_4 _47805_ (.A(_17234_),
    .B(_17235_),
    .C(_17237_),
    .Y(_17239_));
 sky130_vsdinv _47806_ (.A(_17133_),
    .Y(_17240_));
 sky130_fd_sc_hd__a21bo_4 _47807_ (.A1(_17136_),
    .A2(_17240_),
    .B1_N(_17139_),
    .X(_17241_));
 sky130_fd_sc_hd__xnor2_4 _47808_ (.A(_17241_),
    .B(_16799_),
    .Y(_17242_));
 sky130_fd_sc_hd__xor2_4 _47809_ (.A(_17148_),
    .B(_17242_),
    .X(_17243_));
 sky130_fd_sc_hd__a21o_4 _47810_ (.A1(_17238_),
    .A2(_17239_),
    .B1(_17243_),
    .X(_17244_));
 sky130_fd_sc_hd__nand3_4 _47811_ (.A(_17238_),
    .B(_17239_),
    .C(_17243_),
    .Y(_17245_));
 sky130_fd_sc_hd__a21boi_4 _47812_ (.A1(_17146_),
    .A2(_17154_),
    .B1_N(_17147_),
    .Y(_17246_));
 sky130_vsdinv _47813_ (.A(_17246_),
    .Y(_17247_));
 sky130_fd_sc_hd__a21o_4 _47814_ (.A1(_17244_),
    .A2(_17245_),
    .B1(_17247_),
    .X(_17248_));
 sky130_fd_sc_hd__nand3_4 _47815_ (.A(_17244_),
    .B(_17245_),
    .C(_17247_),
    .Y(_17249_));
 sky130_fd_sc_hd__buf_1 _47816_ (.A(_16927_),
    .X(_17250_));
 sky130_fd_sc_hd__a21bo_4 _47817_ (.A1(_17250_),
    .A2(_17152_),
    .B1_N(_17151_),
    .X(_17251_));
 sky130_fd_sc_hd__xor2_4 _47818_ (.A(_17163_),
    .B(_17251_),
    .X(_17252_));
 sky130_fd_sc_hd__xor2_4 _47819_ (.A(_17162_),
    .B(_17252_),
    .X(_17253_));
 sky130_fd_sc_hd__a21o_4 _47820_ (.A1(_17248_),
    .A2(_17249_),
    .B1(_17253_),
    .X(_17254_));
 sky130_fd_sc_hd__nand3_4 _47821_ (.A(_17248_),
    .B(_17249_),
    .C(_17253_),
    .Y(_17255_));
 sky130_fd_sc_hd__nand2_4 _47822_ (.A(_17254_),
    .B(_17255_),
    .Y(_17256_));
 sky130_fd_sc_hd__a21o_4 _47823_ (.A1(_17161_),
    .A2(_17169_),
    .B1(_17256_),
    .X(_17257_));
 sky130_fd_sc_hd__nand3_4 _47824_ (.A(_17256_),
    .B(_17161_),
    .C(_17169_),
    .Y(_17258_));
 sky130_fd_sc_hd__nand2_4 _47825_ (.A(_17257_),
    .B(_17258_),
    .Y(_17259_));
 sky130_fd_sc_hd__buf_1 _47826_ (.A(_16829_),
    .X(_17260_));
 sky130_fd_sc_hd__a21boi_4 _47827_ (.A1(_17260_),
    .A2(_17165_),
    .B1_N(_17164_),
    .Y(_17261_));
 sky130_fd_sc_hd__xor2_4 _47828_ (.A(_16971_),
    .B(_17261_),
    .X(_17262_));
 sky130_fd_sc_hd__xor2_4 _47829_ (.A(_16827_),
    .B(_17262_),
    .X(_17263_));
 sky130_vsdinv _47830_ (.A(_17263_),
    .Y(_17264_));
 sky130_fd_sc_hd__nand2_4 _47831_ (.A(_17259_),
    .B(_17264_),
    .Y(_17265_));
 sky130_fd_sc_hd__nand3_4 _47832_ (.A(_17257_),
    .B(_17258_),
    .C(_17263_),
    .Y(_17266_));
 sky130_fd_sc_hd__nand2_4 _47833_ (.A(_17265_),
    .B(_17266_),
    .Y(_17267_));
 sky130_fd_sc_hd__a21boi_4 _47834_ (.A1(_17172_),
    .A2(_17177_),
    .B1_N(_17174_),
    .Y(_17268_));
 sky130_fd_sc_hd__nand2_4 _47835_ (.A(_17267_),
    .B(_17268_),
    .Y(_17269_));
 sky130_vsdinv _47836_ (.A(_17268_),
    .Y(_17270_));
 sky130_fd_sc_hd__nand3_4 _47837_ (.A(_17265_),
    .B(_17266_),
    .C(_17270_),
    .Y(_17271_));
 sky130_fd_sc_hd__nand2_4 _47838_ (.A(_17269_),
    .B(_17271_),
    .Y(_17272_));
 sky130_fd_sc_hd__buf_1 _47839_ (.A(_16827_),
    .X(_17273_));
 sky130_fd_sc_hd__or2_4 _47840_ (.A(_17071_),
    .B(_17175_),
    .X(_17274_));
 sky130_fd_sc_hd__o21ai_4 _47841_ (.A1(_17273_),
    .A2(_17176_),
    .B1(_17274_),
    .Y(_17275_));
 sky130_fd_sc_hd__xor2_4 _47842_ (.A(_16150_),
    .B(_17275_),
    .X(_17276_));
 sky130_vsdinv _47843_ (.A(_17276_),
    .Y(_17277_));
 sky130_fd_sc_hd__nand2_4 _47844_ (.A(_17272_),
    .B(_17277_),
    .Y(_17278_));
 sky130_fd_sc_hd__nand3_4 _47845_ (.A(_17269_),
    .B(_17271_),
    .C(_17276_),
    .Y(_17279_));
 sky130_fd_sc_hd__nand2_4 _47846_ (.A(_17278_),
    .B(_17279_),
    .Y(_17280_));
 sky130_fd_sc_hd__a21boi_4 _47847_ (.A1(_17183_),
    .A2(_17189_),
    .B1_N(_17186_),
    .Y(_17281_));
 sky130_fd_sc_hd__nand2_4 _47848_ (.A(_17280_),
    .B(_17281_),
    .Y(_17282_));
 sky130_vsdinv _47849_ (.A(_17281_),
    .Y(_17283_));
 sky130_fd_sc_hd__nand3_4 _47850_ (.A(_17278_),
    .B(_17279_),
    .C(_17283_),
    .Y(_17284_));
 sky130_fd_sc_hd__nor2_4 _47851_ (.A(_16852_),
    .B(_17188_),
    .Y(_17285_));
 sky130_fd_sc_hd__a21o_4 _47852_ (.A1(_17282_),
    .A2(_17284_),
    .B1(_17285_),
    .X(_17286_));
 sky130_fd_sc_hd__nand3_4 _47853_ (.A(_17282_),
    .B(_17285_),
    .C(_17284_),
    .Y(_17287_));
 sky130_fd_sc_hd__nand2_4 _47854_ (.A(_17286_),
    .B(_17287_),
    .Y(_17288_));
 sky130_fd_sc_hd__a21boi_4 _47855_ (.A1(_17195_),
    .A2(_17199_),
    .B1_N(_17197_),
    .Y(_17289_));
 sky130_fd_sc_hd__nand2_4 _47856_ (.A(_17288_),
    .B(_17289_),
    .Y(_17290_));
 sky130_vsdinv _47857_ (.A(_17289_),
    .Y(_17291_));
 sky130_fd_sc_hd__nand3_4 _47858_ (.A(_17286_),
    .B(_17287_),
    .C(_17291_),
    .Y(_17292_));
 sky130_fd_sc_hd__nand2_4 _47859_ (.A(_17290_),
    .B(_17292_),
    .Y(_17293_));
 sky130_fd_sc_hd__nand4_4 _47860_ (.A(_16860_),
    .B(_17105_),
    .C(_16994_),
    .D(_17208_),
    .Y(_17294_));
 sky130_fd_sc_hd__a21o_4 _47861_ (.A1(_17201_),
    .A2(_17202_),
    .B1(_17204_),
    .X(_17295_));
 sky130_fd_sc_hd__nand4_4 _47862_ (.A(_17103_),
    .B(_17209_),
    .C(_17295_),
    .D(_17206_),
    .Y(_17296_));
 sky130_fd_sc_hd__o21a_4 _47863_ (.A1(_17103_),
    .A2(_17205_),
    .B1(_17206_),
    .X(_17297_));
 sky130_fd_sc_hd__o21a_4 _47864_ (.A1(_17109_),
    .A2(_17296_),
    .B1(_17297_),
    .X(_17298_));
 sky130_fd_sc_hd__o21ai_4 _47865_ (.A1(_17294_),
    .A2(_16872_),
    .B1(_17298_),
    .Y(_17299_));
 sky130_fd_sc_hd__xnor2_4 _47866_ (.A(_17293_),
    .B(_17299_),
    .Y(_01465_));
 sky130_fd_sc_hd__maj3_4 _47867_ (.A(_17121_),
    .B(_17218_),
    .C(_17219_),
    .X(_17300_));
 sky130_fd_sc_hd__xor2_4 _47868_ (.A(_17300_),
    .B(_17212_),
    .X(_17301_));
 sky130_fd_sc_hd__xor2_4 _47869_ (.A(_17133_),
    .B(_17301_),
    .X(_17302_));
 sky130_vsdinv _47870_ (.A(_17223_),
    .Y(_17303_));
 sky130_fd_sc_hd__nand2_4 _47871_ (.A(_17303_),
    .B(_17230_),
    .Y(_17304_));
 sky130_fd_sc_hd__o21ai_4 _47872_ (.A1(_17221_),
    .A2(_17231_),
    .B1(_17304_),
    .Y(_17305_));
 sky130_fd_sc_hd__o21a_4 _47873_ (.A1(_03610_),
    .A2(_03617_),
    .B1(_16921_),
    .X(_17306_));
 sky130_fd_sc_hd__nand3_4 _47874_ (.A(_03410_),
    .B(_03610_),
    .C(_03617_),
    .Y(_17307_));
 sky130_fd_sc_hd__and2_4 _47875_ (.A(_17306_),
    .B(_17307_),
    .X(_17308_));
 sky130_fd_sc_hd__xor2_4 _47876_ (.A(_17121_),
    .B(_17308_),
    .X(_17309_));
 sky130_fd_sc_hd__and2_4 _47877_ (.A(_17228_),
    .B(_17225_),
    .X(_17310_));
 sky130_fd_sc_hd__a2bb2o_4 _47878_ (.A1_N(_17009_),
    .A2_N(_03637_),
    .B1(_17011_),
    .B2(_17113_),
    .X(_17311_));
 sky130_fd_sc_hd__buf_4 _47879_ (.A(_17113_),
    .X(_17312_));
 sky130_fd_sc_hd__nand4_4 _47880_ (.A(_03394_),
    .B(_17122_),
    .C(_17312_),
    .D(_11387_),
    .Y(_17313_));
 sky130_fd_sc_hd__nand2_4 _47881_ (.A(_17007_),
    .B(_16996_),
    .Y(_17314_));
 sky130_fd_sc_hd__a21bo_4 _47882_ (.A1(_17311_),
    .A2(_17313_),
    .B1_N(_17314_),
    .X(_17315_));
 sky130_fd_sc_hd__buf_1 _47883_ (.A(_16543_),
    .X(_17316_));
 sky130_fd_sc_hd__nand4_4 _47884_ (.A(_17316_),
    .B(_17311_),
    .C(_03625_),
    .D(_17313_),
    .Y(_17317_));
 sky130_fd_sc_hd__and2_4 _47885_ (.A(_17315_),
    .B(_17317_),
    .X(_17318_));
 sky130_fd_sc_hd__xnor2_4 _47886_ (.A(_17310_),
    .B(_17318_),
    .Y(_17319_));
 sky130_fd_sc_hd__xnor2_4 _47887_ (.A(_17309_),
    .B(_17319_),
    .Y(_17320_));
 sky130_fd_sc_hd__xor2_4 _47888_ (.A(_17305_),
    .B(_17320_),
    .X(_17321_));
 sky130_fd_sc_hd__or2_4 _47889_ (.A(_17302_),
    .B(_17321_),
    .X(_17322_));
 sky130_fd_sc_hd__nand2_4 _47890_ (.A(_17321_),
    .B(_17302_),
    .Y(_17323_));
 sky130_fd_sc_hd__a21boi_4 _47891_ (.A1(_17232_),
    .A2(_17216_),
    .B1_N(_17235_),
    .Y(_17324_));
 sky130_vsdinv _47892_ (.A(_17324_),
    .Y(_17325_));
 sky130_fd_sc_hd__a21o_4 _47893_ (.A1(_17322_),
    .A2(_17323_),
    .B1(_17325_),
    .X(_17326_));
 sky130_fd_sc_hd__nand3_4 _47894_ (.A(_17325_),
    .B(_17322_),
    .C(_17323_),
    .Y(_17327_));
 sky130_fd_sc_hd__buf_1 _47895_ (.A(_17240_),
    .X(_17328_));
 sky130_vsdinv _47896_ (.A(_17211_),
    .Y(_17329_));
 sky130_fd_sc_hd__maj3_4 _47897_ (.A(_17328_),
    .B(_17212_),
    .C(_17329_),
    .X(_17330_));
 sky130_fd_sc_hd__buf_1 _47898_ (.A(_16799_),
    .X(_17331_));
 sky130_fd_sc_hd__or2_4 _47899_ (.A(_17330_),
    .B(_17331_),
    .X(_17332_));
 sky130_fd_sc_hd__nand2_4 _47900_ (.A(_17331_),
    .B(_17330_),
    .Y(_17333_));
 sky130_fd_sc_hd__nand2_4 _47901_ (.A(_17332_),
    .B(_17333_),
    .Y(_17334_));
 sky130_fd_sc_hd__xor2_4 _47902_ (.A(_17148_),
    .B(_17334_),
    .X(_17335_));
 sky130_fd_sc_hd__a21o_4 _47903_ (.A1(_17326_),
    .A2(_17327_),
    .B1(_17335_),
    .X(_17336_));
 sky130_fd_sc_hd__nand3_4 _47904_ (.A(_17326_),
    .B(_17335_),
    .C(_17327_),
    .Y(_17337_));
 sky130_fd_sc_hd__a21boi_4 _47905_ (.A1(_17238_),
    .A2(_17243_),
    .B1_N(_17239_),
    .Y(_17338_));
 sky130_vsdinv _47906_ (.A(_17338_),
    .Y(_17339_));
 sky130_fd_sc_hd__a21oi_4 _47907_ (.A1(_17336_),
    .A2(_17337_),
    .B1(_17339_),
    .Y(_17340_));
 sky130_fd_sc_hd__nand3_4 _47908_ (.A(_17336_),
    .B(_17339_),
    .C(_17337_),
    .Y(_17341_));
 sky130_vsdinv _47909_ (.A(_17341_),
    .Y(_17342_));
 sky130_vsdinv _47910_ (.A(_17057_),
    .Y(_17343_));
 sky130_fd_sc_hd__maj3_4 _47911_ (.A(_17250_),
    .B(_16799_),
    .C(_17241_),
    .X(_17344_));
 sky130_fd_sc_hd__or2_4 _47912_ (.A(_17343_),
    .B(_17344_),
    .X(_17345_));
 sky130_fd_sc_hd__buf_1 _47913_ (.A(_17345_),
    .X(_17346_));
 sky130_fd_sc_hd__nand2_4 _47914_ (.A(_17344_),
    .B(_17343_),
    .Y(_17347_));
 sky130_fd_sc_hd__a21o_4 _47915_ (.A1(_17346_),
    .A2(_17347_),
    .B1(_17260_),
    .X(_17348_));
 sky130_fd_sc_hd__nand3_4 _47916_ (.A(_17346_),
    .B(_17260_),
    .C(_17347_),
    .Y(_17349_));
 sky130_fd_sc_hd__and2_4 _47917_ (.A(_17348_),
    .B(_17349_),
    .X(_17350_));
 sky130_vsdinv _47918_ (.A(_17350_),
    .Y(_17351_));
 sky130_fd_sc_hd__o21ai_4 _47919_ (.A1(_17340_),
    .A2(_17342_),
    .B1(_17351_),
    .Y(_17352_));
 sky130_vsdinv _47920_ (.A(_17340_),
    .Y(_17353_));
 sky130_fd_sc_hd__nand3_4 _47921_ (.A(_17353_),
    .B(_17341_),
    .C(_17350_),
    .Y(_17354_));
 sky130_fd_sc_hd__a21boi_4 _47922_ (.A1(_17248_),
    .A2(_17253_),
    .B1_N(_17249_),
    .Y(_17355_));
 sky130_vsdinv _47923_ (.A(_17355_),
    .Y(_17356_));
 sky130_fd_sc_hd__a21o_4 _47924_ (.A1(_17352_),
    .A2(_17354_),
    .B1(_17356_),
    .X(_17357_));
 sky130_fd_sc_hd__nand3_4 _47925_ (.A(_17352_),
    .B(_17354_),
    .C(_17356_),
    .Y(_17358_));
 sky130_fd_sc_hd__maj3_4 _47926_ (.A(_17343_),
    .B(_17251_),
    .C(_16829_),
    .X(_17359_));
 sky130_fd_sc_hd__or2_4 _47927_ (.A(_16971_),
    .B(_17359_),
    .X(_17360_));
 sky130_fd_sc_hd__nand2_4 _47928_ (.A(_17359_),
    .B(_16972_),
    .Y(_17361_));
 sky130_fd_sc_hd__a21oi_4 _47929_ (.A1(_17360_),
    .A2(_17361_),
    .B1(_17083_),
    .Y(_17362_));
 sky130_fd_sc_hd__nand3_4 _47930_ (.A(_17360_),
    .B(_17083_),
    .C(_17361_),
    .Y(_17363_));
 sky130_vsdinv _47931_ (.A(_17363_),
    .Y(_17364_));
 sky130_fd_sc_hd__nor2_4 _47932_ (.A(_17362_),
    .B(_17364_),
    .Y(_17365_));
 sky130_fd_sc_hd__a21o_4 _47933_ (.A1(_17357_),
    .A2(_17358_),
    .B1(_17365_),
    .X(_17366_));
 sky130_fd_sc_hd__nand3_4 _47934_ (.A(_17357_),
    .B(_17358_),
    .C(_17365_),
    .Y(_17367_));
 sky130_fd_sc_hd__nand2_4 _47935_ (.A(_17366_),
    .B(_17367_),
    .Y(_17368_));
 sky130_fd_sc_hd__a21boi_4 _47936_ (.A1(_17258_),
    .A2(_17263_),
    .B1_N(_17257_),
    .Y(_17369_));
 sky130_fd_sc_hd__nand2_4 _47937_ (.A(_17368_),
    .B(_17369_),
    .Y(_17370_));
 sky130_vsdinv _47938_ (.A(_17369_),
    .Y(_17371_));
 sky130_fd_sc_hd__nand3_4 _47939_ (.A(_17371_),
    .B(_17367_),
    .C(_17366_),
    .Y(_17372_));
 sky130_fd_sc_hd__nand2_4 _47940_ (.A(_17370_),
    .B(_17372_),
    .Y(_17373_));
 sky130_fd_sc_hd__maj3_4 _47941_ (.A(_17071_),
    .B(_17261_),
    .C(_17273_),
    .X(_17374_));
 sky130_fd_sc_hd__xor2_4 _47942_ (.A(_16314_),
    .B(_17374_),
    .X(_17375_));
 sky130_vsdinv _47943_ (.A(_17375_),
    .Y(_17376_));
 sky130_fd_sc_hd__nand2_4 _47944_ (.A(_17373_),
    .B(_17376_),
    .Y(_17377_));
 sky130_fd_sc_hd__nand3_4 _47945_ (.A(_17370_),
    .B(_17372_),
    .C(_17375_),
    .Y(_17378_));
 sky130_fd_sc_hd__nand2_4 _47946_ (.A(_17377_),
    .B(_17378_),
    .Y(_17379_));
 sky130_fd_sc_hd__a21boi_4 _47947_ (.A1(_17269_),
    .A2(_17276_),
    .B1_N(_17271_),
    .Y(_17380_));
 sky130_fd_sc_hd__nand2_4 _47948_ (.A(_17379_),
    .B(_17380_),
    .Y(_17381_));
 sky130_vsdinv _47949_ (.A(_17380_),
    .Y(_17382_));
 sky130_fd_sc_hd__nand3_4 _47950_ (.A(_17382_),
    .B(_17377_),
    .C(_17378_),
    .Y(_17383_));
 sky130_fd_sc_hd__nand2_4 _47951_ (.A(_17381_),
    .B(_17383_),
    .Y(_17384_));
 sky130_fd_sc_hd__and2_4 _47952_ (.A(_17275_),
    .B(_17095_),
    .X(_17385_));
 sky130_vsdinv _47953_ (.A(_17385_),
    .Y(_17386_));
 sky130_fd_sc_hd__nand2_4 _47954_ (.A(_17384_),
    .B(_17386_),
    .Y(_17387_));
 sky130_fd_sc_hd__nand3_4 _47955_ (.A(_17381_),
    .B(_17385_),
    .C(_17383_),
    .Y(_17388_));
 sky130_fd_sc_hd__nand2_4 _47956_ (.A(_17387_),
    .B(_17388_),
    .Y(_17389_));
 sky130_fd_sc_hd__nand2_4 _47957_ (.A(_17287_),
    .B(_17284_),
    .Y(_17390_));
 sky130_vsdinv _47958_ (.A(_17390_),
    .Y(_17391_));
 sky130_fd_sc_hd__nand2_4 _47959_ (.A(_17389_),
    .B(_17391_),
    .Y(_17392_));
 sky130_fd_sc_hd__nand3_4 _47960_ (.A(_17387_),
    .B(_17390_),
    .C(_17388_),
    .Y(_17393_));
 sky130_fd_sc_hd__nand2_4 _47961_ (.A(_17392_),
    .B(_17393_),
    .Y(_17394_));
 sky130_fd_sc_hd__a21boi_4 _47962_ (.A1(_17299_),
    .A2(_17290_),
    .B1_N(_17292_),
    .Y(_17395_));
 sky130_fd_sc_hd__xor2_4 _47963_ (.A(_17394_),
    .B(_17395_),
    .X(_01466_));
 sky130_fd_sc_hd__a21boi_4 _47964_ (.A1(_17320_),
    .A2(_17305_),
    .B1_N(_17323_),
    .Y(_17396_));
 sky130_vsdinv _47965_ (.A(_17396_),
    .Y(_17397_));
 sky130_fd_sc_hd__a21bo_4 _47966_ (.A1(_17306_),
    .A2(_17217_),
    .B1_N(_17307_),
    .X(_17398_));
 sky130_fd_sc_hd__a21o_4 _47967_ (.A1(_17138_),
    .A2(_17137_),
    .B1(_17398_),
    .X(_17399_));
 sky130_fd_sc_hd__nand3_4 _47968_ (.A(_17398_),
    .B(_17138_),
    .C(_17137_),
    .Y(_17400_));
 sky130_fd_sc_hd__and2_4 _47969_ (.A(_17399_),
    .B(_17400_),
    .X(_17401_));
 sky130_fd_sc_hd__xor2_4 _47970_ (.A(_17328_),
    .B(_17401_),
    .X(_17402_));
 sky130_vsdinv _47971_ (.A(_17318_),
    .Y(_17403_));
 sky130_fd_sc_hd__buf_8 _47972_ (.A(_17309_),
    .X(_17404_));
 sky130_fd_sc_hd__maj3_4 _47973_ (.A(_17310_),
    .B(_17403_),
    .C(_17404_),
    .X(_17405_));
 sky130_fd_sc_hd__and2_4 _47974_ (.A(_17317_),
    .B(_17313_),
    .X(_17406_));
 sky130_fd_sc_hd__buf_1 _47975_ (.A(_17406_),
    .X(_17407_));
 sky130_fd_sc_hd__nand2_4 _47976_ (.A(_03410_),
    .B(_03625_),
    .Y(_17408_));
 sky130_fd_sc_hd__a2bb2o_4 _47977_ (.A1_N(_17122_),
    .A2_N(_03637_),
    .B1(_17316_),
    .B2(_17312_),
    .X(_17409_));
 sky130_fd_sc_hd__nand4_4 _47978_ (.A(_03398_),
    .B(_17316_),
    .C(_17312_),
    .D(_11388_),
    .Y(_17410_));
 sky130_fd_sc_hd__and2_4 _47979_ (.A(_17409_),
    .B(_17410_),
    .X(_17411_));
 sky130_fd_sc_hd__xor2_4 _47980_ (.A(_17408_),
    .B(_17411_),
    .X(_17412_));
 sky130_fd_sc_hd__xnor2_4 _47981_ (.A(_17407_),
    .B(_17412_),
    .Y(_17413_));
 sky130_fd_sc_hd__xnor2_4 _47982_ (.A(_17404_),
    .B(_17413_),
    .Y(_17414_));
 sky130_fd_sc_hd__xor2_4 _47983_ (.A(_17405_),
    .B(_17414_),
    .X(_17415_));
 sky130_fd_sc_hd__xor2_4 _47984_ (.A(_17402_),
    .B(_17415_),
    .X(_17416_));
 sky130_fd_sc_hd__or2_4 _47985_ (.A(_17397_),
    .B(_17416_),
    .X(_17417_));
 sky130_fd_sc_hd__buf_1 _47986_ (.A(_17417_),
    .X(_17418_));
 sky130_fd_sc_hd__nand2_4 _47987_ (.A(_17416_),
    .B(_17397_),
    .Y(_17419_));
 sky130_vsdinv _47988_ (.A(_17300_),
    .Y(_17420_));
 sky130_fd_sc_hd__maj3_4 _47989_ (.A(_17328_),
    .B(_17212_),
    .C(_17420_),
    .X(_17421_));
 sky130_fd_sc_hd__xnor2_4 _47990_ (.A(_17421_),
    .B(_17331_),
    .Y(_17422_));
 sky130_fd_sc_hd__xor2_4 _47991_ (.A(_17148_),
    .B(_17422_),
    .X(_17423_));
 sky130_fd_sc_hd__a21o_4 _47992_ (.A1(_17418_),
    .A2(_17419_),
    .B1(_17423_),
    .X(_17424_));
 sky130_fd_sc_hd__nand3_4 _47993_ (.A(_17418_),
    .B(_17419_),
    .C(_17423_),
    .Y(_17425_));
 sky130_fd_sc_hd__a21boi_4 _47994_ (.A1(_17326_),
    .A2(_17335_),
    .B1_N(_17327_),
    .Y(_17426_));
 sky130_vsdinv _47995_ (.A(_17426_),
    .Y(_17427_));
 sky130_fd_sc_hd__a21o_4 _47996_ (.A1(_17424_),
    .A2(_17425_),
    .B1(_17427_),
    .X(_17428_));
 sky130_fd_sc_hd__nand3_4 _47997_ (.A(_17427_),
    .B(_17424_),
    .C(_17425_),
    .Y(_17429_));
 sky130_fd_sc_hd__a21boi_4 _47998_ (.A1(_17332_),
    .A2(_17250_),
    .B1_N(_17333_),
    .Y(_17430_));
 sky130_fd_sc_hd__xor2_4 _47999_ (.A(_17343_),
    .B(_17430_),
    .X(_17431_));
 sky130_fd_sc_hd__xor2_4 _48000_ (.A(_17162_),
    .B(_17431_),
    .X(_17432_));
 sky130_fd_sc_hd__a21o_4 _48001_ (.A1(_17428_),
    .A2(_17429_),
    .B1(_17432_),
    .X(_17433_));
 sky130_fd_sc_hd__nand3_4 _48002_ (.A(_17428_),
    .B(_17429_),
    .C(_17432_),
    .Y(_17434_));
 sky130_fd_sc_hd__o21a_4 _48003_ (.A1(_17351_),
    .A2(_17340_),
    .B1(_17341_),
    .X(_17435_));
 sky130_vsdinv _48004_ (.A(_17435_),
    .Y(_17436_));
 sky130_fd_sc_hd__a21o_4 _48005_ (.A1(_17433_),
    .A2(_17434_),
    .B1(_17436_),
    .X(_17437_));
 sky130_fd_sc_hd__nand3_4 _48006_ (.A(_17436_),
    .B(_17433_),
    .C(_17434_),
    .Y(_17438_));
 sky130_fd_sc_hd__a21boi_4 _48007_ (.A1(_17346_),
    .A2(_17260_),
    .B1_N(_17347_),
    .Y(_17439_));
 sky130_fd_sc_hd__xor2_4 _48008_ (.A(_16972_),
    .B(_17439_),
    .X(_17440_));
 sky130_fd_sc_hd__xor2_4 _48009_ (.A(_17273_),
    .B(_17440_),
    .X(_17441_));
 sky130_fd_sc_hd__a21o_4 _48010_ (.A1(_17437_),
    .A2(_17438_),
    .B1(_17441_),
    .X(_17442_));
 sky130_fd_sc_hd__nand3_4 _48011_ (.A(_17437_),
    .B(_17438_),
    .C(_17441_),
    .Y(_17443_));
 sky130_fd_sc_hd__a21boi_4 _48012_ (.A1(_17357_),
    .A2(_17365_),
    .B1_N(_17358_),
    .Y(_17444_));
 sky130_vsdinv _48013_ (.A(_17444_),
    .Y(_17445_));
 sky130_fd_sc_hd__a21o_4 _48014_ (.A1(_17442_),
    .A2(_17443_),
    .B1(_17445_),
    .X(_17446_));
 sky130_fd_sc_hd__nand3_4 _48015_ (.A(_17442_),
    .B(_17443_),
    .C(_17445_),
    .Y(_17447_));
 sky130_fd_sc_hd__a21oi_4 _48016_ (.A1(_17363_),
    .A2(_17361_),
    .B1(_17095_),
    .Y(_17448_));
 sky130_fd_sc_hd__and3_4 _48017_ (.A(_17363_),
    .B(_16150_),
    .C(_17361_),
    .X(_17449_));
 sky130_fd_sc_hd__nor2_4 _48018_ (.A(_17448_),
    .B(_17449_),
    .Y(_17450_));
 sky130_vsdinv _48019_ (.A(_17450_),
    .Y(_17451_));
 sky130_fd_sc_hd__a21o_4 _48020_ (.A1(_17446_),
    .A2(_17447_),
    .B1(_17451_),
    .X(_17452_));
 sky130_fd_sc_hd__nand3_4 _48021_ (.A(_17446_),
    .B(_17447_),
    .C(_17451_),
    .Y(_17453_));
 sky130_fd_sc_hd__a21boi_4 _48022_ (.A1(_17370_),
    .A2(_17375_),
    .B1_N(_17372_),
    .Y(_17454_));
 sky130_vsdinv _48023_ (.A(_17454_),
    .Y(_17455_));
 sky130_fd_sc_hd__a21oi_4 _48024_ (.A1(_17452_),
    .A2(_17453_),
    .B1(_17455_),
    .Y(_17456_));
 sky130_vsdinv _48025_ (.A(_17456_),
    .Y(_17457_));
 sky130_fd_sc_hd__nand3_4 _48026_ (.A(_17452_),
    .B(_17455_),
    .C(_17453_),
    .Y(_17458_));
 sky130_fd_sc_hd__nor2_4 _48027_ (.A(_16852_),
    .B(_17374_),
    .Y(_17459_));
 sky130_fd_sc_hd__a21o_4 _48028_ (.A1(_17457_),
    .A2(_17458_),
    .B1(_17459_),
    .X(_17460_));
 sky130_fd_sc_hd__nand3_4 _48029_ (.A(_17457_),
    .B(_17459_),
    .C(_17458_),
    .Y(_17461_));
 sky130_fd_sc_hd__nand2_4 _48030_ (.A(_17460_),
    .B(_17461_),
    .Y(_17462_));
 sky130_fd_sc_hd__a21boi_4 _48031_ (.A1(_17381_),
    .A2(_17385_),
    .B1_N(_17383_),
    .Y(_17463_));
 sky130_fd_sc_hd__nand2_4 _48032_ (.A(_17462_),
    .B(_17463_),
    .Y(_17464_));
 sky130_vsdinv _48033_ (.A(_17463_),
    .Y(_17465_));
 sky130_fd_sc_hd__nand3_4 _48034_ (.A(_17460_),
    .B(_17465_),
    .C(_17461_),
    .Y(_17466_));
 sky130_fd_sc_hd__nand2_4 _48035_ (.A(_17464_),
    .B(_17466_),
    .Y(_17467_));
 sky130_fd_sc_hd__nor2_4 _48036_ (.A(_17293_),
    .B(_17394_),
    .Y(_17468_));
 sky130_fd_sc_hd__nand2_4 _48037_ (.A(_17299_),
    .B(_17468_),
    .Y(_17469_));
 sky130_fd_sc_hd__maj3_4 _48038_ (.A(_17292_),
    .B(_17389_),
    .C(_17391_),
    .X(_17470_));
 sky130_fd_sc_hd__nand2_4 _48039_ (.A(_17469_),
    .B(_17470_),
    .Y(_17471_));
 sky130_fd_sc_hd__xnor2_4 _48040_ (.A(_17467_),
    .B(_17471_),
    .Y(_01467_));
 sky130_vsdinv _48041_ (.A(_17467_),
    .Y(_17472_));
 sky130_fd_sc_hd__nand2_4 _48042_ (.A(_17471_),
    .B(_17472_),
    .Y(_17473_));
 sky130_fd_sc_hd__maj3_4 _48043_ (.A(_17071_),
    .B(_17439_),
    .C(_17273_),
    .X(_17474_));
 sky130_vsdinv _48044_ (.A(_17474_),
    .Y(_17475_));
 sky130_fd_sc_hd__a21o_4 _48045_ (.A1(_17453_),
    .A2(_17447_),
    .B1(_17475_),
    .X(_17476_));
 sky130_fd_sc_hd__nand3_4 _48046_ (.A(_17453_),
    .B(_17447_),
    .C(_17475_),
    .Y(_17477_));
 sky130_fd_sc_hd__nand2_4 _48047_ (.A(_14757_),
    .B(_15781_),
    .Y(_17478_));
 sky130_fd_sc_hd__a21boi_4 _48048_ (.A1(_13480_),
    .A2(_15783_),
    .B1_N(_17478_),
    .Y(_17479_));
 sky130_vsdinv _48049_ (.A(_17479_),
    .Y(_17480_));
 sky130_fd_sc_hd__a21o_4 _48050_ (.A1(_17476_),
    .A2(_17477_),
    .B1(_17480_),
    .X(_17481_));
 sky130_fd_sc_hd__nand3_4 _48051_ (.A(_17476_),
    .B(_17477_),
    .C(_17480_),
    .Y(_17482_));
 sky130_vsdinv _48052_ (.A(_17449_),
    .Y(_17483_));
 sky130_fd_sc_hd__a21o_4 _48053_ (.A1(_17481_),
    .A2(_17482_),
    .B1(_17483_),
    .X(_17484_));
 sky130_fd_sc_hd__nand3_4 _48054_ (.A(_17481_),
    .B(_17483_),
    .C(_17482_),
    .Y(_17485_));
 sky130_fd_sc_hd__a21boi_4 _48055_ (.A1(_15376_),
    .A2(_15377_),
    .B1_N(_16567_),
    .Y(_17486_));
 sky130_fd_sc_hd__a21oi_4 _48056_ (.A1(_16266_),
    .A2(_16566_),
    .B1(_17486_),
    .Y(_17487_));
 sky130_fd_sc_hd__maj3_4 _48057_ (.A(_17163_),
    .B(_17430_),
    .C(_17162_),
    .X(_17488_));
 sky130_fd_sc_hd__xor2_4 _48058_ (.A(_17487_),
    .B(_17488_),
    .X(_17489_));
 sky130_fd_sc_hd__nand2_4 _48059_ (.A(_16680_),
    .B(_16922_),
    .Y(_17490_));
 sky130_fd_sc_hd__o21ai_4 _48060_ (.A1(_16923_),
    .A2(_16680_),
    .B1(_17490_),
    .Y(_17491_));
 sky130_fd_sc_hd__maj3_4 _48061_ (.A(_17250_),
    .B(_17331_),
    .C(_17421_),
    .X(_17492_));
 sky130_fd_sc_hd__xor2_4 _48062_ (.A(_17491_),
    .B(_17492_),
    .X(_17493_));
 sky130_vsdinv _48063_ (.A(_17408_),
    .Y(_17494_));
 sky130_fd_sc_hd__a21boi_4 _48064_ (.A1(_17409_),
    .A2(_17494_),
    .B1_N(_17410_),
    .Y(_17495_));
 sky130_fd_sc_hd__or2_4 _48065_ (.A(_17405_),
    .B(_17414_),
    .X(_17496_));
 sky130_fd_sc_hd__a21bo_4 _48066_ (.A1(_17415_),
    .A2(_17402_),
    .B1_N(_17496_),
    .X(_17497_));
 sky130_fd_sc_hd__or2_4 _48067_ (.A(_17495_),
    .B(_17497_),
    .X(_17498_));
 sky130_fd_sc_hd__nand2_4 _48068_ (.A(_17497_),
    .B(_17495_),
    .Y(_17499_));
 sky130_fd_sc_hd__a21boi_4 _48069_ (.A1(_17399_),
    .A2(_17328_),
    .B1_N(_17400_),
    .Y(_17500_));
 sky130_vsdinv _48070_ (.A(_17500_),
    .Y(_17501_));
 sky130_fd_sc_hd__a21o_4 _48071_ (.A1(_17498_),
    .A2(_17499_),
    .B1(_17501_),
    .X(_17502_));
 sky130_fd_sc_hd__nand3_4 _48072_ (.A(_17498_),
    .B(_17501_),
    .C(_17499_),
    .Y(_17503_));
 sky130_fd_sc_hd__nand2_4 _48073_ (.A(_03410_),
    .B(_17312_),
    .Y(_17504_));
 sky130_fd_sc_hd__maj3_4 _48074_ (.A(_17404_),
    .B(_17412_),
    .C(_17407_),
    .X(_17505_));
 sky130_fd_sc_hd__xnor2_4 _48075_ (.A(_17504_),
    .B(_17505_),
    .Y(_17506_));
 sky130_fd_sc_hd__xor2_4 _48076_ (.A(_17494_),
    .B(_17404_),
    .X(_17507_));
 sky130_fd_sc_hd__nor2_4 _48077_ (.A(_17316_),
    .B(_03637_),
    .Y(_17508_));
 sky130_fd_sc_hd__xor2_4 _48078_ (.A(_17508_),
    .B(_17402_),
    .X(_17509_));
 sky130_fd_sc_hd__xor2_4 _48079_ (.A(_17507_),
    .B(_17509_),
    .X(_17510_));
 sky130_fd_sc_hd__xnor2_4 _48080_ (.A(_17506_),
    .B(_17510_),
    .Y(_17511_));
 sky130_fd_sc_hd__a21o_4 _48081_ (.A1(_17502_),
    .A2(_17503_),
    .B1(_17511_),
    .X(_17512_));
 sky130_fd_sc_hd__nand3_4 _48082_ (.A(_17502_),
    .B(_17511_),
    .C(_17503_),
    .Y(_17513_));
 sky130_fd_sc_hd__a21boi_4 _48083_ (.A1(_17418_),
    .A2(_17423_),
    .B1_N(_17419_),
    .Y(_17514_));
 sky130_vsdinv _48084_ (.A(_17514_),
    .Y(_17515_));
 sky130_fd_sc_hd__a21o_4 _48085_ (.A1(_17512_),
    .A2(_17513_),
    .B1(_17515_),
    .X(_17516_));
 sky130_fd_sc_hd__nand3_4 _48086_ (.A(_17512_),
    .B(_17515_),
    .C(_17513_),
    .Y(_17517_));
 sky130_fd_sc_hd__nand2_4 _48087_ (.A(_17516_),
    .B(_17517_),
    .Y(_17518_));
 sky130_fd_sc_hd__or2_4 _48088_ (.A(_17493_),
    .B(_17518_),
    .X(_17519_));
 sky130_fd_sc_hd__nand2_4 _48089_ (.A(_17518_),
    .B(_17493_),
    .Y(_17520_));
 sky130_fd_sc_hd__a21boi_4 _48090_ (.A1(_17428_),
    .A2(_17432_),
    .B1_N(_17429_),
    .Y(_17521_));
 sky130_vsdinv _48091_ (.A(_17521_),
    .Y(_17522_));
 sky130_fd_sc_hd__a21o_4 _48092_ (.A1(_17519_),
    .A2(_17520_),
    .B1(_17522_),
    .X(_17523_));
 sky130_fd_sc_hd__nand3_4 _48093_ (.A(_17519_),
    .B(_17522_),
    .C(_17520_),
    .Y(_17524_));
 sky130_fd_sc_hd__nand2_4 _48094_ (.A(_17523_),
    .B(_17524_),
    .Y(_17525_));
 sky130_fd_sc_hd__or2_4 _48095_ (.A(_17489_),
    .B(_17525_),
    .X(_17526_));
 sky130_fd_sc_hd__nand2_4 _48096_ (.A(_17525_),
    .B(_17489_),
    .Y(_17527_));
 sky130_fd_sc_hd__a21boi_4 _48097_ (.A1(_17437_),
    .A2(_17441_),
    .B1_N(_17438_),
    .Y(_17528_));
 sky130_vsdinv _48098_ (.A(_17528_),
    .Y(_17529_));
 sky130_fd_sc_hd__a21o_4 _48099_ (.A1(_17526_),
    .A2(_17527_),
    .B1(_17529_),
    .X(_17530_));
 sky130_fd_sc_hd__nand3_4 _48100_ (.A(_17526_),
    .B(_17529_),
    .C(_17527_),
    .Y(_17531_));
 sky130_fd_sc_hd__and2_4 _48101_ (.A(_17530_),
    .B(_17531_),
    .X(_17532_));
 sky130_vsdinv _48102_ (.A(_17532_),
    .Y(_17533_));
 sky130_fd_sc_hd__nand3_4 _48103_ (.A(_17461_),
    .B(_17458_),
    .C(_17533_),
    .Y(_17534_));
 sky130_vsdinv _48104_ (.A(_17459_),
    .Y(_17535_));
 sky130_fd_sc_hd__o21ai_4 _48105_ (.A1(_17535_),
    .A2(_17456_),
    .B1(_17458_),
    .Y(_17536_));
 sky130_fd_sc_hd__nand2_4 _48106_ (.A(_17536_),
    .B(_17532_),
    .Y(_17537_));
 sky130_fd_sc_hd__nand2_4 _48107_ (.A(_17534_),
    .B(_17537_),
    .Y(_17538_));
 sky130_fd_sc_hd__a21o_4 _48108_ (.A1(_17484_),
    .A2(_17485_),
    .B1(_17538_),
    .X(_17539_));
 sky130_fd_sc_hd__nand3_4 _48109_ (.A(_17538_),
    .B(_17484_),
    .C(_17485_),
    .Y(_17540_));
 sky130_fd_sc_hd__nand2_4 _48110_ (.A(_17539_),
    .B(_17540_),
    .Y(_17541_));
 sky130_vsdinv _48111_ (.A(_17541_),
    .Y(_17542_));
 sky130_fd_sc_hd__a21oi_4 _48112_ (.A1(_17473_),
    .A2(_17466_),
    .B1(_17542_),
    .Y(_17543_));
 sky130_vsdinv _48113_ (.A(_17466_),
    .Y(_17544_));
 sky130_fd_sc_hd__a21oi_4 _48114_ (.A1(_17469_),
    .A2(_17470_),
    .B1(_17467_),
    .Y(_17545_));
 sky130_fd_sc_hd__nor3_4 _48115_ (.A(_17544_),
    .B(_17541_),
    .C(_17545_),
    .Y(_17546_));
 sky130_fd_sc_hd__nor2_4 _48116_ (.A(_17543_),
    .B(_17546_),
    .Y(_01468_));
 sky130_fd_sc_hd__a21oi_4 _48117_ (.A1(_06046_),
    .A2(_06048_),
    .B1(_05986_),
    .Y(_17547_));
 sky130_fd_sc_hd__nor2_4 _48118_ (.A(_17547_),
    .B(_06122_),
    .Y(_01414_));
 sky130_fd_sc_hd__buf_1 _48119_ (.A(_03467_),
    .X(_17548_));
 sky130_fd_sc_hd__buf_1 _48120_ (.A(_17548_),
    .X(_17549_));
 sky130_fd_sc_hd__nor3_4 _48121_ (.A(_21344_),
    .B(_17549_),
    .C(_05616_),
    .Y(_24285_));
 sky130_fd_sc_hd__nor2_4 _48122_ (.A(_03428_),
    .B(_03697_),
    .Y(_17550_));
 sky130_fd_sc_hd__o21a_4 _48123_ (.A1(_04546_),
    .A2(_17550_),
    .B1(_21127_),
    .X(_17551_));
 sky130_fd_sc_hd__buf_1 _48124_ (.A(_21153_),
    .X(_17552_));
 sky130_fd_sc_hd__buf_1 _48125_ (.A(_17552_),
    .X(_17553_));
 sky130_fd_sc_hd__buf_1 _48126_ (.A(_17553_),
    .X(_17554_));
 sky130_fd_sc_hd__buf_1 _48127_ (.A(_21168_),
    .X(_17555_));
 sky130_fd_sc_hd__and4_4 _48128_ (.A(_17551_),
    .B(_17554_),
    .C(_21145_),
    .D(_17555_),
    .X(_24296_));
 sky130_fd_sc_hd__buf_1 _48129_ (.A(_18608_),
    .X(_17556_));
 sky130_fd_sc_hd__buf_1 _48130_ (.A(_17556_),
    .X(_17557_));
 sky130_fd_sc_hd__buf_1 _48131_ (.A(_17557_),
    .X(_17558_));
 sky130_fd_sc_hd__buf_1 _48132_ (.A(_18629_),
    .X(_17559_));
 sky130_fd_sc_hd__buf_1 _48133_ (.A(_03424_),
    .X(_17560_));
 sky130_fd_sc_hd__nand2_4 _48134_ (.A(_18619_),
    .B(_17560_),
    .Y(_17561_));
 sky130_fd_sc_hd__o21a_4 _48135_ (.A1(_17559_),
    .A2(_21389_),
    .B1(_17561_),
    .X(_17562_));
 sky130_fd_sc_hd__buf_1 _48136_ (.A(_21122_),
    .X(_17563_));
 sky130_fd_sc_hd__buf_1 _48137_ (.A(_17563_),
    .X(_17564_));
 sky130_fd_sc_hd__a21bo_4 _48138_ (.A1(_17562_),
    .A2(_17564_),
    .B1_N(_05440_),
    .X(_17565_));
 sky130_fd_sc_hd__nor4_4 _48139_ (.A(_17558_),
    .B(_03450_),
    .C(_17549_),
    .D(_17565_),
    .Y(_24307_));
 sky130_fd_sc_hd__buf_1 _48140_ (.A(_18622_),
    .X(_17566_));
 sky130_fd_sc_hd__buf_1 _48141_ (.A(_17566_),
    .X(_17567_));
 sky130_fd_sc_hd__buf_1 _48142_ (.A(_03424_),
    .X(_17568_));
 sky130_fd_sc_hd__buf_1 _48143_ (.A(_17568_),
    .X(_17569_));
 sky130_fd_sc_hd__buf_1 _48144_ (.A(_17569_),
    .X(_17570_));
 sky130_fd_sc_hd__o21ai_4 _48145_ (.A1(_17570_),
    .A2(_21367_),
    .B1(_18633_),
    .Y(_17571_));
 sky130_fd_sc_hd__buf_1 _48146_ (.A(_18629_),
    .X(_17572_));
 sky130_fd_sc_hd__nand2_4 _48147_ (.A(_17572_),
    .B(_21397_),
    .Y(_17573_));
 sky130_vsdinv _48148_ (.A(_17573_),
    .Y(_17574_));
 sky130_fd_sc_hd__buf_1 _48149_ (.A(_03424_),
    .X(_17575_));
 sky130_fd_sc_hd__buf_1 _48150_ (.A(_17575_),
    .X(_17576_));
 sky130_fd_sc_hd__nor2_4 _48151_ (.A(_17576_),
    .B(_21409_),
    .Y(_17577_));
 sky130_fd_sc_hd__buf_1 _48152_ (.A(_21122_),
    .X(_17578_));
 sky130_fd_sc_hd__buf_1 _48153_ (.A(_17578_),
    .X(_17579_));
 sky130_fd_sc_hd__o21a_4 _48154_ (.A1(_17574_),
    .A2(_17577_),
    .B1(_17579_),
    .X(_17580_));
 sky130_fd_sc_hd__a21o_4 _48155_ (.A1(_17567_),
    .A2(_17571_),
    .B1(_17580_),
    .X(_17581_));
 sky130_fd_sc_hd__and4_4 _48156_ (.A(_17581_),
    .B(_17554_),
    .C(_21145_),
    .D(_01521_),
    .X(_24310_));
 sky130_fd_sc_hd__buf_1 _48157_ (.A(_17560_),
    .X(_17582_));
 sky130_fd_sc_hd__buf_1 _48158_ (.A(_17582_),
    .X(_17583_));
 sky130_fd_sc_hd__buf_1 _48159_ (.A(_17572_),
    .X(_17584_));
 sky130_fd_sc_hd__nand2_4 _48160_ (.A(_17584_),
    .B(_21408_),
    .Y(_17585_));
 sky130_fd_sc_hd__o21ai_4 _48161_ (.A1(_17583_),
    .A2(_21435_),
    .B1(_17585_),
    .Y(_17586_));
 sky130_fd_sc_hd__buf_1 _48162_ (.A(_17564_),
    .X(_17587_));
 sky130_fd_sc_hd__nand2_4 _48163_ (.A(_17586_),
    .B(_17587_),
    .Y(_17588_));
 sky130_fd_sc_hd__o21ai_4 _48164_ (.A1(_21125_),
    .A2(_17562_),
    .B1(_17588_),
    .Y(_17589_));
 sky130_fd_sc_hd__buf_1 _48165_ (.A(_21140_),
    .X(_17590_));
 sky130_fd_sc_hd__buf_1 _48166_ (.A(_17590_),
    .X(_17591_));
 sky130_fd_sc_hd__buf_1 _48167_ (.A(_03446_),
    .X(_17592_));
 sky130_fd_sc_hd__nand4_4 _48168_ (.A(_18300_),
    .B(_21109_),
    .C(_21125_),
    .D(_17592_),
    .Y(_17593_));
 sky130_fd_sc_hd__a21bo_4 _48169_ (.A1(_17589_),
    .A2(_17591_),
    .B1_N(_17593_),
    .X(_17594_));
 sky130_fd_sc_hd__buf_1 _48170_ (.A(_21168_),
    .X(_17595_));
 sky130_fd_sc_hd__and3_4 _48171_ (.A(_17594_),
    .B(_21156_),
    .C(_17595_),
    .X(_24311_));
 sky130_fd_sc_hd__nand2_4 _48172_ (.A(_17584_),
    .B(_21434_),
    .Y(_17596_));
 sky130_fd_sc_hd__o21ai_4 _48173_ (.A1(_17583_),
    .A2(_21455_),
    .B1(_17596_),
    .Y(_17597_));
 sky130_fd_sc_hd__o21a_4 _48174_ (.A1(_17574_),
    .A2(_17577_),
    .B1(_17566_),
    .X(_17598_));
 sky130_fd_sc_hd__a21o_4 _48175_ (.A1(_17587_),
    .A2(_17597_),
    .B1(_17598_),
    .X(_17599_));
 sky130_fd_sc_hd__buf_1 _48176_ (.A(_17578_),
    .X(_17600_));
 sky130_fd_sc_hd__buf_1 _48177_ (.A(_17600_),
    .X(_17601_));
 sky130_fd_sc_hd__nand3_4 _48178_ (.A(_17571_),
    .B(_17601_),
    .C(_17592_),
    .Y(_17602_));
 sky130_fd_sc_hd__a21bo_4 _48179_ (.A1(_17599_),
    .A2(_17591_),
    .B1_N(_17602_),
    .X(_17603_));
 sky130_fd_sc_hd__and3_4 _48180_ (.A(_17603_),
    .B(_17554_),
    .C(_17555_),
    .X(_24312_));
 sky130_fd_sc_hd__buf_1 _48181_ (.A(_18622_),
    .X(_17604_));
 sky130_fd_sc_hd__buf_1 _48182_ (.A(_17604_),
    .X(_17605_));
 sky130_fd_sc_hd__nand2_4 _48183_ (.A(_17559_),
    .B(_18582_),
    .Y(_17606_));
 sky130_vsdinv _48184_ (.A(_17606_),
    .Y(_17607_));
 sky130_fd_sc_hd__buf_1 _48185_ (.A(_17575_),
    .X(_17608_));
 sky130_fd_sc_hd__nor2_4 _48186_ (.A(_17608_),
    .B(_21471_),
    .Y(_17609_));
 sky130_fd_sc_hd__o21a_4 _48187_ (.A1(_17607_),
    .A2(_17609_),
    .B1(_17579_),
    .X(_17610_));
 sky130_fd_sc_hd__a21o_4 _48188_ (.A1(_17605_),
    .A2(_17586_),
    .B1(_17610_),
    .X(_17611_));
 sky130_fd_sc_hd__or2_4 _48189_ (.A(_21141_),
    .B(_17565_),
    .X(_17612_));
 sky130_fd_sc_hd__a21bo_4 _48190_ (.A1(_24246_),
    .A2(_17611_),
    .B1_N(_17612_),
    .X(_17613_));
 sky130_fd_sc_hd__and3_4 _48191_ (.A(_17613_),
    .B(_17554_),
    .C(_17555_),
    .X(_24313_));
 sky130_fd_sc_hd__buf_1 _48192_ (.A(_17591_),
    .X(_17614_));
 sky130_fd_sc_hd__nand2_4 _48193_ (.A(_18630_),
    .B(_21479_),
    .Y(_17615_));
 sky130_vsdinv _48194_ (.A(_17615_),
    .Y(_17616_));
 sky130_fd_sc_hd__buf_1 _48195_ (.A(_17560_),
    .X(_17617_));
 sky130_fd_sc_hd__nor2_4 _48196_ (.A(_17617_),
    .B(_21486_),
    .Y(_17618_));
 sky130_fd_sc_hd__o21a_4 _48197_ (.A1(_17616_),
    .A2(_17618_),
    .B1(_17579_),
    .X(_17619_));
 sky130_fd_sc_hd__a21o_4 _48198_ (.A1(_17567_),
    .A2(_17597_),
    .B1(_17619_),
    .X(_17620_));
 sky130_fd_sc_hd__buf_1 _48199_ (.A(_03447_),
    .X(_17621_));
 sky130_fd_sc_hd__and2_4 _48200_ (.A(_17581_),
    .B(_17621_),
    .X(_17622_));
 sky130_fd_sc_hd__a21o_4 _48201_ (.A1(_17614_),
    .A2(_17620_),
    .B1(_17622_),
    .X(_17623_));
 sky130_fd_sc_hd__nand3_4 _48202_ (.A(_17623_),
    .B(_01518_),
    .C(_01521_),
    .Y(_17624_));
 sky130_vsdinv _48203_ (.A(_17624_),
    .Y(_24314_));
 sky130_fd_sc_hd__buf_1 _48204_ (.A(_03458_),
    .X(_17625_));
 sky130_fd_sc_hd__buf_1 _48205_ (.A(_03446_),
    .X(_17626_));
 sky130_fd_sc_hd__buf_1 _48206_ (.A(_17626_),
    .X(_17627_));
 sky130_fd_sc_hd__buf_1 _48207_ (.A(_17627_),
    .X(_17628_));
 sky130_fd_sc_hd__buf_1 _48208_ (.A(_17563_),
    .X(_17629_));
 sky130_fd_sc_hd__buf_1 _48209_ (.A(_17629_),
    .X(_17630_));
 sky130_fd_sc_hd__buf_1 _48210_ (.A(_17576_),
    .X(_17631_));
 sky130_fd_sc_hd__buf_1 _48211_ (.A(_17568_),
    .X(_17632_));
 sky130_fd_sc_hd__buf_1 _48212_ (.A(_17632_),
    .X(_17633_));
 sky130_fd_sc_hd__nand2_4 _48213_ (.A(_17633_),
    .B(_21493_),
    .Y(_17634_));
 sky130_fd_sc_hd__o21ai_4 _48214_ (.A1(_17631_),
    .A2(_21506_),
    .B1(_17634_),
    .Y(_17635_));
 sky130_fd_sc_hd__o21a_4 _48215_ (.A1(_17607_),
    .A2(_17609_),
    .B1(_03438_),
    .X(_17636_));
 sky130_fd_sc_hd__a21o_4 _48216_ (.A1(_17630_),
    .A2(_17635_),
    .B1(_17636_),
    .X(_17637_));
 sky130_fd_sc_hd__buf_1 _48217_ (.A(_24245_),
    .X(_17638_));
 sky130_fd_sc_hd__and2_4 _48218_ (.A(_17637_),
    .B(_17638_),
    .X(_17639_));
 sky130_fd_sc_hd__a21oi_4 _48219_ (.A1(_17628_),
    .A2(_17589_),
    .B1(_17639_),
    .Y(_17640_));
 sky130_fd_sc_hd__buf_1 _48220_ (.A(_17556_),
    .X(_17641_));
 sky130_fd_sc_hd__nand4_4 _48221_ (.A(_21351_),
    .B(_05595_),
    .C(_17641_),
    .D(_01492_),
    .Y(_17642_));
 sky130_fd_sc_hd__o21ai_4 _48222_ (.A1(_17625_),
    .A2(_17640_),
    .B1(_17642_),
    .Y(_17643_));
 sky130_fd_sc_hd__buf_1 _48223_ (.A(_21167_),
    .X(_17644_));
 sky130_fd_sc_hd__buf_1 _48224_ (.A(_17644_),
    .X(_17645_));
 sky130_fd_sc_hd__and2_4 _48225_ (.A(_17643_),
    .B(_17645_),
    .X(_24315_));
 sky130_fd_sc_hd__buf_1 _48226_ (.A(_21142_),
    .X(_17646_));
 sky130_fd_sc_hd__nand2_4 _48227_ (.A(_03425_),
    .B(_18660_),
    .Y(_17647_));
 sky130_fd_sc_hd__o21a_4 _48228_ (.A1(_17559_),
    .A2(_21529_),
    .B1(_17647_),
    .X(_17648_));
 sky130_fd_sc_hd__buf_1 _48229_ (.A(_17604_),
    .X(_17649_));
 sky130_fd_sc_hd__buf_1 _48230_ (.A(_17649_),
    .X(_17650_));
 sky130_fd_sc_hd__o21ai_4 _48231_ (.A1(_17616_),
    .A2(_17618_),
    .B1(_17650_),
    .Y(_17651_));
 sky130_fd_sc_hd__o21ai_4 _48232_ (.A1(_03440_),
    .A2(_17648_),
    .B1(_17651_),
    .Y(_17652_));
 sky130_fd_sc_hd__and2_4 _48233_ (.A(_17599_),
    .B(_03448_),
    .X(_17653_));
 sky130_fd_sc_hd__a21o_4 _48234_ (.A1(_17646_),
    .A2(_17652_),
    .B1(_17653_),
    .X(_17654_));
 sky130_fd_sc_hd__and4_4 _48235_ (.A(_17571_),
    .B(_21126_),
    .C(_03458_),
    .D(_17646_),
    .X(_17655_));
 sky130_fd_sc_hd__a21o_4 _48236_ (.A1(_17654_),
    .A2(_21155_),
    .B1(_17655_),
    .X(_17656_));
 sky130_fd_sc_hd__and2_4 _48237_ (.A(_17656_),
    .B(_17645_),
    .X(_24316_));
 sky130_fd_sc_hd__buf_1 _48238_ (.A(_17605_),
    .X(_17657_));
 sky130_fd_sc_hd__nand2_4 _48239_ (.A(_03425_),
    .B(_18651_),
    .Y(_17658_));
 sky130_vsdinv _48240_ (.A(_17658_),
    .Y(_17659_));
 sky130_fd_sc_hd__nor2_4 _48241_ (.A(_17582_),
    .B(_21546_),
    .Y(_17660_));
 sky130_fd_sc_hd__buf_1 _48242_ (.A(_21123_),
    .X(_17661_));
 sky130_fd_sc_hd__buf_1 _48243_ (.A(_17661_),
    .X(_17662_));
 sky130_fd_sc_hd__o21a_4 _48244_ (.A1(_17659_),
    .A2(_17660_),
    .B1(_17662_),
    .X(_17663_));
 sky130_fd_sc_hd__a21o_4 _48245_ (.A1(_17657_),
    .A2(_17635_),
    .B1(_17663_),
    .X(_17664_));
 sky130_fd_sc_hd__and2_4 _48246_ (.A(_17611_),
    .B(_17621_),
    .X(_17665_));
 sky130_fd_sc_hd__a21o_4 _48247_ (.A1(_17614_),
    .A2(_17664_),
    .B1(_17665_),
    .X(_17666_));
 sky130_fd_sc_hd__buf_1 _48248_ (.A(_17552_),
    .X(_17667_));
 sky130_fd_sc_hd__buf_1 _48249_ (.A(_17592_),
    .X(_17668_));
 sky130_fd_sc_hd__buf_1 _48250_ (.A(_17668_),
    .X(_17669_));
 sky130_fd_sc_hd__nor3_4 _48251_ (.A(_01494_),
    .B(_17669_),
    .C(_17565_),
    .Y(_17670_));
 sky130_fd_sc_hd__a21o_4 _48252_ (.A1(_17666_),
    .A2(_17667_),
    .B1(_17670_),
    .X(_17671_));
 sky130_fd_sc_hd__and2_4 _48253_ (.A(_17671_),
    .B(_17645_),
    .X(_24286_));
 sky130_fd_sc_hd__buf_1 _48254_ (.A(_17578_),
    .X(_17672_));
 sky130_fd_sc_hd__nand2_4 _48255_ (.A(_17632_),
    .B(_21545_),
    .Y(_17673_));
 sky130_fd_sc_hd__o21ai_4 _48256_ (.A1(_03426_),
    .A2(_21564_),
    .B1(_17673_),
    .Y(_17674_));
 sky130_fd_sc_hd__nor2_4 _48257_ (.A(_17578_),
    .B(_17648_),
    .Y(_17675_));
 sky130_fd_sc_hd__a21o_4 _48258_ (.A1(_17672_),
    .A2(_17674_),
    .B1(_17675_),
    .X(_17676_));
 sky130_fd_sc_hd__and2_4 _48259_ (.A(_17620_),
    .B(_03448_),
    .X(_17677_));
 sky130_fd_sc_hd__a21o_4 _48260_ (.A1(_17646_),
    .A2(_17676_),
    .B1(_17677_),
    .X(_17678_));
 sky130_fd_sc_hd__buf_1 _48261_ (.A(_18608_),
    .X(_17679_));
 sky130_fd_sc_hd__buf_1 _48262_ (.A(_17679_),
    .X(_17680_));
 sky130_fd_sc_hd__nand3_4 _48263_ (.A(_17581_),
    .B(_17680_),
    .C(_01492_),
    .Y(_17681_));
 sky130_fd_sc_hd__a21bo_4 _48264_ (.A1(_17678_),
    .A2(_21155_),
    .B1_N(_17681_),
    .X(_17682_));
 sky130_fd_sc_hd__and2_4 _48265_ (.A(_17682_),
    .B(_17645_),
    .X(_24287_));
 sky130_fd_sc_hd__buf_1 _48266_ (.A(_01491_),
    .X(_17683_));
 sky130_fd_sc_hd__buf_1 _48267_ (.A(_18629_),
    .X(_17684_));
 sky130_fd_sc_hd__nand2_4 _48268_ (.A(_17684_),
    .B(_18657_),
    .Y(_17685_));
 sky130_fd_sc_hd__o21ai_4 _48269_ (.A1(_17633_),
    .A2(_21580_),
    .B1(_17685_),
    .Y(_17686_));
 sky130_fd_sc_hd__o21a_4 _48270_ (.A1(_17659_),
    .A2(_17660_),
    .B1(_17604_),
    .X(_17687_));
 sky130_fd_sc_hd__a21o_4 _48271_ (.A1(_17600_),
    .A2(_17686_),
    .B1(_17687_),
    .X(_17688_));
 sky130_fd_sc_hd__buf_1 _48272_ (.A(_03447_),
    .X(_17689_));
 sky130_fd_sc_hd__and2_4 _48273_ (.A(_17637_),
    .B(_17689_),
    .X(_17690_));
 sky130_fd_sc_hd__a21o_4 _48274_ (.A1(_17683_),
    .A2(_17688_),
    .B1(_17690_),
    .X(_17691_));
 sky130_fd_sc_hd__buf_1 _48275_ (.A(_17556_),
    .X(_17692_));
 sky130_fd_sc_hd__and2_4 _48276_ (.A(_17594_),
    .B(_17692_),
    .X(_17693_));
 sky130_fd_sc_hd__a21o_4 _48277_ (.A1(_17691_),
    .A2(_21155_),
    .B1(_17693_),
    .X(_17694_));
 sky130_fd_sc_hd__buf_1 _48278_ (.A(_17644_),
    .X(_17695_));
 sky130_fd_sc_hd__and2_4 _48279_ (.A(_17694_),
    .B(_17695_),
    .X(_24288_));
 sky130_fd_sc_hd__buf_1 _48280_ (.A(_18623_),
    .X(_17696_));
 sky130_fd_sc_hd__buf_1 _48281_ (.A(_17696_),
    .X(_17697_));
 sky130_fd_sc_hd__nand2_4 _48282_ (.A(_17572_),
    .B(_18646_),
    .Y(_17698_));
 sky130_vsdinv _48283_ (.A(_17698_),
    .Y(_17699_));
 sky130_fd_sc_hd__buf_1 _48284_ (.A(_03425_),
    .X(_17700_));
 sky130_fd_sc_hd__nor2_4 _48285_ (.A(_17700_),
    .B(_21602_),
    .Y(_17701_));
 sky130_fd_sc_hd__o21a_4 _48286_ (.A1(_17699_),
    .A2(_17701_),
    .B1(_21124_),
    .X(_17702_));
 sky130_fd_sc_hd__a21o_4 _48287_ (.A1(_17697_),
    .A2(_17674_),
    .B1(_17702_),
    .X(_17703_));
 sky130_fd_sc_hd__buf_1 _48288_ (.A(_24245_),
    .X(_17704_));
 sky130_fd_sc_hd__and2_4 _48289_ (.A(_17703_),
    .B(_17704_),
    .X(_17705_));
 sky130_fd_sc_hd__a21o_4 _48290_ (.A1(_17628_),
    .A2(_17652_),
    .B1(_17705_),
    .X(_17706_));
 sky130_fd_sc_hd__and2_4 _48291_ (.A(_17603_),
    .B(_17692_),
    .X(_17707_));
 sky130_fd_sc_hd__a21o_4 _48292_ (.A1(_17706_),
    .A2(_17667_),
    .B1(_17707_),
    .X(_17708_));
 sky130_fd_sc_hd__and2_4 _48293_ (.A(_17708_),
    .B(_17695_),
    .X(_24289_));
 sky130_fd_sc_hd__buf_1 _48294_ (.A(_01494_),
    .X(_17709_));
 sky130_fd_sc_hd__buf_1 _48295_ (.A(_17626_),
    .X(_17710_));
 sky130_fd_sc_hd__buf_1 _48296_ (.A(_17710_),
    .X(_17711_));
 sky130_fd_sc_hd__buf_1 _48297_ (.A(_17566_),
    .X(_17712_));
 sky130_fd_sc_hd__nand2_4 _48298_ (.A(_17684_),
    .B(_21601_),
    .Y(_17713_));
 sky130_vsdinv _48299_ (.A(_17713_),
    .Y(_17714_));
 sky130_fd_sc_hd__nor2_4 _48300_ (.A(_18631_),
    .B(_21622_),
    .Y(_17715_));
 sky130_fd_sc_hd__o21a_4 _48301_ (.A1(_17714_),
    .A2(_17715_),
    .B1(_17672_),
    .X(_17716_));
 sky130_fd_sc_hd__a21o_4 _48302_ (.A1(_17712_),
    .A2(_17686_),
    .B1(_17716_),
    .X(_17717_));
 sky130_fd_sc_hd__buf_1 _48303_ (.A(_21141_),
    .X(_17718_));
 sky130_fd_sc_hd__and2_4 _48304_ (.A(_17717_),
    .B(_17718_),
    .X(_17719_));
 sky130_fd_sc_hd__a21o_4 _48305_ (.A1(_17711_),
    .A2(_17664_),
    .B1(_17719_),
    .X(_17720_));
 sky130_fd_sc_hd__and2_4 _48306_ (.A(_17613_),
    .B(_17692_),
    .X(_17721_));
 sky130_fd_sc_hd__a21o_4 _48307_ (.A1(_17709_),
    .A2(_17720_),
    .B1(_17721_),
    .X(_17722_));
 sky130_fd_sc_hd__and2_4 _48308_ (.A(_17722_),
    .B(_17695_),
    .X(_24290_));
 sky130_fd_sc_hd__buf_1 _48309_ (.A(_17641_),
    .X(_17723_));
 sky130_fd_sc_hd__buf_1 _48310_ (.A(_17564_),
    .X(_17724_));
 sky130_fd_sc_hd__nand2_4 _48311_ (.A(_17632_),
    .B(_18638_),
    .Y(_17725_));
 sky130_fd_sc_hd__o21ai_4 _48312_ (.A1(_17570_),
    .A2(_21640_),
    .B1(_17725_),
    .Y(_17726_));
 sky130_fd_sc_hd__o21a_4 _48313_ (.A1(_17699_),
    .A2(_17701_),
    .B1(_17566_),
    .X(_17727_));
 sky130_fd_sc_hd__a21o_4 _48314_ (.A1(_17724_),
    .A2(_17726_),
    .B1(_17727_),
    .X(_17728_));
 sky130_fd_sc_hd__and2_4 _48315_ (.A(_17676_),
    .B(_17626_),
    .X(_17729_));
 sky130_fd_sc_hd__a21o_4 _48316_ (.A1(_24246_),
    .A2(_17728_),
    .B1(_17729_),
    .X(_17730_));
 sky130_fd_sc_hd__buf_1 _48317_ (.A(_21153_),
    .X(_17731_));
 sky130_fd_sc_hd__and2_4 _48318_ (.A(_17730_),
    .B(_17731_),
    .X(_17732_));
 sky130_fd_sc_hd__a21o_4 _48319_ (.A1(_17723_),
    .A2(_17623_),
    .B1(_17732_),
    .X(_17733_));
 sky130_fd_sc_hd__and2_4 _48320_ (.A(_17733_),
    .B(_17695_),
    .X(_24291_));
 sky130_fd_sc_hd__buf_1 _48321_ (.A(_17641_),
    .X(_17734_));
 sky130_fd_sc_hd__buf_1 _48322_ (.A(_21142_),
    .X(_17735_));
 sky130_fd_sc_hd__nand2_4 _48323_ (.A(_17632_),
    .B(_18642_),
    .Y(_17736_));
 sky130_fd_sc_hd__o21ai_4 _48324_ (.A1(_17583_),
    .A2(_21654_),
    .B1(_17736_),
    .Y(_17737_));
 sky130_fd_sc_hd__buf_1 _48325_ (.A(_17604_),
    .X(_17738_));
 sky130_fd_sc_hd__o21a_4 _48326_ (.A1(_17714_),
    .A2(_17715_),
    .B1(_17738_),
    .X(_17739_));
 sky130_fd_sc_hd__a21o_4 _48327_ (.A1(_17601_),
    .A2(_17737_),
    .B1(_17739_),
    .X(_17740_));
 sky130_fd_sc_hd__buf_1 _48328_ (.A(_03447_),
    .X(_17741_));
 sky130_fd_sc_hd__and2_4 _48329_ (.A(_17688_),
    .B(_17741_),
    .X(_17742_));
 sky130_fd_sc_hd__a211o_4 _48330_ (.A1(_17735_),
    .A2(_17740_),
    .B1(_17679_),
    .C1(_17742_),
    .X(_17743_));
 sky130_vsdinv _48331_ (.A(_17743_),
    .Y(_17744_));
 sky130_fd_sc_hd__a211o_4 _48332_ (.A1(_17734_),
    .A2(_17640_),
    .B1(_17548_),
    .C1(_17744_),
    .X(_17745_));
 sky130_fd_sc_hd__o41ai_4 _48333_ (.A1(_21344_),
    .A2(_17558_),
    .A3(_17595_),
    .A4(_05605_),
    .B1(_17745_),
    .Y(_24292_));
 sky130_fd_sc_hd__buf_1 _48334_ (.A(_18602_),
    .X(_17746_));
 sky130_fd_sc_hd__buf_1 _48335_ (.A(_17746_),
    .X(_17747_));
 sky130_fd_sc_hd__nand2_4 _48336_ (.A(_17654_),
    .B(_17625_),
    .Y(_17748_));
 sky130_fd_sc_hd__buf_1 _48337_ (.A(_17741_),
    .X(_17749_));
 sky130_fd_sc_hd__nand2_4 _48338_ (.A(_18630_),
    .B(_18710_),
    .Y(_17750_));
 sky130_vsdinv _48339_ (.A(_17750_),
    .Y(_17751_));
 sky130_fd_sc_hd__nor2_4 _48340_ (.A(_17617_),
    .B(_21671_),
    .Y(_17752_));
 sky130_fd_sc_hd__buf_1 _48341_ (.A(_17563_),
    .X(_17753_));
 sky130_fd_sc_hd__o21a_4 _48342_ (.A1(_17751_),
    .A2(_17752_),
    .B1(_17753_),
    .X(_17754_));
 sky130_fd_sc_hd__a21o_4 _48343_ (.A1(_17649_),
    .A2(_17726_),
    .B1(_17754_),
    .X(_17755_));
 sky130_fd_sc_hd__and2_4 _48344_ (.A(_17755_),
    .B(_21142_),
    .X(_17756_));
 sky130_fd_sc_hd__a21o_4 _48345_ (.A1(_17749_),
    .A2(_17703_),
    .B1(_17756_),
    .X(_17757_));
 sky130_fd_sc_hd__buf_1 _48346_ (.A(_17552_),
    .X(_17758_));
 sky130_fd_sc_hd__nand2_4 _48347_ (.A(_17757_),
    .B(_17758_),
    .Y(_17759_));
 sky130_fd_sc_hd__buf_1 _48348_ (.A(_03467_),
    .X(_17760_));
 sky130_fd_sc_hd__a21oi_4 _48349_ (.A1(_17748_),
    .A2(_17759_),
    .B1(_17760_),
    .Y(_17761_));
 sky130_fd_sc_hd__a41o_4 _48350_ (.A1(_21156_),
    .A2(_21145_),
    .A3(_17747_),
    .A4(_17551_),
    .B1(_17761_),
    .X(_24293_));
 sky130_fd_sc_hd__nand2_4 _48351_ (.A(_17666_),
    .B(_03459_),
    .Y(_17762_));
 sky130_fd_sc_hd__nand2_4 _48352_ (.A(_17560_),
    .B(_18714_),
    .Y(_17763_));
 sky130_vsdinv _48353_ (.A(_17763_),
    .Y(_17764_));
 sky130_fd_sc_hd__nor2_4 _48354_ (.A(_17576_),
    .B(_21687_),
    .Y(_17765_));
 sky130_fd_sc_hd__o21a_4 _48355_ (.A1(_17764_),
    .A2(_17765_),
    .B1(_17661_),
    .X(_17766_));
 sky130_fd_sc_hd__a21o_4 _48356_ (.A1(_17567_),
    .A2(_17737_),
    .B1(_17766_),
    .X(_17767_));
 sky130_fd_sc_hd__buf_1 _48357_ (.A(_21141_),
    .X(_17768_));
 sky130_fd_sc_hd__and2_4 _48358_ (.A(_17767_),
    .B(_17768_),
    .X(_17769_));
 sky130_fd_sc_hd__a21o_4 _48359_ (.A1(_03449_),
    .A2(_17717_),
    .B1(_17769_),
    .X(_17770_));
 sky130_fd_sc_hd__nand2_4 _48360_ (.A(_17770_),
    .B(_17758_),
    .Y(_17771_));
 sky130_fd_sc_hd__buf_1 _48361_ (.A(_03467_),
    .X(_17772_));
 sky130_fd_sc_hd__a21o_4 _48362_ (.A1(_17762_),
    .A2(_17771_),
    .B1(_17772_),
    .X(_17773_));
 sky130_fd_sc_hd__o41ai_4 _48363_ (.A1(_17558_),
    .A2(_03450_),
    .A3(_17595_),
    .A4(_17565_),
    .B1(_17773_),
    .Y(_24294_));
 sky130_fd_sc_hd__nand2_4 _48364_ (.A(_17678_),
    .B(_17625_),
    .Y(_17774_));
 sky130_fd_sc_hd__nand2_4 _48365_ (.A(_17568_),
    .B(_18705_),
    .Y(_17775_));
 sky130_fd_sc_hd__o21ai_4 _48366_ (.A1(_03427_),
    .A2(_21707_),
    .B1(_17775_),
    .Y(_17776_));
 sky130_fd_sc_hd__o21a_4 _48367_ (.A1(_17751_),
    .A2(_17752_),
    .B1(_17649_),
    .X(_17777_));
 sky130_fd_sc_hd__a21o_4 _48368_ (.A1(_17601_),
    .A2(_17776_),
    .B1(_17777_),
    .X(_17778_));
 sky130_fd_sc_hd__and2_4 _48369_ (.A(_17728_),
    .B(_03448_),
    .X(_17779_));
 sky130_fd_sc_hd__a21o_4 _48370_ (.A1(_21143_),
    .A2(_17778_),
    .B1(_17779_),
    .X(_17780_));
 sky130_fd_sc_hd__nand2_4 _48371_ (.A(_17780_),
    .B(_17758_),
    .Y(_17781_));
 sky130_fd_sc_hd__a21oi_4 _48372_ (.A1(_17774_),
    .A2(_17781_),
    .B1(_17772_),
    .Y(_17782_));
 sky130_fd_sc_hd__a41o_4 _48373_ (.A1(_21156_),
    .A2(_21144_),
    .A3(_17747_),
    .A4(_17581_),
    .B1(_17782_),
    .X(_24295_));
 sky130_fd_sc_hd__buf_1 _48374_ (.A(_17772_),
    .X(_17783_));
 sky130_fd_sc_hd__buf_1 _48375_ (.A(_17617_),
    .X(_17784_));
 sky130_fd_sc_hd__nand2_4 _48376_ (.A(_17569_),
    .B(_18694_),
    .Y(_17785_));
 sky130_fd_sc_hd__o21ai_4 _48377_ (.A1(_17784_),
    .A2(_21722_),
    .B1(_17785_),
    .Y(_17786_));
 sky130_fd_sc_hd__o21a_4 _48378_ (.A1(_17764_),
    .A2(_17765_),
    .B1(_17738_),
    .X(_17787_));
 sky130_fd_sc_hd__a21oi_4 _48379_ (.A1(_21125_),
    .A2(_17786_),
    .B1(_17787_),
    .Y(_17788_));
 sky130_fd_sc_hd__nand2_4 _48380_ (.A(_17740_),
    .B(_17749_),
    .Y(_17789_));
 sky130_fd_sc_hd__o21ai_4 _48381_ (.A1(_17628_),
    .A2(_17788_),
    .B1(_17789_),
    .Y(_17790_));
 sky130_fd_sc_hd__nand2_4 _48382_ (.A(_17790_),
    .B(_17553_),
    .Y(_17791_));
 sky130_fd_sc_hd__a21boi_4 _48383_ (.A1(_17691_),
    .A2(_17558_),
    .B1_N(_17791_),
    .Y(_17792_));
 sky130_fd_sc_hd__buf_1 _48384_ (.A(_17553_),
    .X(_17793_));
 sky130_fd_sc_hd__buf_1 _48385_ (.A(_18602_),
    .X(_17794_));
 sky130_fd_sc_hd__buf_1 _48386_ (.A(_17794_),
    .X(_17795_));
 sky130_fd_sc_hd__nand3_4 _48387_ (.A(_17594_),
    .B(_17793_),
    .C(_17795_),
    .Y(_17796_));
 sky130_fd_sc_hd__o21ai_4 _48388_ (.A1(_17783_),
    .A2(_17792_),
    .B1(_17796_),
    .Y(_24297_));
 sky130_fd_sc_hd__nand2_4 _48389_ (.A(_17706_),
    .B(_17723_),
    .Y(_17797_));
 sky130_fd_sc_hd__buf_1 _48390_ (.A(_17627_),
    .X(_17798_));
 sky130_fd_sc_hd__buf_1 _48391_ (.A(_17696_),
    .X(_17799_));
 sky130_fd_sc_hd__nand2_4 _48392_ (.A(_17684_),
    .B(_18666_),
    .Y(_17800_));
 sky130_vsdinv _48393_ (.A(_17800_),
    .Y(_17801_));
 sky130_fd_sc_hd__nor2_4 _48394_ (.A(_18631_),
    .B(_21740_),
    .Y(_17802_));
 sky130_fd_sc_hd__o21a_4 _48395_ (.A1(_17801_),
    .A2(_17802_),
    .B1(_17672_),
    .X(_17803_));
 sky130_fd_sc_hd__a21o_4 _48396_ (.A1(_17799_),
    .A2(_17776_),
    .B1(_17803_),
    .X(_17804_));
 sky130_fd_sc_hd__and2_4 _48397_ (.A(_17804_),
    .B(_17638_),
    .X(_17805_));
 sky130_fd_sc_hd__a21o_4 _48398_ (.A1(_17798_),
    .A2(_17755_),
    .B1(_17805_),
    .X(_17806_));
 sky130_fd_sc_hd__buf_1 _48399_ (.A(_17731_),
    .X(_17807_));
 sky130_fd_sc_hd__nand2_4 _48400_ (.A(_17806_),
    .B(_17807_),
    .Y(_17808_));
 sky130_fd_sc_hd__buf_1 _48401_ (.A(_17794_),
    .X(_17809_));
 sky130_fd_sc_hd__a21o_4 _48402_ (.A1(_17797_),
    .A2(_17808_),
    .B1(_17809_),
    .X(_17810_));
 sky130_fd_sc_hd__nand3_4 _48403_ (.A(_17603_),
    .B(_17793_),
    .C(_17747_),
    .Y(_17811_));
 sky130_fd_sc_hd__nand2_4 _48404_ (.A(_17810_),
    .B(_17811_),
    .Y(_24298_));
 sky130_fd_sc_hd__nand2_4 _48405_ (.A(_17720_),
    .B(_17723_),
    .Y(_17812_));
 sky130_fd_sc_hd__buf_1 _48406_ (.A(_17710_),
    .X(_17813_));
 sky130_fd_sc_hd__nand2_4 _48407_ (.A(_17684_),
    .B(_21739_),
    .Y(_17814_));
 sky130_vsdinv _48408_ (.A(_17814_),
    .Y(_17815_));
 sky130_fd_sc_hd__nor2_4 _48409_ (.A(_18631_),
    .B(_21751_),
    .Y(_17816_));
 sky130_fd_sc_hd__o21a_4 _48410_ (.A1(_17815_),
    .A2(_17816_),
    .B1(_17672_),
    .X(_17817_));
 sky130_fd_sc_hd__a21o_4 _48411_ (.A1(_17799_),
    .A2(_17786_),
    .B1(_17817_),
    .X(_17818_));
 sky130_fd_sc_hd__and2_4 _48412_ (.A(_17818_),
    .B(_17638_),
    .X(_17819_));
 sky130_fd_sc_hd__a21o_4 _48413_ (.A1(_17813_),
    .A2(_17767_),
    .B1(_17819_),
    .X(_17820_));
 sky130_fd_sc_hd__nand2_4 _48414_ (.A(_17820_),
    .B(_17807_),
    .Y(_17821_));
 sky130_fd_sc_hd__a21o_4 _48415_ (.A1(_17812_),
    .A2(_17821_),
    .B1(_17809_),
    .X(_17822_));
 sky130_fd_sc_hd__nand3_4 _48416_ (.A(_17613_),
    .B(_17793_),
    .C(_17795_),
    .Y(_17823_));
 sky130_fd_sc_hd__nand2_4 _48417_ (.A(_17822_),
    .B(_17823_),
    .Y(_24299_));
 sky130_fd_sc_hd__nand2_4 _48418_ (.A(_17569_),
    .B(_18676_),
    .Y(_17824_));
 sky130_fd_sc_hd__o21ai_4 _48419_ (.A1(_03427_),
    .A2(_21766_),
    .B1(_17824_),
    .Y(_17825_));
 sky130_fd_sc_hd__o21a_4 _48420_ (.A1(_17801_),
    .A2(_17802_),
    .B1(_03438_),
    .X(_17826_));
 sky130_fd_sc_hd__a21o_4 _48421_ (.A1(_17662_),
    .A2(_17825_),
    .B1(_17826_),
    .X(_17827_));
 sky130_fd_sc_hd__and2_4 _48422_ (.A(_17827_),
    .B(_17704_),
    .X(_17828_));
 sky130_fd_sc_hd__a21o_4 _48423_ (.A1(_17628_),
    .A2(_17778_),
    .B1(_17828_),
    .X(_17829_));
 sky130_fd_sc_hd__nand2_4 _48424_ (.A(_17829_),
    .B(_17709_),
    .Y(_17830_));
 sky130_fd_sc_hd__buf_1 _48425_ (.A(_17692_),
    .X(_17831_));
 sky130_fd_sc_hd__nand2_4 _48426_ (.A(_17730_),
    .B(_17831_),
    .Y(_17832_));
 sky130_fd_sc_hd__a21o_4 _48427_ (.A1(_17830_),
    .A2(_17832_),
    .B1(_17809_),
    .X(_17833_));
 sky130_fd_sc_hd__nand3_4 _48428_ (.A(_17623_),
    .B(_17793_),
    .C(_17795_),
    .Y(_17834_));
 sky130_fd_sc_hd__nand2_4 _48429_ (.A(_17833_),
    .B(_17834_),
    .Y(_24300_));
 sky130_fd_sc_hd__a211o_4 _48430_ (.A1(_17735_),
    .A2(_17740_),
    .B1(_24249_),
    .C1(_17742_),
    .X(_17835_));
 sky130_fd_sc_hd__nand2_4 _48431_ (.A(_17582_),
    .B(_18688_),
    .Y(_17836_));
 sky130_vsdinv _48432_ (.A(_17836_),
    .Y(_17837_));
 sky130_fd_sc_hd__nor2_4 _48433_ (.A(_17633_),
    .B(_18728_),
    .Y(_17838_));
 sky130_fd_sc_hd__o21a_4 _48434_ (.A1(_17837_),
    .A2(_17838_),
    .B1(_21124_),
    .X(_17839_));
 sky130_fd_sc_hd__o21a_4 _48435_ (.A1(_17815_),
    .A2(_17816_),
    .B1(_17738_),
    .X(_17840_));
 sky130_fd_sc_hd__or3_4 _48436_ (.A(_17592_),
    .B(_17839_),
    .C(_17840_),
    .X(_17841_));
 sky130_fd_sc_hd__nand2_4 _48437_ (.A(_17788_),
    .B(_17668_),
    .Y(_17842_));
 sky130_fd_sc_hd__a21o_4 _48438_ (.A1(_17841_),
    .A2(_17842_),
    .B1(_03458_),
    .X(_17843_));
 sky130_fd_sc_hd__a21o_4 _48439_ (.A1(_17835_),
    .A2(_17843_),
    .B1(_17746_),
    .X(_17844_));
 sky130_fd_sc_hd__o21ai_4 _48440_ (.A1(_01521_),
    .A2(_17643_),
    .B1(_17844_),
    .Y(_17845_));
 sky130_vsdinv _48441_ (.A(_17845_),
    .Y(_24301_));
 sky130_fd_sc_hd__buf_1 _48442_ (.A(_17556_),
    .X(_17846_));
 sky130_fd_sc_hd__buf_1 _48443_ (.A(_17846_),
    .X(_17847_));
 sky130_fd_sc_hd__nand2_4 _48444_ (.A(_17757_),
    .B(_17847_),
    .Y(_17848_));
 sky130_fd_sc_hd__nand2_4 _48445_ (.A(_17804_),
    .B(_17813_),
    .Y(_17849_));
 sky130_fd_sc_hd__buf_1 _48446_ (.A(_03438_),
    .X(_17850_));
 sky130_fd_sc_hd__buf_1 _48447_ (.A(_17850_),
    .X(_17851_));
 sky130_fd_sc_hd__nand2_4 _48448_ (.A(_17582_),
    .B(_18731_),
    .Y(_17852_));
 sky130_vsdinv _48449_ (.A(_17852_),
    .Y(_17853_));
 sky130_fd_sc_hd__buf_1 _48450_ (.A(_17584_),
    .X(_17854_));
 sky130_fd_sc_hd__nor2_4 _48451_ (.A(_17854_),
    .B(_21793_),
    .Y(_17855_));
 sky130_fd_sc_hd__o21a_4 _48452_ (.A1(_17853_),
    .A2(_17855_),
    .B1(_17630_),
    .X(_17856_));
 sky130_fd_sc_hd__a21o_4 _48453_ (.A1(_17851_),
    .A2(_17825_),
    .B1(_17856_),
    .X(_17857_));
 sky130_fd_sc_hd__buf_1 _48454_ (.A(_24246_),
    .X(_17858_));
 sky130_fd_sc_hd__nand2_4 _48455_ (.A(_17857_),
    .B(_17858_),
    .Y(_17859_));
 sky130_fd_sc_hd__a21o_4 _48456_ (.A1(_17849_),
    .A2(_17859_),
    .B1(_17557_),
    .X(_17860_));
 sky130_fd_sc_hd__a21oi_4 _48457_ (.A1(_17848_),
    .A2(_17860_),
    .B1(_17795_),
    .Y(_17861_));
 sky130_fd_sc_hd__a21o_4 _48458_ (.A1(_17549_),
    .A2(_17656_),
    .B1(_17861_),
    .X(_24302_));
 sky130_fd_sc_hd__buf_1 _48459_ (.A(_17548_),
    .X(_17862_));
 sky130_fd_sc_hd__nand2_4 _48460_ (.A(_17770_),
    .B(_17847_),
    .Y(_17863_));
 sky130_fd_sc_hd__nand2_4 _48461_ (.A(_17818_),
    .B(_17813_),
    .Y(_17864_));
 sky130_fd_sc_hd__buf_1 _48462_ (.A(_17630_),
    .X(_17865_));
 sky130_fd_sc_hd__buf_1 _48463_ (.A(_17784_),
    .X(_17866_));
 sky130_fd_sc_hd__nand2_4 _48464_ (.A(_17568_),
    .B(_18764_),
    .Y(_17867_));
 sky130_fd_sc_hd__o21ai_4 _48465_ (.A1(_17866_),
    .A2(_21804_),
    .B1(_17867_),
    .Y(_17868_));
 sky130_fd_sc_hd__o21a_4 _48466_ (.A1(_17837_),
    .A2(_17838_),
    .B1(_03439_),
    .X(_17869_));
 sky130_fd_sc_hd__a21o_4 _48467_ (.A1(_17865_),
    .A2(_17868_),
    .B1(_17869_),
    .X(_17870_));
 sky130_fd_sc_hd__nand2_4 _48468_ (.A(_17870_),
    .B(_17858_),
    .Y(_17871_));
 sky130_fd_sc_hd__a21o_4 _48469_ (.A1(_17864_),
    .A2(_17871_),
    .B1(_17557_),
    .X(_17872_));
 sky130_fd_sc_hd__buf_1 _48470_ (.A(_17746_),
    .X(_17873_));
 sky130_fd_sc_hd__a21oi_4 _48471_ (.A1(_17863_),
    .A2(_17872_),
    .B1(_17873_),
    .Y(_17874_));
 sky130_fd_sc_hd__a21o_4 _48472_ (.A1(_17862_),
    .A2(_17671_),
    .B1(_17874_),
    .X(_24303_));
 sky130_fd_sc_hd__nand2_4 _48473_ (.A(_17780_),
    .B(_17847_),
    .Y(_17875_));
 sky130_fd_sc_hd__nand2_4 _48474_ (.A(_17827_),
    .B(_17813_),
    .Y(_17876_));
 sky130_fd_sc_hd__nand2_4 _48475_ (.A(_17569_),
    .B(_18720_),
    .Y(_17877_));
 sky130_fd_sc_hd__o21ai_4 _48476_ (.A1(_17854_),
    .A2(_21822_),
    .B1(_17877_),
    .Y(_17878_));
 sky130_fd_sc_hd__o21a_4 _48477_ (.A1(_17853_),
    .A2(_17855_),
    .B1(_03439_),
    .X(_17879_));
 sky130_fd_sc_hd__a21o_4 _48478_ (.A1(_17865_),
    .A2(_17878_),
    .B1(_17879_),
    .X(_17880_));
 sky130_fd_sc_hd__buf_1 _48479_ (.A(_17591_),
    .X(_17881_));
 sky130_fd_sc_hd__nand2_4 _48480_ (.A(_17880_),
    .B(_17881_),
    .Y(_17882_));
 sky130_fd_sc_hd__buf_1 _48481_ (.A(_17679_),
    .X(_17883_));
 sky130_fd_sc_hd__a21o_4 _48482_ (.A1(_17876_),
    .A2(_17882_),
    .B1(_17883_),
    .X(_17884_));
 sky130_fd_sc_hd__a21oi_4 _48483_ (.A1(_17875_),
    .A2(_17884_),
    .B1(_17873_),
    .Y(_17885_));
 sky130_fd_sc_hd__a21o_4 _48484_ (.A1(_17862_),
    .A2(_17682_),
    .B1(_17885_),
    .X(_24304_));
 sky130_fd_sc_hd__buf_1 _48485_ (.A(_03468_),
    .X(_17886_));
 sky130_fd_sc_hd__nand2_4 _48486_ (.A(_17790_),
    .B(_17847_),
    .Y(_17887_));
 sky130_fd_sc_hd__nand2_4 _48487_ (.A(_17868_),
    .B(_03440_),
    .Y(_17888_));
 sky130_fd_sc_hd__nand2_4 _48488_ (.A(_17570_),
    .B(_18757_),
    .Y(_17889_));
 sky130_fd_sc_hd__o21ai_4 _48489_ (.A1(_03428_),
    .A2(_21834_),
    .B1(_17889_),
    .Y(_17890_));
 sky130_fd_sc_hd__nand2_4 _48490_ (.A(_17890_),
    .B(_21126_),
    .Y(_17891_));
 sky130_fd_sc_hd__a21oi_4 _48491_ (.A1(_17888_),
    .A2(_17891_),
    .B1(_17669_),
    .Y(_17892_));
 sky130_fd_sc_hd__o21a_4 _48492_ (.A1(_17839_),
    .A2(_17840_),
    .B1(_03449_),
    .X(_17893_));
 sky130_fd_sc_hd__buf_1 _48493_ (.A(_17731_),
    .X(_17894_));
 sky130_fd_sc_hd__o21ai_4 _48494_ (.A1(_17892_),
    .A2(_17893_),
    .B1(_17894_),
    .Y(_17895_));
 sky130_fd_sc_hd__a21oi_4 _48495_ (.A1(_17887_),
    .A2(_17895_),
    .B1(_17873_),
    .Y(_17896_));
 sky130_fd_sc_hd__a21o_4 _48496_ (.A1(_17694_),
    .A2(_17886_),
    .B1(_17896_),
    .X(_24305_));
 sky130_fd_sc_hd__buf_1 _48497_ (.A(_17846_),
    .X(_17897_));
 sky130_fd_sc_hd__nand2_4 _48498_ (.A(_17806_),
    .B(_17897_),
    .Y(_17898_));
 sky130_fd_sc_hd__buf_1 _48499_ (.A(_17710_),
    .X(_17899_));
 sky130_fd_sc_hd__nand2_4 _48500_ (.A(_17857_),
    .B(_17899_),
    .Y(_17900_));
 sky130_fd_sc_hd__buf_1 _48501_ (.A(_17850_),
    .X(_17901_));
 sky130_fd_sc_hd__nand2_4 _48502_ (.A(_17878_),
    .B(_17901_),
    .Y(_17902_));
 sky130_fd_sc_hd__nand2_4 _48503_ (.A(_17584_),
    .B(_18746_),
    .Y(_17903_));
 sky130_fd_sc_hd__o21ai_4 _48504_ (.A1(_17854_),
    .A2(_21854_),
    .B1(_17903_),
    .Y(_17904_));
 sky130_fd_sc_hd__buf_1 _48505_ (.A(_17662_),
    .X(_17905_));
 sky130_fd_sc_hd__nand2_4 _48506_ (.A(_17904_),
    .B(_17905_),
    .Y(_17906_));
 sky130_fd_sc_hd__buf_1 _48507_ (.A(_17741_),
    .X(_17907_));
 sky130_fd_sc_hd__a21o_4 _48508_ (.A1(_17902_),
    .A2(_17906_),
    .B1(_17907_),
    .X(_17908_));
 sky130_fd_sc_hd__a21o_4 _48509_ (.A1(_17900_),
    .A2(_17908_),
    .B1(_17883_),
    .X(_17909_));
 sky130_fd_sc_hd__a21oi_4 _48510_ (.A1(_17898_),
    .A2(_17909_),
    .B1(_17873_),
    .Y(_17910_));
 sky130_fd_sc_hd__a21o_4 _48511_ (.A1(_17862_),
    .A2(_17708_),
    .B1(_17910_),
    .X(_24306_));
 sky130_fd_sc_hd__buf_1 _48512_ (.A(_03468_),
    .X(_17911_));
 sky130_fd_sc_hd__nand2_4 _48513_ (.A(_17820_),
    .B(_17897_),
    .Y(_17912_));
 sky130_fd_sc_hd__nand2_4 _48514_ (.A(_17870_),
    .B(_17899_),
    .Y(_17913_));
 sky130_fd_sc_hd__nand2_4 _48515_ (.A(_21109_),
    .B(_21869_),
    .Y(_17914_));
 sky130_fd_sc_hd__nand2_4 _48516_ (.A(_17633_),
    .B(_18751_),
    .Y(_17915_));
 sky130_fd_sc_hd__buf_1 _48517_ (.A(_17738_),
    .X(_17916_));
 sky130_fd_sc_hd__a21o_4 _48518_ (.A1(_17914_),
    .A2(_17915_),
    .B1(_17916_),
    .X(_17917_));
 sky130_fd_sc_hd__nand2_4 _48519_ (.A(_17890_),
    .B(_17657_),
    .Y(_17918_));
 sky130_fd_sc_hd__a21o_4 _48520_ (.A1(_17917_),
    .A2(_17918_),
    .B1(_17907_),
    .X(_17919_));
 sky130_fd_sc_hd__a21o_4 _48521_ (.A1(_17913_),
    .A2(_17919_),
    .B1(_17883_),
    .X(_17920_));
 sky130_fd_sc_hd__buf_1 _48522_ (.A(_17746_),
    .X(_17921_));
 sky130_fd_sc_hd__a21oi_4 _48523_ (.A1(_17912_),
    .A2(_17920_),
    .B1(_17921_),
    .Y(_17922_));
 sky130_fd_sc_hd__a21o_4 _48524_ (.A1(_17722_),
    .A2(_17911_),
    .B1(_17922_),
    .X(_24308_));
 sky130_fd_sc_hd__nand2_4 _48525_ (.A(_17829_),
    .B(_17897_),
    .Y(_17923_));
 sky130_fd_sc_hd__nand2_4 _48526_ (.A(_17880_),
    .B(_17899_),
    .Y(_17924_));
 sky130_fd_sc_hd__and2_4 _48527_ (.A(_17904_),
    .B(_17916_),
    .X(_17925_));
 sky130_fd_sc_hd__nor2_4 _48528_ (.A(_17631_),
    .B(_05413_),
    .Y(_17926_));
 sky130_vsdinv _48529_ (.A(_17926_),
    .Y(_17927_));
 sky130_fd_sc_hd__nand2_4 _48530_ (.A(_17559_),
    .B(pcpi_rs1[30]),
    .Y(_17928_));
 sky130_fd_sc_hd__a21oi_4 _48531_ (.A1(_17927_),
    .A2(_17928_),
    .B1(_03440_),
    .Y(_17929_));
 sky130_fd_sc_hd__o21ai_4 _48532_ (.A1(_17925_),
    .A2(_17929_),
    .B1(_17614_),
    .Y(_17930_));
 sky130_fd_sc_hd__a21o_4 _48533_ (.A1(_17924_),
    .A2(_17930_),
    .B1(_17883_),
    .X(_17931_));
 sky130_fd_sc_hd__a21oi_4 _48534_ (.A1(_17923_),
    .A2(_17931_),
    .B1(_17921_),
    .Y(_17932_));
 sky130_fd_sc_hd__a21o_4 _48535_ (.A1(_17733_),
    .A2(_17911_),
    .B1(_17932_),
    .X(_24309_));
 sky130_fd_sc_hd__o21ai_4 _48536_ (.A1(_21109_),
    .A2(_05413_),
    .B1(_17914_),
    .Y(_17933_));
 sky130_fd_sc_hd__o21ai_4 _48537_ (.A1(_17784_),
    .A2(_21834_),
    .B1(_17915_),
    .Y(_17934_));
 sky130_fd_sc_hd__and2_4 _48538_ (.A(_17934_),
    .B(_17724_),
    .X(_17935_));
 sky130_fd_sc_hd__a21o_4 _48539_ (.A1(_17933_),
    .A2(_17650_),
    .B1(_17935_),
    .X(_17936_));
 sky130_fd_sc_hd__o21ai_4 _48540_ (.A1(_17631_),
    .A2(_21804_),
    .B1(_17889_),
    .Y(_17937_));
 sky130_fd_sc_hd__o21ai_4 _48541_ (.A1(_17572_),
    .A2(_18728_),
    .B1(_17867_),
    .Y(_17938_));
 sky130_fd_sc_hd__and2_4 _48542_ (.A(_17938_),
    .B(_17661_),
    .X(_17939_));
 sky130_fd_sc_hd__a21o_4 _48543_ (.A1(_17799_),
    .A2(_17937_),
    .B1(_17939_),
    .X(_17940_));
 sky130_fd_sc_hd__and2_4 _48544_ (.A(_17940_),
    .B(_17638_),
    .X(_17941_));
 sky130_fd_sc_hd__a21o_4 _48545_ (.A1(_17798_),
    .A2(_17936_),
    .B1(_17941_),
    .X(_17942_));
 sky130_fd_sc_hd__buf_1 _48546_ (.A(_17575_),
    .X(_17943_));
 sky130_fd_sc_hd__o21ai_4 _48547_ (.A1(_17943_),
    .A2(_18673_),
    .B1(_17836_),
    .Y(_17944_));
 sky130_fd_sc_hd__o21ai_4 _48548_ (.A1(_17943_),
    .A2(_21722_),
    .B1(_17814_),
    .Y(_17945_));
 sky130_fd_sc_hd__buf_1 _48549_ (.A(_17563_),
    .X(_17946_));
 sky130_fd_sc_hd__and2_4 _48550_ (.A(_17945_),
    .B(_17946_),
    .X(_17947_));
 sky130_fd_sc_hd__a21o_4 _48551_ (.A1(_17697_),
    .A2(_17944_),
    .B1(_17947_),
    .X(_17948_));
 sky130_fd_sc_hd__o21ai_4 _48552_ (.A1(_17608_),
    .A2(_21687_),
    .B1(_17785_),
    .Y(_17949_));
 sky130_fd_sc_hd__o21ai_4 _48553_ (.A1(_18630_),
    .A2(_21654_),
    .B1(_17763_),
    .Y(_17950_));
 sky130_fd_sc_hd__and2_4 _48554_ (.A(_17950_),
    .B(_21123_),
    .X(_17951_));
 sky130_fd_sc_hd__a21o_4 _48555_ (.A1(_17696_),
    .A2(_17949_),
    .B1(_17951_),
    .X(_17952_));
 sky130_fd_sc_hd__and2_4 _48556_ (.A(_17952_),
    .B(_17590_),
    .X(_17953_));
 sky130_fd_sc_hd__a21o_4 _48557_ (.A1(_17627_),
    .A2(_17948_),
    .B1(_17953_),
    .X(_17954_));
 sky130_fd_sc_hd__and2_4 _48558_ (.A(_17954_),
    .B(_21154_),
    .X(_17955_));
 sky130_fd_sc_hd__a21o_4 _48559_ (.A1(_17734_),
    .A2(_17942_),
    .B1(_17955_),
    .X(_17956_));
 sky130_fd_sc_hd__buf_1 _48560_ (.A(_17689_),
    .X(_17957_));
 sky130_fd_sc_hd__o21ai_4 _48561_ (.A1(_03426_),
    .A2(_21622_),
    .B1(_17736_),
    .Y(_17958_));
 sky130_fd_sc_hd__o21ai_4 _48562_ (.A1(_03426_),
    .A2(_21580_),
    .B1(_17713_),
    .Y(_17959_));
 sky130_fd_sc_hd__and2_4 _48563_ (.A(_17959_),
    .B(_17629_),
    .X(_17960_));
 sky130_fd_sc_hd__a21o_4 _48564_ (.A1(_17712_),
    .A2(_17958_),
    .B1(_17960_),
    .X(_17961_));
 sky130_fd_sc_hd__o21ai_4 _48565_ (.A1(_17700_),
    .A2(_21546_),
    .B1(_17685_),
    .Y(_17962_));
 sky130_fd_sc_hd__o21ai_4 _48566_ (.A1(_17700_),
    .A2(_21506_),
    .B1(_17658_),
    .Y(_17963_));
 sky130_fd_sc_hd__and2_4 _48567_ (.A(_17963_),
    .B(_17753_),
    .X(_17964_));
 sky130_fd_sc_hd__a21o_4 _48568_ (.A1(_17605_),
    .A2(_17962_),
    .B1(_17964_),
    .X(_17965_));
 sky130_fd_sc_hd__and2_4 _48569_ (.A(_17965_),
    .B(_17768_),
    .X(_17966_));
 sky130_fd_sc_hd__a21o_4 _48570_ (.A1(_17957_),
    .A2(_17961_),
    .B1(_17966_),
    .X(_17967_));
 sky130_fd_sc_hd__nand2_4 _48571_ (.A(_17967_),
    .B(_17897_),
    .Y(_17968_));
 sky130_fd_sc_hd__o21ai_4 _48572_ (.A1(_17631_),
    .A2(_21471_),
    .B1(_17634_),
    .Y(_17969_));
 sky130_fd_sc_hd__o21ai_4 _48573_ (.A1(_03427_),
    .A2(_21435_),
    .B1(_17606_),
    .Y(_17970_));
 sky130_fd_sc_hd__and2_4 _48574_ (.A(_17970_),
    .B(_17662_),
    .X(_17971_));
 sky130_fd_sc_hd__a21o_4 _48575_ (.A1(_17851_),
    .A2(_17969_),
    .B1(_17971_),
    .X(_17972_));
 sky130_fd_sc_hd__nand2_4 _48576_ (.A(_17972_),
    .B(_17899_),
    .Y(_17973_));
 sky130_fd_sc_hd__o21ai_4 _48577_ (.A1(_17866_),
    .A2(_21389_),
    .B1(_17585_),
    .Y(_17974_));
 sky130_fd_sc_hd__nand2_4 _48578_ (.A(_17974_),
    .B(_17901_),
    .Y(_17975_));
 sky130_fd_sc_hd__o21ai_4 _48579_ (.A1(_03428_),
    .A2(_21344_),
    .B1(_17561_),
    .Y(_17976_));
 sky130_fd_sc_hd__nand2_4 _48580_ (.A(_17976_),
    .B(_17905_),
    .Y(_17977_));
 sky130_fd_sc_hd__a21o_4 _48581_ (.A1(_17975_),
    .A2(_17977_),
    .B1(_17907_),
    .X(_17978_));
 sky130_fd_sc_hd__buf_1 _48582_ (.A(_17679_),
    .X(_17979_));
 sky130_fd_sc_hd__a21o_4 _48583_ (.A1(_17973_),
    .A2(_17978_),
    .B1(_17979_),
    .X(_17980_));
 sky130_fd_sc_hd__a21oi_4 _48584_ (.A1(_17968_),
    .A2(_17980_),
    .B1(_17921_),
    .Y(_17981_));
 sky130_fd_sc_hd__a21o_4 _48585_ (.A1(_17956_),
    .A2(_17911_),
    .B1(_17981_),
    .X(_24317_));
 sky130_fd_sc_hd__o21ai_4 _48586_ (.A1(_17583_),
    .A2(_18758_),
    .B1(_17903_),
    .Y(_17982_));
 sky130_fd_sc_hd__o21ai_4 _48587_ (.A1(_17943_),
    .A2(_21793_),
    .B1(_17877_),
    .Y(_17983_));
 sky130_fd_sc_hd__and2_4 _48588_ (.A(_17983_),
    .B(_17946_),
    .X(_17984_));
 sky130_fd_sc_hd__a21o_4 _48589_ (.A1(_17799_),
    .A2(_17982_),
    .B1(_17984_),
    .X(_17985_));
 sky130_fd_sc_hd__nor2_4 _48590_ (.A(instr_sra),
    .B(instr_srai),
    .Y(_17986_));
 sky130_fd_sc_hd__nor3_4 _48591_ (.A(_17661_),
    .B(_05412_),
    .C(_17986_),
    .Y(_17987_));
 sky130_fd_sc_hd__o21ai_4 _48592_ (.A1(_17617_),
    .A2(_21854_),
    .B1(_17928_),
    .Y(_17988_));
 sky130_fd_sc_hd__and2_4 _48593_ (.A(_17988_),
    .B(_17564_),
    .X(_17989_));
 sky130_fd_sc_hd__a211o_4 _48594_ (.A1(_17649_),
    .A2(_17926_),
    .B1(_17987_),
    .C1(_17989_),
    .X(_17990_));
 sky130_fd_sc_hd__and2_4 _48595_ (.A(_17990_),
    .B(_17621_),
    .X(_17991_));
 sky130_fd_sc_hd__a21o_4 _48596_ (.A1(_17858_),
    .A2(_17985_),
    .B1(_17991_),
    .X(_17992_));
 sky130_fd_sc_hd__o21ai_4 _48597_ (.A1(_17608_),
    .A2(_21766_),
    .B1(_17852_),
    .Y(_17993_));
 sky130_fd_sc_hd__o21ai_4 _48598_ (.A1(_17943_),
    .A2(_21740_),
    .B1(_17824_),
    .Y(_17994_));
 sky130_fd_sc_hd__and2_4 _48599_ (.A(_17994_),
    .B(_17946_),
    .X(_17995_));
 sky130_fd_sc_hd__a21o_4 _48600_ (.A1(_17697_),
    .A2(_17993_),
    .B1(_17995_),
    .X(_17996_));
 sky130_fd_sc_hd__o21ai_4 _48601_ (.A1(_17608_),
    .A2(_21707_),
    .B1(_17800_),
    .Y(_17997_));
 sky130_fd_sc_hd__o21ai_4 _48602_ (.A1(_17575_),
    .A2(_21671_),
    .B1(_17775_),
    .Y(_17998_));
 sky130_fd_sc_hd__and2_4 _48603_ (.A(_17998_),
    .B(_21123_),
    .X(_17999_));
 sky130_fd_sc_hd__a21o_4 _48604_ (.A1(_17696_),
    .A2(_17997_),
    .B1(_17999_),
    .X(_18000_));
 sky130_fd_sc_hd__and2_4 _48605_ (.A(_18000_),
    .B(_17590_),
    .X(_18001_));
 sky130_fd_sc_hd__a21o_4 _48606_ (.A1(_17627_),
    .A2(_17996_),
    .B1(_18001_),
    .X(_18002_));
 sky130_fd_sc_hd__and2_4 _48607_ (.A(_18002_),
    .B(_21154_),
    .X(_18003_));
 sky130_fd_sc_hd__a21o_4 _48608_ (.A1(_17734_),
    .A2(_17992_),
    .B1(_18003_),
    .X(_18004_));
 sky130_fd_sc_hd__o21ai_4 _48609_ (.A1(_17700_),
    .A2(_21563_),
    .B1(_17698_),
    .Y(_18005_));
 sky130_fd_sc_hd__o21ai_4 _48610_ (.A1(_17784_),
    .A2(_21529_),
    .B1(_17673_),
    .Y(_18006_));
 sky130_fd_sc_hd__and2_4 _48611_ (.A(_18006_),
    .B(_17724_),
    .X(_18007_));
 sky130_fd_sc_hd__a21o_4 _48612_ (.A1(_17650_),
    .A2(_18005_),
    .B1(_18007_),
    .X(_18008_));
 sky130_fd_sc_hd__o21ai_4 _48613_ (.A1(_17570_),
    .A2(_21640_),
    .B1(_17750_),
    .Y(_18009_));
 sky130_fd_sc_hd__o21ai_4 _48614_ (.A1(_17576_),
    .A2(_21602_),
    .B1(_17725_),
    .Y(_18010_));
 sky130_fd_sc_hd__and2_4 _48615_ (.A(_18010_),
    .B(_17629_),
    .X(_18011_));
 sky130_fd_sc_hd__a21o_4 _48616_ (.A1(_17712_),
    .A2(_18009_),
    .B1(_18011_),
    .X(_18012_));
 sky130_fd_sc_hd__and2_4 _48617_ (.A(_18012_),
    .B(_17621_),
    .X(_18013_));
 sky130_fd_sc_hd__a21o_4 _48618_ (.A1(_17614_),
    .A2(_18008_),
    .B1(_18013_),
    .X(_18014_));
 sky130_fd_sc_hd__buf_1 _48619_ (.A(_17846_),
    .X(_18015_));
 sky130_fd_sc_hd__nand2_4 _48620_ (.A(_18014_),
    .B(_18015_),
    .Y(_18016_));
 sky130_fd_sc_hd__o21ai_4 _48621_ (.A1(_17854_),
    .A2(_21455_),
    .B1(_17615_),
    .Y(_18017_));
 sky130_vsdinv _48622_ (.A(_17647_),
    .Y(_18018_));
 sky130_fd_sc_hd__o21a_4 _48623_ (.A1(_18018_),
    .A2(_17618_),
    .B1(_17850_),
    .X(_18019_));
 sky130_fd_sc_hd__a21o_4 _48624_ (.A1(_17865_),
    .A2(_18017_),
    .B1(_18019_),
    .X(_18020_));
 sky130_fd_sc_hd__buf_1 _48625_ (.A(_17710_),
    .X(_18021_));
 sky130_fd_sc_hd__nand2_4 _48626_ (.A(_18020_),
    .B(_18021_),
    .Y(_18022_));
 sky130_fd_sc_hd__o21ai_4 _48627_ (.A1(_17574_),
    .A2(_17550_),
    .B1(_17865_),
    .Y(_18023_));
 sky130_fd_sc_hd__o21ai_4 _48628_ (.A1(_17866_),
    .A2(_21409_),
    .B1(_17596_),
    .Y(_18024_));
 sky130_fd_sc_hd__nand2_4 _48629_ (.A(_18024_),
    .B(_17657_),
    .Y(_18025_));
 sky130_fd_sc_hd__a21o_4 _48630_ (.A1(_18023_),
    .A2(_18025_),
    .B1(_17907_),
    .X(_18026_));
 sky130_fd_sc_hd__a21o_4 _48631_ (.A1(_18022_),
    .A2(_18026_),
    .B1(_17979_),
    .X(_18027_));
 sky130_fd_sc_hd__a21oi_4 _48632_ (.A1(_18016_),
    .A2(_18027_),
    .B1(_17921_),
    .Y(_18028_));
 sky130_fd_sc_hd__a21o_4 _48633_ (.A1(_18004_),
    .A2(_17911_),
    .B1(_18028_),
    .X(_24328_));
 sky130_fd_sc_hd__and2_4 _48634_ (.A(_17937_),
    .B(_17587_),
    .X(_18029_));
 sky130_fd_sc_hd__a21o_4 _48635_ (.A1(_17657_),
    .A2(_17934_),
    .B1(_18029_),
    .X(_18030_));
 sky130_fd_sc_hd__a21oi_4 _48636_ (.A1(_17933_),
    .A2(_17601_),
    .B1(_17987_),
    .Y(_18031_));
 sky130_fd_sc_hd__nor2_4 _48637_ (.A(_17735_),
    .B(_18031_),
    .Y(_18032_));
 sky130_fd_sc_hd__a21o_4 _48638_ (.A1(_18030_),
    .A2(_17858_),
    .B1(_18032_),
    .X(_18033_));
 sky130_fd_sc_hd__and2_4 _48639_ (.A(_17949_),
    .B(_17946_),
    .X(_18034_));
 sky130_fd_sc_hd__a21o_4 _48640_ (.A1(_17697_),
    .A2(_17945_),
    .B1(_18034_),
    .X(_18035_));
 sky130_fd_sc_hd__and2_4 _48641_ (.A(_17938_),
    .B(_18623_),
    .X(_18036_));
 sky130_fd_sc_hd__a21o_4 _48642_ (.A1(_21124_),
    .A2(_17944_),
    .B1(_18036_),
    .X(_18037_));
 sky130_fd_sc_hd__and2_4 _48643_ (.A(_18037_),
    .B(_17626_),
    .X(_18038_));
 sky130_fd_sc_hd__a21o_4 _48644_ (.A1(_01491_),
    .A2(_18035_),
    .B1(_18038_),
    .X(_18039_));
 sky130_fd_sc_hd__and2_4 _48645_ (.A(_18039_),
    .B(_21154_),
    .X(_18040_));
 sky130_fd_sc_hd__a21o_4 _48646_ (.A1(_17734_),
    .A2(_18033_),
    .B1(_18040_),
    .X(_18041_));
 sky130_fd_sc_hd__and2_4 _48647_ (.A(_17958_),
    .B(_17629_),
    .X(_18042_));
 sky130_fd_sc_hd__a21o_4 _48648_ (.A1(_17712_),
    .A2(_17950_),
    .B1(_18042_),
    .X(_18043_));
 sky130_fd_sc_hd__and2_4 _48649_ (.A(_17962_),
    .B(_17753_),
    .X(_18044_));
 sky130_fd_sc_hd__a21o_4 _48650_ (.A1(_17567_),
    .A2(_17959_),
    .B1(_18044_),
    .X(_18045_));
 sky130_fd_sc_hd__and2_4 _48651_ (.A(_18045_),
    .B(_17768_),
    .X(_18046_));
 sky130_fd_sc_hd__a21o_4 _48652_ (.A1(_03449_),
    .A2(_18043_),
    .B1(_18046_),
    .X(_18047_));
 sky130_fd_sc_hd__nand2_4 _48653_ (.A(_18047_),
    .B(_18015_),
    .Y(_18048_));
 sky130_fd_sc_hd__and2_4 _48654_ (.A(_17969_),
    .B(_17587_),
    .X(_18049_));
 sky130_fd_sc_hd__a21o_4 _48655_ (.A1(_17851_),
    .A2(_17963_),
    .B1(_18049_),
    .X(_18050_));
 sky130_fd_sc_hd__nand2_4 _48656_ (.A(_18050_),
    .B(_18021_),
    .Y(_18051_));
 sky130_fd_sc_hd__nand2_4 _48657_ (.A(_17970_),
    .B(_17901_),
    .Y(_18052_));
 sky130_fd_sc_hd__nand2_4 _48658_ (.A(_17974_),
    .B(_17905_),
    .Y(_18053_));
 sky130_fd_sc_hd__a21o_4 _48659_ (.A1(_18052_),
    .A2(_18053_),
    .B1(_17668_),
    .X(_18054_));
 sky130_fd_sc_hd__a21o_4 _48660_ (.A1(_18051_),
    .A2(_18054_),
    .B1(_17979_),
    .X(_18055_));
 sky130_fd_sc_hd__buf_1 _48661_ (.A(_17794_),
    .X(_18056_));
 sky130_fd_sc_hd__a21oi_4 _48662_ (.A1(_18048_),
    .A2(_18055_),
    .B1(_18056_),
    .Y(_18057_));
 sky130_fd_sc_hd__a21o_4 _48663_ (.A1(_18041_),
    .A2(_17747_),
    .B1(_18057_),
    .X(_24339_));
 sky130_fd_sc_hd__and2_4 _48664_ (.A(_17997_),
    .B(_17600_),
    .X(_18058_));
 sky130_fd_sc_hd__a21o_4 _48665_ (.A1(_17916_),
    .A2(_17994_),
    .B1(_18058_),
    .X(_18059_));
 sky130_fd_sc_hd__and2_4 _48666_ (.A(_17993_),
    .B(_17579_),
    .X(_18060_));
 sky130_fd_sc_hd__a21o_4 _48667_ (.A1(_17850_),
    .A2(_17983_),
    .B1(_18060_),
    .X(_18061_));
 sky130_fd_sc_hd__and2_4 _48668_ (.A(_18061_),
    .B(_17689_),
    .X(_18062_));
 sky130_fd_sc_hd__a21o_4 _48669_ (.A1(_17683_),
    .A2(_18059_),
    .B1(_18062_),
    .X(_18063_));
 sky130_fd_sc_hd__buf_1 _48670_ (.A(_17552_),
    .X(_18064_));
 sky130_fd_sc_hd__and2_4 _48671_ (.A(_17982_),
    .B(_17724_),
    .X(_18065_));
 sky130_fd_sc_hd__a21o_4 _48672_ (.A1(_17650_),
    .A2(_17988_),
    .B1(_18065_),
    .X(_18066_));
 sky130_fd_sc_hd__buf_1 _48673_ (.A(_17986_),
    .X(_18067_));
 sky130_fd_sc_hd__o21ai_4 _48674_ (.A1(_17866_),
    .A2(_03439_),
    .B1(_18067_),
    .Y(_18068_));
 sky130_fd_sc_hd__and3_4 _48675_ (.A(_18068_),
    .B(_17741_),
    .C(_21905_),
    .X(_18069_));
 sky130_fd_sc_hd__a21oi_4 _48676_ (.A1(_18066_),
    .A2(_17646_),
    .B1(_18069_),
    .Y(_18070_));
 sky130_fd_sc_hd__nor2_4 _48677_ (.A(_18064_),
    .B(_18070_),
    .Y(_18071_));
 sky130_fd_sc_hd__a21o_4 _48678_ (.A1(_18063_),
    .A2(_17667_),
    .B1(_18071_),
    .X(_18072_));
 sky130_fd_sc_hd__and2_4 _48679_ (.A(_18009_),
    .B(_17600_),
    .X(_18073_));
 sky130_fd_sc_hd__a21o_4 _48680_ (.A1(_17916_),
    .A2(_17998_),
    .B1(_18073_),
    .X(_18074_));
 sky130_fd_sc_hd__and2_4 _48681_ (.A(_18005_),
    .B(_17753_),
    .X(_18075_));
 sky130_fd_sc_hd__a21o_4 _48682_ (.A1(_17605_),
    .A2(_18010_),
    .B1(_18075_),
    .X(_18076_));
 sky130_fd_sc_hd__and2_4 _48683_ (.A(_18076_),
    .B(_17718_),
    .X(_18077_));
 sky130_fd_sc_hd__a21o_4 _48684_ (.A1(_17711_),
    .A2(_18074_),
    .B1(_18077_),
    .X(_18078_));
 sky130_fd_sc_hd__nand2_4 _48685_ (.A(_18078_),
    .B(_18015_),
    .Y(_18079_));
 sky130_fd_sc_hd__o21a_4 _48686_ (.A1(_18018_),
    .A2(_17618_),
    .B1(_17630_),
    .X(_18080_));
 sky130_fd_sc_hd__a21o_4 _48687_ (.A1(_17901_),
    .A2(_18006_),
    .B1(_18080_),
    .X(_18081_));
 sky130_fd_sc_hd__nand2_4 _48688_ (.A(_18081_),
    .B(_18021_),
    .Y(_18082_));
 sky130_fd_sc_hd__nand2_4 _48689_ (.A(_18017_),
    .B(_17851_),
    .Y(_18083_));
 sky130_fd_sc_hd__nand2_4 _48690_ (.A(_18024_),
    .B(_17905_),
    .Y(_18084_));
 sky130_fd_sc_hd__a21o_4 _48691_ (.A1(_18083_),
    .A2(_18084_),
    .B1(_17668_),
    .X(_18085_));
 sky130_fd_sc_hd__a21o_4 _48692_ (.A1(_18082_),
    .A2(_18085_),
    .B1(_17979_),
    .X(_18086_));
 sky130_fd_sc_hd__a21oi_4 _48693_ (.A1(_18079_),
    .A2(_18086_),
    .B1(_18056_),
    .Y(_18087_));
 sky130_fd_sc_hd__a21o_4 _48694_ (.A1(_17862_),
    .A2(_18072_),
    .B1(_18087_),
    .X(_24342_));
 sky130_fd_sc_hd__buf_1 _48695_ (.A(_17548_),
    .X(_18088_));
 sky130_fd_sc_hd__and2_4 _48696_ (.A(_17948_),
    .B(_17704_),
    .X(_18089_));
 sky130_fd_sc_hd__a21o_4 _48697_ (.A1(_17798_),
    .A2(_17940_),
    .B1(_18089_),
    .X(_18090_));
 sky130_fd_sc_hd__nor3_4 _48698_ (.A(_17590_),
    .B(_05413_),
    .C(_18067_),
    .Y(_18091_));
 sky130_fd_sc_hd__a21oi_4 _48699_ (.A1(_17936_),
    .A2(_21143_),
    .B1(_18091_),
    .Y(_18092_));
 sky130_fd_sc_hd__nor2_4 _48700_ (.A(_18064_),
    .B(_18092_),
    .Y(_18093_));
 sky130_fd_sc_hd__a21o_4 _48701_ (.A1(_18090_),
    .A2(_17667_),
    .B1(_18093_),
    .X(_18094_));
 sky130_fd_sc_hd__and2_4 _48702_ (.A(_17961_),
    .B(_17718_),
    .X(_18095_));
 sky130_fd_sc_hd__a21o_4 _48703_ (.A1(_17957_),
    .A2(_17952_),
    .B1(_18095_),
    .X(_18096_));
 sky130_fd_sc_hd__nand2_4 _48704_ (.A(_18096_),
    .B(_18015_),
    .Y(_18097_));
 sky130_fd_sc_hd__nand2_4 _48705_ (.A(_17965_),
    .B(_18021_),
    .Y(_18098_));
 sky130_fd_sc_hd__nand2_4 _48706_ (.A(_17972_),
    .B(_17881_),
    .Y(_18099_));
 sky130_fd_sc_hd__a21o_4 _48707_ (.A1(_18098_),
    .A2(_18099_),
    .B1(_17680_),
    .X(_18100_));
 sky130_fd_sc_hd__a21oi_4 _48708_ (.A1(_18097_),
    .A2(_18100_),
    .B1(_18056_),
    .Y(_18101_));
 sky130_fd_sc_hd__a21o_4 _48709_ (.A1(_18088_),
    .A2(_18094_),
    .B1(_18101_),
    .X(_24343_));
 sky130_fd_sc_hd__and2_4 _48710_ (.A(_17985_),
    .B(_17689_),
    .X(_18102_));
 sky130_fd_sc_hd__a21o_4 _48711_ (.A1(_17683_),
    .A2(_17996_),
    .B1(_18102_),
    .X(_18103_));
 sky130_fd_sc_hd__a21oi_4 _48712_ (.A1(_17990_),
    .A2(_21143_),
    .B1(_18091_),
    .Y(_18104_));
 sky130_fd_sc_hd__nor2_4 _48713_ (.A(_18064_),
    .B(_18104_),
    .Y(_18105_));
 sky130_fd_sc_hd__a21o_4 _48714_ (.A1(_18103_),
    .A2(_17807_),
    .B1(_18105_),
    .X(_18106_));
 sky130_fd_sc_hd__and2_4 _48715_ (.A(_18012_),
    .B(_17718_),
    .X(_18107_));
 sky130_fd_sc_hd__a21o_4 _48716_ (.A1(_17957_),
    .A2(_18000_),
    .B1(_18107_),
    .X(_18108_));
 sky130_fd_sc_hd__buf_1 _48717_ (.A(_17846_),
    .X(_18109_));
 sky130_fd_sc_hd__nand2_4 _48718_ (.A(_18108_),
    .B(_18109_),
    .Y(_18110_));
 sky130_fd_sc_hd__nand2_4 _48719_ (.A(_18008_),
    .B(_17711_),
    .Y(_18111_));
 sky130_fd_sc_hd__nand2_4 _48720_ (.A(_18020_),
    .B(_17881_),
    .Y(_18112_));
 sky130_fd_sc_hd__a21o_4 _48721_ (.A1(_18111_),
    .A2(_18112_),
    .B1(_17680_),
    .X(_18113_));
 sky130_fd_sc_hd__a21oi_4 _48722_ (.A1(_18110_),
    .A2(_18113_),
    .B1(_18056_),
    .Y(_18114_));
 sky130_fd_sc_hd__a21o_4 _48723_ (.A1(_18088_),
    .A2(_18106_),
    .B1(_18114_),
    .X(_24344_));
 sky130_fd_sc_hd__and2_4 _48724_ (.A(_18037_),
    .B(_17704_),
    .X(_18115_));
 sky130_fd_sc_hd__a21o_4 _48725_ (.A1(_17798_),
    .A2(_18030_),
    .B1(_18115_),
    .X(_18116_));
 sky130_vsdinv _48726_ (.A(_18091_),
    .Y(_18117_));
 sky130_fd_sc_hd__o21a_4 _48727_ (.A1(_17749_),
    .A2(_18031_),
    .B1(_18117_),
    .X(_18118_));
 sky130_fd_sc_hd__nor2_4 _48728_ (.A(_18064_),
    .B(_18118_),
    .Y(_18119_));
 sky130_fd_sc_hd__a21o_4 _48729_ (.A1(_18116_),
    .A2(_17807_),
    .B1(_18119_),
    .X(_18120_));
 sky130_fd_sc_hd__and2_4 _48730_ (.A(_18043_),
    .B(_17768_),
    .X(_18121_));
 sky130_fd_sc_hd__a21o_4 _48731_ (.A1(_17957_),
    .A2(_18035_),
    .B1(_18121_),
    .X(_18122_));
 sky130_fd_sc_hd__nand2_4 _48732_ (.A(_18122_),
    .B(_18109_),
    .Y(_18123_));
 sky130_fd_sc_hd__nand2_4 _48733_ (.A(_18045_),
    .B(_17711_),
    .Y(_18124_));
 sky130_fd_sc_hd__nand2_4 _48734_ (.A(_18050_),
    .B(_17881_),
    .Y(_18125_));
 sky130_fd_sc_hd__a21o_4 _48735_ (.A1(_18124_),
    .A2(_18125_),
    .B1(_17680_),
    .X(_18126_));
 sky130_fd_sc_hd__buf_1 _48736_ (.A(_17794_),
    .X(_18127_));
 sky130_fd_sc_hd__a21oi_4 _48737_ (.A1(_18123_),
    .A2(_18126_),
    .B1(_18127_),
    .Y(_18128_));
 sky130_fd_sc_hd__a21o_4 _48738_ (.A1(_18088_),
    .A2(_18120_),
    .B1(_18128_),
    .X(_24345_));
 sky130_fd_sc_hd__buf_1 _48739_ (.A(_17644_),
    .X(_18129_));
 sky130_fd_sc_hd__and2_4 _48740_ (.A(_18061_),
    .B(_01491_),
    .X(_18130_));
 sky130_fd_sc_hd__a21o_4 _48741_ (.A1(_17669_),
    .A2(_18066_),
    .B1(_18130_),
    .X(_18131_));
 sky130_fd_sc_hd__buf_1 _48742_ (.A(_18067_),
    .X(_18132_));
 sky130_fd_sc_hd__a21boi_4 _48743_ (.A1(_05595_),
    .A2(_17683_),
    .B1_N(_18132_),
    .Y(_18133_));
 sky130_fd_sc_hd__nor3_4 _48744_ (.A(_17758_),
    .B(_05414_),
    .C(_18133_),
    .Y(_18134_));
 sky130_fd_sc_hd__a21oi_4 _48745_ (.A1(_18131_),
    .A2(_01518_),
    .B1(_18134_),
    .Y(_18135_));
 sky130_fd_sc_hd__nand2_4 _48746_ (.A(_18076_),
    .B(_17669_),
    .Y(_18136_));
 sky130_fd_sc_hd__nand2_4 _48747_ (.A(_18081_),
    .B(_01492_),
    .Y(_18137_));
 sky130_fd_sc_hd__a21oi_4 _48748_ (.A1(_18136_),
    .A2(_18137_),
    .B1(_17723_),
    .Y(_18138_));
 sky130_fd_sc_hd__and2_4 _48749_ (.A(_18074_),
    .B(_17735_),
    .X(_18139_));
 sky130_fd_sc_hd__and2_4 _48750_ (.A(_18059_),
    .B(_17749_),
    .X(_18140_));
 sky130_fd_sc_hd__o21a_4 _48751_ (.A1(_18139_),
    .A2(_18140_),
    .B1(_17625_),
    .X(_18141_));
 sky130_fd_sc_hd__o21ai_4 _48752_ (.A1(_18138_),
    .A2(_18141_),
    .B1(_17595_),
    .Y(_18142_));
 sky130_fd_sc_hd__o21ai_4 _48753_ (.A1(_18129_),
    .A2(_18135_),
    .B1(_18142_),
    .Y(_24346_));
 sky130_fd_sc_hd__nor3_4 _48754_ (.A(_24249_),
    .B(_05414_),
    .C(_18067_),
    .Y(_18143_));
 sky130_fd_sc_hd__a21oi_4 _48755_ (.A1(_17942_),
    .A2(_01518_),
    .B1(_18143_),
    .Y(_18144_));
 sky130_fd_sc_hd__nand2_4 _48756_ (.A(_17954_),
    .B(_17831_),
    .Y(_18145_));
 sky130_fd_sc_hd__nand2_4 _48757_ (.A(_17967_),
    .B(_17894_),
    .Y(_18146_));
 sky130_fd_sc_hd__a21o_4 _48758_ (.A1(_18145_),
    .A2(_18146_),
    .B1(_17760_),
    .X(_18147_));
 sky130_fd_sc_hd__o21ai_4 _48759_ (.A1(_18129_),
    .A2(_18144_),
    .B1(_18147_),
    .Y(_24347_));
 sky130_fd_sc_hd__a21oi_4 _48760_ (.A1(_17992_),
    .A2(_17709_),
    .B1(_18143_),
    .Y(_18148_));
 sky130_fd_sc_hd__nand2_4 _48761_ (.A(_18002_),
    .B(_03459_),
    .Y(_18149_));
 sky130_fd_sc_hd__nand2_4 _48762_ (.A(_18014_),
    .B(_17894_),
    .Y(_18150_));
 sky130_fd_sc_hd__a21o_4 _48763_ (.A1(_18149_),
    .A2(_18150_),
    .B1(_17760_),
    .X(_18151_));
 sky130_fd_sc_hd__o21ai_4 _48764_ (.A1(_18129_),
    .A2(_18148_),
    .B1(_18151_),
    .Y(_24348_));
 sky130_fd_sc_hd__a21oi_4 _48765_ (.A1(_18033_),
    .A2(_17709_),
    .B1(_18143_),
    .Y(_18152_));
 sky130_fd_sc_hd__nand2_4 _48766_ (.A(_18039_),
    .B(_03459_),
    .Y(_18153_));
 sky130_fd_sc_hd__nand2_4 _48767_ (.A(_18047_),
    .B(_17894_),
    .Y(_18154_));
 sky130_fd_sc_hd__a21o_4 _48768_ (.A1(_18153_),
    .A2(_18154_),
    .B1(_17760_),
    .X(_18155_));
 sky130_fd_sc_hd__o21ai_4 _48769_ (.A1(_18129_),
    .A2(_18152_),
    .B1(_18155_),
    .Y(_24318_));
 sky130_fd_sc_hd__buf_1 _48770_ (.A(_17641_),
    .X(_18156_));
 sky130_vsdinv _48771_ (.A(_18143_),
    .Y(_18157_));
 sky130_fd_sc_hd__o21ai_4 _48772_ (.A1(_18156_),
    .A2(_18070_),
    .B1(_18157_),
    .Y(_18158_));
 sky130_fd_sc_hd__nand2_4 _48773_ (.A(_18063_),
    .B(_18109_),
    .Y(_18159_));
 sky130_fd_sc_hd__buf_1 _48774_ (.A(_17731_),
    .X(_18160_));
 sky130_fd_sc_hd__nand2_4 _48775_ (.A(_18078_),
    .B(_18160_),
    .Y(_18161_));
 sky130_fd_sc_hd__a21oi_4 _48776_ (.A1(_18159_),
    .A2(_18161_),
    .B1(_18127_),
    .Y(_18162_));
 sky130_fd_sc_hd__a21o_4 _48777_ (.A1(_18088_),
    .A2(_18158_),
    .B1(_18162_),
    .X(_24319_));
 sky130_fd_sc_hd__o21ai_4 _48778_ (.A1(_18156_),
    .A2(_18092_),
    .B1(_18157_),
    .Y(_18163_));
 sky130_fd_sc_hd__nand2_4 _48779_ (.A(_18090_),
    .B(_18109_),
    .Y(_18164_));
 sky130_fd_sc_hd__nand2_4 _48780_ (.A(_18096_),
    .B(_18160_),
    .Y(_18165_));
 sky130_fd_sc_hd__a21oi_4 _48781_ (.A1(_18164_),
    .A2(_18165_),
    .B1(_18127_),
    .Y(_18166_));
 sky130_fd_sc_hd__a21o_4 _48782_ (.A1(_17886_),
    .A2(_18163_),
    .B1(_18166_),
    .X(_24320_));
 sky130_fd_sc_hd__o21ai_4 _48783_ (.A1(_18156_),
    .A2(_18104_),
    .B1(_18157_),
    .Y(_18167_));
 sky130_fd_sc_hd__nand2_4 _48784_ (.A(_18103_),
    .B(_17831_),
    .Y(_18168_));
 sky130_fd_sc_hd__nand2_4 _48785_ (.A(_18108_),
    .B(_18160_),
    .Y(_18169_));
 sky130_fd_sc_hd__a21oi_4 _48786_ (.A1(_18168_),
    .A2(_18169_),
    .B1(_18127_),
    .Y(_18170_));
 sky130_fd_sc_hd__a21o_4 _48787_ (.A1(_17886_),
    .A2(_18167_),
    .B1(_18170_),
    .X(_24321_));
 sky130_fd_sc_hd__o21ai_4 _48788_ (.A1(_18156_),
    .A2(_18118_),
    .B1(_18157_),
    .Y(_18171_));
 sky130_fd_sc_hd__nand2_4 _48789_ (.A(_18116_),
    .B(_17831_),
    .Y(_18172_));
 sky130_fd_sc_hd__nand2_4 _48790_ (.A(_18122_),
    .B(_18160_),
    .Y(_18173_));
 sky130_fd_sc_hd__a21oi_4 _48791_ (.A1(_18172_),
    .A2(_18173_),
    .B1(_17809_),
    .Y(_18174_));
 sky130_fd_sc_hd__a21o_4 _48792_ (.A1(_17886_),
    .A2(_18171_),
    .B1(_18174_),
    .X(_24322_));
 sky130_fd_sc_hd__a211o_4 _48793_ (.A1(_03450_),
    .A2(_18066_),
    .B1(_17553_),
    .C1(_18130_),
    .X(_18175_));
 sky130_fd_sc_hd__a211o_4 _48794_ (.A1(_21144_),
    .A2(_18074_),
    .B1(_17557_),
    .C1(_18140_),
    .X(_18176_));
 sky130_fd_sc_hd__nand3_4 _48795_ (.A(_18175_),
    .B(_18176_),
    .C(_17555_),
    .Y(_18177_));
 sky130_fd_sc_hd__nand2_4 _48796_ (.A(_03468_),
    .B(_21906_),
    .Y(_18178_));
 sky130_fd_sc_hd__a21o_4 _48797_ (.A1(_05616_),
    .A2(_18132_),
    .B1(_18178_),
    .X(_18179_));
 sky130_fd_sc_hd__nand2_4 _48798_ (.A(_18177_),
    .B(_18179_),
    .Y(_24323_));
 sky130_fd_sc_hd__nor3_4 _48799_ (.A(_21166_),
    .B(_05414_),
    .C(_18132_),
    .Y(_18180_));
 sky130_fd_sc_hd__buf_1 _48800_ (.A(_18180_),
    .X(_18181_));
 sky130_fd_sc_hd__buf_1 _48801_ (.A(_18181_),
    .X(_18182_));
 sky130_fd_sc_hd__a21o_4 _48802_ (.A1(_17956_),
    .A2(_21169_),
    .B1(_18182_),
    .X(_24324_));
 sky130_fd_sc_hd__a21o_4 _48803_ (.A1(_18004_),
    .A2(_21169_),
    .B1(_18182_),
    .X(_24325_));
 sky130_fd_sc_hd__a21o_4 _48804_ (.A1(_18041_),
    .A2(_21169_),
    .B1(_18182_),
    .X(_24326_));
 sky130_fd_sc_hd__buf_1 _48805_ (.A(_17644_),
    .X(_18183_));
 sky130_fd_sc_hd__a21o_4 _48806_ (.A1(_18072_),
    .A2(_18183_),
    .B1(_18182_),
    .X(_24327_));
 sky130_fd_sc_hd__buf_1 _48807_ (.A(_18180_),
    .X(_18184_));
 sky130_fd_sc_hd__a21o_4 _48808_ (.A1(_18094_),
    .A2(_18183_),
    .B1(_18184_),
    .X(_24329_));
 sky130_fd_sc_hd__a21o_4 _48809_ (.A1(_18106_),
    .A2(_18183_),
    .B1(_18184_),
    .X(_24330_));
 sky130_fd_sc_hd__a21o_4 _48810_ (.A1(_18120_),
    .A2(_18183_),
    .B1(_18184_),
    .X(_24331_));
 sky130_vsdinv _48811_ (.A(_18132_),
    .Y(_18185_));
 sky130_fd_sc_hd__nand3_4 _48812_ (.A(_18185_),
    .B(_17772_),
    .C(_21906_),
    .Y(_18186_));
 sky130_fd_sc_hd__o21ai_4 _48813_ (.A1(_17783_),
    .A2(_18135_),
    .B1(_18186_),
    .Y(_24332_));
 sky130_fd_sc_hd__o21ai_4 _48814_ (.A1(_17783_),
    .A2(_18144_),
    .B1(_18186_),
    .Y(_24333_));
 sky130_fd_sc_hd__o21ai_4 _48815_ (.A1(_17783_),
    .A2(_18148_),
    .B1(_18186_),
    .Y(_24334_));
 sky130_fd_sc_hd__o21ai_4 _48816_ (.A1(_17549_),
    .A2(_18152_),
    .B1(_18186_),
    .Y(_24335_));
 sky130_fd_sc_hd__buf_1 _48817_ (.A(_21168_),
    .X(_18187_));
 sky130_fd_sc_hd__a21o_4 _48818_ (.A1(_18158_),
    .A2(_18187_),
    .B1(_18184_),
    .X(_24336_));
 sky130_fd_sc_hd__a21o_4 _48819_ (.A1(_18163_),
    .A2(_18187_),
    .B1(_18181_),
    .X(_24337_));
 sky130_fd_sc_hd__a21o_4 _48820_ (.A1(_18167_),
    .A2(_18187_),
    .B1(_18181_),
    .X(_24338_));
 sky130_fd_sc_hd__a21o_4 _48821_ (.A1(_18171_),
    .A2(_18187_),
    .B1(_18181_),
    .X(_24340_));
 sky130_fd_sc_hd__o21a_4 _48822_ (.A1(_18185_),
    .A2(_05626_),
    .B1(_21906_),
    .X(_24341_));
 sky130_fd_sc_hd__conb_1 _48823_ (.LO(mem_la_addr[0]));
 sky130_fd_sc_hd__conb_1 _48824_ (.LO(mem_la_addr[1]));
 sky130_fd_sc_hd__conb_1 _48825_ (.LO(trace_valid));
 sky130_fd_sc_hd__buf_2 _48826_ (.A(mem_la_wdata[0]),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__buf_2 _48827_ (.A(mem_la_wdata[1]),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__buf_2 _48828_ (.A(mem_la_wdata[2]),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__buf_2 _48829_ (.A(mem_la_wdata[3]),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__buf_2 _48830_ (.A(mem_la_wdata[4]),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__buf_2 _48831_ (.A(mem_la_wdata[5]),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__buf_2 _48832_ (.A(mem_la_wdata[6]),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__buf_2 _48833_ (.A(mem_la_wdata[7]),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__buf_2 _48834_ (.A(zero_),
    .X(trace_data[0]));
 sky130_fd_sc_hd__buf_2 _48835_ (.A(zero_),
    .X(trace_data[1]));
 sky130_fd_sc_hd__buf_2 _48836_ (.A(zero_),
    .X(trace_data[2]));
 sky130_fd_sc_hd__buf_2 _48837_ (.A(zero_),
    .X(trace_data[3]));
 sky130_fd_sc_hd__buf_2 _48838_ (.A(zero_),
    .X(trace_data[4]));
 sky130_fd_sc_hd__buf_2 _48839_ (.A(zero_),
    .X(trace_data[5]));
 sky130_fd_sc_hd__buf_2 _48840_ (.A(zero_),
    .X(trace_data[6]));
 sky130_fd_sc_hd__buf_2 _48841_ (.A(zero_),
    .X(trace_data[7]));
 sky130_fd_sc_hd__buf_2 _48842_ (.A(zero_),
    .X(trace_data[8]));
 sky130_fd_sc_hd__buf_2 _48843_ (.A(zero_),
    .X(trace_data[9]));
 sky130_fd_sc_hd__buf_2 _48844_ (.A(zero_),
    .X(trace_data[10]));
 sky130_fd_sc_hd__buf_2 _48845_ (.A(zero_),
    .X(trace_data[11]));
 sky130_fd_sc_hd__buf_2 _48846_ (.A(zero_),
    .X(trace_data[12]));
 sky130_fd_sc_hd__buf_2 _48847_ (.A(zero_),
    .X(trace_data[13]));
 sky130_fd_sc_hd__buf_2 _48848_ (.A(zero_),
    .X(trace_data[14]));
 sky130_fd_sc_hd__buf_2 _48849_ (.A(zero_),
    .X(trace_data[15]));
 sky130_fd_sc_hd__buf_2 _48850_ (.A(zero_),
    .X(trace_data[16]));
 sky130_fd_sc_hd__buf_2 _48851_ (.A(zero_),
    .X(trace_data[17]));
 sky130_fd_sc_hd__buf_2 _48852_ (.A(zero_),
    .X(trace_data[18]));
 sky130_fd_sc_hd__buf_2 _48853_ (.A(zero_),
    .X(trace_data[19]));
 sky130_fd_sc_hd__buf_2 _48854_ (.A(zero_),
    .X(trace_data[20]));
 sky130_fd_sc_hd__buf_2 _48855_ (.A(zero_),
    .X(trace_data[21]));
 sky130_fd_sc_hd__buf_2 _48856_ (.A(zero_),
    .X(trace_data[22]));
 sky130_fd_sc_hd__buf_2 _48857_ (.A(zero_),
    .X(trace_data[23]));
 sky130_fd_sc_hd__buf_2 _48858_ (.A(zero_),
    .X(trace_data[24]));
 sky130_fd_sc_hd__buf_2 _48859_ (.A(zero_),
    .X(trace_data[25]));
 sky130_fd_sc_hd__buf_2 _48860_ (.A(zero_),
    .X(trace_data[26]));
 sky130_fd_sc_hd__buf_2 _48861_ (.A(zero_),
    .X(trace_data[27]));
 sky130_fd_sc_hd__buf_2 _48862_ (.A(zero_),
    .X(trace_data[28]));
 sky130_fd_sc_hd__buf_2 _48863_ (.A(zero_),
    .X(trace_data[29]));
 sky130_fd_sc_hd__buf_2 _48864_ (.A(zero_),
    .X(trace_data[30]));
 sky130_fd_sc_hd__buf_2 _48865_ (.A(zero_),
    .X(trace_data[31]));
 sky130_fd_sc_hd__buf_2 _48866_ (.A(zero_),
    .X(trace_data[32]));
 sky130_fd_sc_hd__buf_2 _48867_ (.A(zero_),
    .X(trace_data[33]));
 sky130_fd_sc_hd__buf_2 _48868_ (.A(zero_),
    .X(trace_data[34]));
 sky130_fd_sc_hd__buf_2 _48869_ (.A(zero_),
    .X(trace_data[35]));
 sky130_fd_sc_hd__dfxtp_4 _48870_ (.CLK(clk_0_0),
    .D(_00833_),
    .Q(\cpuregs[12][0] ));
 sky130_fd_sc_hd__dfxtp_4 _48871_ (.CLK(clk_0_0),
    .D(_00844_),
    .Q(\cpuregs[12][1] ));
 sky130_fd_sc_hd__dfxtp_4 _48872_ (.CLK(clk_0_0),
    .D(_00855_),
    .Q(\cpuregs[12][2] ));
 sky130_fd_sc_hd__dfxtp_4 _48873_ (.CLK(clk_0_0),
    .D(_00858_),
    .Q(\cpuregs[12][3] ));
 sky130_fd_sc_hd__dfxtp_4 _48874_ (.CLK(clk_0_0),
    .D(_00859_),
    .Q(\cpuregs[12][4] ));
 sky130_fd_sc_hd__dfxtp_4 _48875_ (.CLK(clk_0_0),
    .D(_00860_),
    .Q(\cpuregs[12][5] ));
 sky130_fd_sc_hd__dfxtp_4 _48876_ (.CLK(clk_0_0),
    .D(_00861_),
    .Q(\cpuregs[12][6] ));
 sky130_fd_sc_hd__dfxtp_4 _48877_ (.CLK(clk_0_0),
    .D(_00862_),
    .Q(\cpuregs[12][7] ));
 sky130_fd_sc_hd__dfxtp_4 _48878_ (.CLK(clk_0_0),
    .D(_00863_),
    .Q(\cpuregs[12][8] ));
 sky130_fd_sc_hd__dfxtp_4 _48879_ (.CLK(clk_0_0),
    .D(_00864_),
    .Q(\cpuregs[12][9] ));
 sky130_fd_sc_hd__dfxtp_4 _48880_ (.CLK(clk_0_0),
    .D(_00834_),
    .Q(\cpuregs[12][10] ));
 sky130_fd_sc_hd__dfxtp_4 _48881_ (.CLK(clk_0_0),
    .D(_00835_),
    .Q(\cpuregs[12][11] ));
 sky130_fd_sc_hd__dfxtp_4 _48882_ (.CLK(clk_0_0),
    .D(_00836_),
    .Q(\cpuregs[12][12] ));
 sky130_fd_sc_hd__dfxtp_4 _48883_ (.CLK(clk_0_0),
    .D(_00837_),
    .Q(\cpuregs[12][13] ));
 sky130_fd_sc_hd__dfxtp_4 _48884_ (.CLK(clk_0_0),
    .D(_00838_),
    .Q(\cpuregs[12][14] ));
 sky130_fd_sc_hd__dfxtp_4 _48885_ (.CLK(clk_0_0),
    .D(_00839_),
    .Q(\cpuregs[12][15] ));
 sky130_fd_sc_hd__dfxtp_4 _48886_ (.CLK(clk_0_16),
    .D(_00840_),
    .Q(\cpuregs[12][16] ));
 sky130_fd_sc_hd__dfxtp_4 _48887_ (.CLK(clk_0_16),
    .D(_00841_),
    .Q(\cpuregs[12][17] ));
 sky130_fd_sc_hd__dfxtp_4 _48888_ (.CLK(clk_0_16),
    .D(_00842_),
    .Q(\cpuregs[12][18] ));
 sky130_fd_sc_hd__dfxtp_4 _48889_ (.CLK(clk_0_16),
    .D(_00843_),
    .Q(\cpuregs[12][19] ));
 sky130_fd_sc_hd__dfxtp_4 _48890_ (.CLK(clk_0_16),
    .D(_00845_),
    .Q(\cpuregs[12][20] ));
 sky130_fd_sc_hd__dfxtp_4 _48891_ (.CLK(clk_0_16),
    .D(_00846_),
    .Q(\cpuregs[12][21] ));
 sky130_fd_sc_hd__dfxtp_4 _48892_ (.CLK(clk_0_16),
    .D(_00847_),
    .Q(\cpuregs[12][22] ));
 sky130_fd_sc_hd__dfxtp_4 _48893_ (.CLK(clk_0_16),
    .D(_00848_),
    .Q(\cpuregs[12][23] ));
 sky130_fd_sc_hd__dfxtp_4 _48894_ (.CLK(clk_0_16),
    .D(_00849_),
    .Q(\cpuregs[12][24] ));
 sky130_fd_sc_hd__dfxtp_4 _48895_ (.CLK(clk_0_16),
    .D(_00850_),
    .Q(\cpuregs[12][25] ));
 sky130_fd_sc_hd__dfxtp_4 _48896_ (.CLK(clk_0_16),
    .D(_00851_),
    .Q(\cpuregs[12][26] ));
 sky130_fd_sc_hd__dfxtp_4 _48897_ (.CLK(clk_0_16),
    .D(_00852_),
    .Q(\cpuregs[12][27] ));
 sky130_fd_sc_hd__dfxtp_4 _48898_ (.CLK(clk_0_16),
    .D(_00853_),
    .Q(\cpuregs[12][28] ));
 sky130_fd_sc_hd__dfxtp_4 _48899_ (.CLK(clk_0_16),
    .D(_00854_),
    .Q(\cpuregs[12][29] ));
 sky130_fd_sc_hd__dfxtp_4 _48900_ (.CLK(clk_0_16),
    .D(_00856_),
    .Q(\cpuregs[12][30] ));
 sky130_fd_sc_hd__dfxtp_4 _48901_ (.CLK(clk_0_16),
    .D(_00857_),
    .Q(\cpuregs[12][31] ));
 sky130_fd_sc_hd__dfxtp_4 _48902_ (.CLK(clk_0_32),
    .D(_00666_),
    .Q(\mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_4 _48903_ (.CLK(clk_0_32),
    .D(_00667_),
    .Q(\mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_4 _48904_ (.CLK(clk_0_32),
    .D(_00668_),
    .Q(\mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_4 _48905_ (.CLK(clk_0_32),
    .D(_01345_),
    .Q(\cpuregs[9][0] ));
 sky130_fd_sc_hd__dfxtp_4 _48906_ (.CLK(clk_0_32),
    .D(_01356_),
    .Q(\cpuregs[9][1] ));
 sky130_fd_sc_hd__dfxtp_4 _48907_ (.CLK(clk_0_32),
    .D(_01367_),
    .Q(\cpuregs[9][2] ));
 sky130_fd_sc_hd__dfxtp_4 _48908_ (.CLK(clk_0_32),
    .D(_01370_),
    .Q(\cpuregs[9][3] ));
 sky130_fd_sc_hd__dfxtp_4 _48909_ (.CLK(clk_0_32),
    .D(_01371_),
    .Q(\cpuregs[9][4] ));
 sky130_fd_sc_hd__dfxtp_4 _48910_ (.CLK(clk_0_32),
    .D(_01372_),
    .Q(\cpuregs[9][5] ));
 sky130_fd_sc_hd__dfxtp_4 _48911_ (.CLK(clk_0_32),
    .D(_01373_),
    .Q(\cpuregs[9][6] ));
 sky130_fd_sc_hd__dfxtp_4 _48912_ (.CLK(clk_0_32),
    .D(_01374_),
    .Q(\cpuregs[9][7] ));
 sky130_fd_sc_hd__dfxtp_4 _48913_ (.CLK(clk_0_32),
    .D(_01375_),
    .Q(\cpuregs[9][8] ));
 sky130_fd_sc_hd__dfxtp_4 _48914_ (.CLK(clk_0_32),
    .D(_01376_),
    .Q(\cpuregs[9][9] ));
 sky130_fd_sc_hd__dfxtp_4 _48915_ (.CLK(clk_0_32),
    .D(_01346_),
    .Q(\cpuregs[9][10] ));
 sky130_fd_sc_hd__dfxtp_4 _48916_ (.CLK(clk_0_32),
    .D(_01347_),
    .Q(\cpuregs[9][11] ));
 sky130_fd_sc_hd__dfxtp_4 _48917_ (.CLK(clk_0_32),
    .D(_01348_),
    .Q(\cpuregs[9][12] ));
 sky130_fd_sc_hd__dfxtp_4 _48918_ (.CLK(clk_0_48),
    .D(_01349_),
    .Q(\cpuregs[9][13] ));
 sky130_fd_sc_hd__dfxtp_4 _48919_ (.CLK(clk_0_48),
    .D(_01350_),
    .Q(\cpuregs[9][14] ));
 sky130_fd_sc_hd__dfxtp_4 _48920_ (.CLK(clk_0_48),
    .D(_01351_),
    .Q(\cpuregs[9][15] ));
 sky130_fd_sc_hd__dfxtp_4 _48921_ (.CLK(clk_0_48),
    .D(_01352_),
    .Q(\cpuregs[9][16] ));
 sky130_fd_sc_hd__dfxtp_4 _48922_ (.CLK(clk_0_48),
    .D(_01353_),
    .Q(\cpuregs[9][17] ));
 sky130_fd_sc_hd__dfxtp_4 _48923_ (.CLK(clk_0_48),
    .D(_01354_),
    .Q(\cpuregs[9][18] ));
 sky130_fd_sc_hd__dfxtp_4 _48924_ (.CLK(clk_0_48),
    .D(_01355_),
    .Q(\cpuregs[9][19] ));
 sky130_fd_sc_hd__dfxtp_4 _48925_ (.CLK(clk_0_48),
    .D(_01357_),
    .Q(\cpuregs[9][20] ));
 sky130_fd_sc_hd__dfxtp_4 _48926_ (.CLK(clk_0_48),
    .D(_01358_),
    .Q(\cpuregs[9][21] ));
 sky130_fd_sc_hd__dfxtp_4 _48927_ (.CLK(clk_0_48),
    .D(_01359_),
    .Q(\cpuregs[9][22] ));
 sky130_fd_sc_hd__dfxtp_4 _48928_ (.CLK(clk_0_48),
    .D(_01360_),
    .Q(\cpuregs[9][23] ));
 sky130_fd_sc_hd__dfxtp_4 _48929_ (.CLK(clk_0_48),
    .D(_01361_),
    .Q(\cpuregs[9][24] ));
 sky130_fd_sc_hd__dfxtp_4 _48930_ (.CLK(clk_0_48),
    .D(_01362_),
    .Q(\cpuregs[9][25] ));
 sky130_fd_sc_hd__dfxtp_4 _48931_ (.CLK(clk_0_48),
    .D(_01363_),
    .Q(\cpuregs[9][26] ));
 sky130_fd_sc_hd__dfxtp_4 _48932_ (.CLK(clk_0_48),
    .D(_01364_),
    .Q(\cpuregs[9][27] ));
 sky130_fd_sc_hd__dfxtp_4 _48933_ (.CLK(clk_0_48),
    .D(_01365_),
    .Q(\cpuregs[9][28] ));
 sky130_fd_sc_hd__dfxtp_4 _48934_ (.CLK(clk_0_64),
    .D(_01366_),
    .Q(\cpuregs[9][29] ));
 sky130_fd_sc_hd__dfxtp_4 _48935_ (.CLK(clk_0_64),
    .D(_01368_),
    .Q(\cpuregs[9][30] ));
 sky130_fd_sc_hd__dfxtp_4 _48936_ (.CLK(clk_0_64),
    .D(_01369_),
    .Q(\cpuregs[9][31] ));
 sky130_fd_sc_hd__dfxtp_4 _48937_ (.CLK(clk_0_64),
    .D(_00865_),
    .Q(\cpuregs[13][0] ));
 sky130_fd_sc_hd__dfxtp_4 _48938_ (.CLK(clk_0_64),
    .D(_00876_),
    .Q(\cpuregs[13][1] ));
 sky130_fd_sc_hd__dfxtp_4 _48939_ (.CLK(clk_0_64),
    .D(_00887_),
    .Q(\cpuregs[13][2] ));
 sky130_fd_sc_hd__dfxtp_4 _48940_ (.CLK(clk_0_64),
    .D(_00890_),
    .Q(\cpuregs[13][3] ));
 sky130_fd_sc_hd__dfxtp_4 _48941_ (.CLK(clk_0_64),
    .D(_00891_),
    .Q(\cpuregs[13][4] ));
 sky130_fd_sc_hd__dfxtp_4 _48942_ (.CLK(clk_0_64),
    .D(_00892_),
    .Q(\cpuregs[13][5] ));
 sky130_fd_sc_hd__dfxtp_4 _48943_ (.CLK(clk_0_64),
    .D(_00893_),
    .Q(\cpuregs[13][6] ));
 sky130_fd_sc_hd__dfxtp_4 _48944_ (.CLK(clk_0_64),
    .D(_00894_),
    .Q(\cpuregs[13][7] ));
 sky130_fd_sc_hd__dfxtp_4 _48945_ (.CLK(clk_0_64),
    .D(_00895_),
    .Q(\cpuregs[13][8] ));
 sky130_fd_sc_hd__dfxtp_4 _48946_ (.CLK(clk_0_64),
    .D(_00896_),
    .Q(\cpuregs[13][9] ));
 sky130_fd_sc_hd__dfxtp_4 _48947_ (.CLK(clk_0_64),
    .D(_00866_),
    .Q(\cpuregs[13][10] ));
 sky130_fd_sc_hd__dfxtp_4 _48948_ (.CLK(clk_0_64),
    .D(_00867_),
    .Q(\cpuregs[13][11] ));
 sky130_fd_sc_hd__dfxtp_4 _48949_ (.CLK(clk_0_64),
    .D(_00868_),
    .Q(\cpuregs[13][12] ));
 sky130_fd_sc_hd__dfxtp_4 _48950_ (.CLK(clk_0_80),
    .D(_00869_),
    .Q(\cpuregs[13][13] ));
 sky130_fd_sc_hd__dfxtp_4 _48951_ (.CLK(clk_0_80),
    .D(_00870_),
    .Q(\cpuregs[13][14] ));
 sky130_fd_sc_hd__dfxtp_4 _48952_ (.CLK(clk_0_80),
    .D(_00871_),
    .Q(\cpuregs[13][15] ));
 sky130_fd_sc_hd__dfxtp_4 _48953_ (.CLK(clk_0_80),
    .D(_00872_),
    .Q(\cpuregs[13][16] ));
 sky130_fd_sc_hd__dfxtp_4 _48954_ (.CLK(clk_0_80),
    .D(_00873_),
    .Q(\cpuregs[13][17] ));
 sky130_fd_sc_hd__dfxtp_4 _48955_ (.CLK(clk_0_80),
    .D(_00874_),
    .Q(\cpuregs[13][18] ));
 sky130_fd_sc_hd__dfxtp_4 _48956_ (.CLK(clk_0_80),
    .D(_00875_),
    .Q(\cpuregs[13][19] ));
 sky130_fd_sc_hd__dfxtp_4 _48957_ (.CLK(clk_0_80),
    .D(_00877_),
    .Q(\cpuregs[13][20] ));
 sky130_fd_sc_hd__dfxtp_4 _48958_ (.CLK(clk_0_80),
    .D(_00878_),
    .Q(\cpuregs[13][21] ));
 sky130_fd_sc_hd__dfxtp_4 _48959_ (.CLK(clk_0_80),
    .D(_00879_),
    .Q(\cpuregs[13][22] ));
 sky130_fd_sc_hd__dfxtp_4 _48960_ (.CLK(clk_0_80),
    .D(_00880_),
    .Q(\cpuregs[13][23] ));
 sky130_fd_sc_hd__dfxtp_4 _48961_ (.CLK(clk_0_80),
    .D(_00881_),
    .Q(\cpuregs[13][24] ));
 sky130_fd_sc_hd__dfxtp_4 _48962_ (.CLK(clk_0_80),
    .D(_00882_),
    .Q(\cpuregs[13][25] ));
 sky130_fd_sc_hd__dfxtp_4 _48963_ (.CLK(clk_0_80),
    .D(_00883_),
    .Q(\cpuregs[13][26] ));
 sky130_fd_sc_hd__dfxtp_4 _48964_ (.CLK(clk_0_80),
    .D(_00884_),
    .Q(\cpuregs[13][27] ));
 sky130_fd_sc_hd__dfxtp_4 _48965_ (.CLK(clk_0_80),
    .D(_00885_),
    .Q(\cpuregs[13][28] ));
 sky130_fd_sc_hd__dfxtp_4 _48966_ (.CLK(clk_0_96),
    .D(_00886_),
    .Q(\cpuregs[13][29] ));
 sky130_fd_sc_hd__dfxtp_4 _48967_ (.CLK(clk_0_96),
    .D(_00888_),
    .Q(\cpuregs[13][30] ));
 sky130_fd_sc_hd__dfxtp_4 _48968_ (.CLK(clk_0_96),
    .D(_00889_),
    .Q(\cpuregs[13][31] ));
 sky130_fd_sc_hd__dfxtp_4 _48969_ (.CLK(clk_0_96),
    .D(_00897_),
    .Q(\cpuregs[14][0] ));
 sky130_fd_sc_hd__dfxtp_4 _48970_ (.CLK(clk_0_96),
    .D(_00908_),
    .Q(\cpuregs[14][1] ));
 sky130_fd_sc_hd__dfxtp_4 _48971_ (.CLK(clk_0_96),
    .D(_00919_),
    .Q(\cpuregs[14][2] ));
 sky130_fd_sc_hd__dfxtp_4 _48972_ (.CLK(clk_0_96),
    .D(_00922_),
    .Q(\cpuregs[14][3] ));
 sky130_fd_sc_hd__dfxtp_4 _48973_ (.CLK(clk_0_96),
    .D(_00923_),
    .Q(\cpuregs[14][4] ));
 sky130_fd_sc_hd__dfxtp_4 _48974_ (.CLK(clk_0_96),
    .D(_00924_),
    .Q(\cpuregs[14][5] ));
 sky130_fd_sc_hd__dfxtp_4 _48975_ (.CLK(clk_0_96),
    .D(_00925_),
    .Q(\cpuregs[14][6] ));
 sky130_fd_sc_hd__dfxtp_4 _48976_ (.CLK(clk_0_96),
    .D(_00926_),
    .Q(\cpuregs[14][7] ));
 sky130_fd_sc_hd__dfxtp_4 _48977_ (.CLK(clk_0_96),
    .D(_00927_),
    .Q(\cpuregs[14][8] ));
 sky130_fd_sc_hd__dfxtp_4 _48978_ (.CLK(clk_0_96),
    .D(_00928_),
    .Q(\cpuregs[14][9] ));
 sky130_fd_sc_hd__dfxtp_4 _48979_ (.CLK(clk_0_96),
    .D(_00898_),
    .Q(\cpuregs[14][10] ));
 sky130_fd_sc_hd__dfxtp_4 _48980_ (.CLK(clk_0_96),
    .D(_00899_),
    .Q(\cpuregs[14][11] ));
 sky130_fd_sc_hd__dfxtp_4 _48981_ (.CLK(clk_0_96),
    .D(_00900_),
    .Q(\cpuregs[14][12] ));
 sky130_fd_sc_hd__dfxtp_4 _48982_ (.CLK(clk_0_112),
    .D(_00901_),
    .Q(\cpuregs[14][13] ));
 sky130_fd_sc_hd__dfxtp_4 _48983_ (.CLK(clk_0_112),
    .D(_00902_),
    .Q(\cpuregs[14][14] ));
 sky130_fd_sc_hd__dfxtp_4 _48984_ (.CLK(clk_0_112),
    .D(_00903_),
    .Q(\cpuregs[14][15] ));
 sky130_fd_sc_hd__dfxtp_4 _48985_ (.CLK(clk_0_112),
    .D(_00904_),
    .Q(\cpuregs[14][16] ));
 sky130_fd_sc_hd__dfxtp_4 _48986_ (.CLK(clk_0_112),
    .D(_00905_),
    .Q(\cpuregs[14][17] ));
 sky130_fd_sc_hd__dfxtp_4 _48987_ (.CLK(clk_0_112),
    .D(_00906_),
    .Q(\cpuregs[14][18] ));
 sky130_fd_sc_hd__dfxtp_4 _48988_ (.CLK(clk_0_112),
    .D(_00907_),
    .Q(\cpuregs[14][19] ));
 sky130_fd_sc_hd__dfxtp_4 _48989_ (.CLK(clk_0_112),
    .D(_00909_),
    .Q(\cpuregs[14][20] ));
 sky130_fd_sc_hd__dfxtp_4 _48990_ (.CLK(clk_0_112),
    .D(_00910_),
    .Q(\cpuregs[14][21] ));
 sky130_fd_sc_hd__dfxtp_4 _48991_ (.CLK(clk_0_112),
    .D(_00911_),
    .Q(\cpuregs[14][22] ));
 sky130_fd_sc_hd__dfxtp_4 _48992_ (.CLK(clk_0_112),
    .D(_00912_),
    .Q(\cpuregs[14][23] ));
 sky130_fd_sc_hd__dfxtp_4 _48993_ (.CLK(clk_0_112),
    .D(_00913_),
    .Q(\cpuregs[14][24] ));
 sky130_fd_sc_hd__dfxtp_4 _48994_ (.CLK(clk_0_112),
    .D(_00914_),
    .Q(\cpuregs[14][25] ));
 sky130_fd_sc_hd__dfxtp_4 _48995_ (.CLK(clk_0_112),
    .D(_00915_),
    .Q(\cpuregs[14][26] ));
 sky130_fd_sc_hd__dfxtp_4 _48996_ (.CLK(clk_0_112),
    .D(_00916_),
    .Q(\cpuregs[14][27] ));
 sky130_fd_sc_hd__dfxtp_4 _48997_ (.CLK(clk_0_112),
    .D(_00917_),
    .Q(\cpuregs[14][28] ));
 sky130_fd_sc_hd__dfxtp_4 _48998_ (.CLK(clk_0_128),
    .D(_00918_),
    .Q(\cpuregs[14][29] ));
 sky130_fd_sc_hd__dfxtp_4 _48999_ (.CLK(clk_0_128),
    .D(_00920_),
    .Q(\cpuregs[14][30] ));
 sky130_fd_sc_hd__dfxtp_4 _49000_ (.CLK(clk_0_128),
    .D(_00921_),
    .Q(\cpuregs[14][31] ));
 sky130_fd_sc_hd__dfxtp_4 _49001_ (.CLK(clk_0_128),
    .D(_01153_),
    .Q(\cpuregs[3][0] ));
 sky130_fd_sc_hd__dfxtp_4 _49002_ (.CLK(clk_0_128),
    .D(_01164_),
    .Q(\cpuregs[3][1] ));
 sky130_fd_sc_hd__dfxtp_4 _49003_ (.CLK(clk_0_128),
    .D(_01175_),
    .Q(\cpuregs[3][2] ));
 sky130_fd_sc_hd__dfxtp_4 _49004_ (.CLK(clk_0_128),
    .D(_01178_),
    .Q(\cpuregs[3][3] ));
 sky130_fd_sc_hd__dfxtp_4 _49005_ (.CLK(clk_0_128),
    .D(_01179_),
    .Q(\cpuregs[3][4] ));
 sky130_fd_sc_hd__dfxtp_4 _49006_ (.CLK(clk_0_128),
    .D(_01180_),
    .Q(\cpuregs[3][5] ));
 sky130_fd_sc_hd__dfxtp_4 _49007_ (.CLK(clk_0_128),
    .D(_01181_),
    .Q(\cpuregs[3][6] ));
 sky130_fd_sc_hd__dfxtp_4 _49008_ (.CLK(clk_0_128),
    .D(_01182_),
    .Q(\cpuregs[3][7] ));
 sky130_fd_sc_hd__dfxtp_4 _49009_ (.CLK(clk_0_128),
    .D(_01183_),
    .Q(\cpuregs[3][8] ));
 sky130_fd_sc_hd__dfxtp_4 _49010_ (.CLK(clk_0_128),
    .D(_01184_),
    .Q(\cpuregs[3][9] ));
 sky130_fd_sc_hd__dfxtp_4 _49011_ (.CLK(clk_0_128),
    .D(_01154_),
    .Q(\cpuregs[3][10] ));
 sky130_fd_sc_hd__dfxtp_4 _49012_ (.CLK(clk_0_128),
    .D(_01155_),
    .Q(\cpuregs[3][11] ));
 sky130_fd_sc_hd__dfxtp_4 _49013_ (.CLK(clk_0_128),
    .D(_01156_),
    .Q(\cpuregs[3][12] ));
 sky130_fd_sc_hd__dfxtp_4 _49014_ (.CLK(clk_0_144),
    .D(_01157_),
    .Q(\cpuregs[3][13] ));
 sky130_fd_sc_hd__dfxtp_4 _49015_ (.CLK(clk_0_144),
    .D(_01158_),
    .Q(\cpuregs[3][14] ));
 sky130_fd_sc_hd__dfxtp_4 _49016_ (.CLK(clk_0_144),
    .D(_01159_),
    .Q(\cpuregs[3][15] ));
 sky130_fd_sc_hd__dfxtp_4 _49017_ (.CLK(clk_0_144),
    .D(_01160_),
    .Q(\cpuregs[3][16] ));
 sky130_fd_sc_hd__dfxtp_4 _49018_ (.CLK(clk_0_144),
    .D(_01161_),
    .Q(\cpuregs[3][17] ));
 sky130_fd_sc_hd__dfxtp_4 _49019_ (.CLK(clk_0_144),
    .D(_01162_),
    .Q(\cpuregs[3][18] ));
 sky130_fd_sc_hd__dfxtp_4 _49020_ (.CLK(clk_0_144),
    .D(_01163_),
    .Q(\cpuregs[3][19] ));
 sky130_fd_sc_hd__dfxtp_4 _49021_ (.CLK(clk_0_144),
    .D(_01165_),
    .Q(\cpuregs[3][20] ));
 sky130_fd_sc_hd__dfxtp_4 _49022_ (.CLK(clk_0_144),
    .D(_01166_),
    .Q(\cpuregs[3][21] ));
 sky130_fd_sc_hd__dfxtp_4 _49023_ (.CLK(clk_0_144),
    .D(_01167_),
    .Q(\cpuregs[3][22] ));
 sky130_fd_sc_hd__dfxtp_4 _49024_ (.CLK(clk_0_144),
    .D(_01168_),
    .Q(\cpuregs[3][23] ));
 sky130_fd_sc_hd__dfxtp_4 _49025_ (.CLK(clk_0_144),
    .D(_01169_),
    .Q(\cpuregs[3][24] ));
 sky130_fd_sc_hd__dfxtp_4 _49026_ (.CLK(clk_0_144),
    .D(_01170_),
    .Q(\cpuregs[3][25] ));
 sky130_fd_sc_hd__dfxtp_4 _49027_ (.CLK(clk_0_144),
    .D(_01171_),
    .Q(\cpuregs[3][26] ));
 sky130_fd_sc_hd__dfxtp_4 _49028_ (.CLK(clk_0_144),
    .D(_01172_),
    .Q(\cpuregs[3][27] ));
 sky130_fd_sc_hd__dfxtp_4 _49029_ (.CLK(clk_0_144),
    .D(_01173_),
    .Q(\cpuregs[3][28] ));
 sky130_fd_sc_hd__dfxtp_4 _49030_ (.CLK(clk_0_160),
    .D(_01174_),
    .Q(\cpuregs[3][29] ));
 sky130_fd_sc_hd__dfxtp_4 _49031_ (.CLK(clk_0_160),
    .D(_01176_),
    .Q(\cpuregs[3][30] ));
 sky130_fd_sc_hd__dfxtp_4 _49032_ (.CLK(clk_0_160),
    .D(_01177_),
    .Q(\cpuregs[3][31] ));
 sky130_fd_sc_hd__dfxtp_4 _49033_ (.CLK(clk_0_160),
    .D(_00929_),
    .Q(\cpuregs[15][0] ));
 sky130_fd_sc_hd__dfxtp_4 _49034_ (.CLK(clk_0_160),
    .D(_00940_),
    .Q(\cpuregs[15][1] ));
 sky130_fd_sc_hd__dfxtp_4 _49035_ (.CLK(clk_0_160),
    .D(_00951_),
    .Q(\cpuregs[15][2] ));
 sky130_fd_sc_hd__dfxtp_4 _49036_ (.CLK(clk_0_160),
    .D(_00954_),
    .Q(\cpuregs[15][3] ));
 sky130_fd_sc_hd__dfxtp_4 _49037_ (.CLK(clk_0_160),
    .D(_00955_),
    .Q(\cpuregs[15][4] ));
 sky130_fd_sc_hd__dfxtp_4 _49038_ (.CLK(clk_0_160),
    .D(_00956_),
    .Q(\cpuregs[15][5] ));
 sky130_fd_sc_hd__dfxtp_4 _49039_ (.CLK(clk_0_160),
    .D(_00957_),
    .Q(\cpuregs[15][6] ));
 sky130_fd_sc_hd__dfxtp_4 _49040_ (.CLK(clk_0_160),
    .D(_00958_),
    .Q(\cpuregs[15][7] ));
 sky130_fd_sc_hd__dfxtp_4 _49041_ (.CLK(clk_0_160),
    .D(_00959_),
    .Q(\cpuregs[15][8] ));
 sky130_fd_sc_hd__dfxtp_4 _49042_ (.CLK(clk_0_160),
    .D(_00960_),
    .Q(\cpuregs[15][9] ));
 sky130_fd_sc_hd__dfxtp_4 _49043_ (.CLK(clk_0_160),
    .D(_00930_),
    .Q(\cpuregs[15][10] ));
 sky130_fd_sc_hd__dfxtp_4 _49044_ (.CLK(clk_0_160),
    .D(_00931_),
    .Q(\cpuregs[15][11] ));
 sky130_fd_sc_hd__dfxtp_4 _49045_ (.CLK(clk_0_160),
    .D(_00932_),
    .Q(\cpuregs[15][12] ));
 sky130_fd_sc_hd__dfxtp_4 _49046_ (.CLK(clk_0_176),
    .D(_00933_),
    .Q(\cpuregs[15][13] ));
 sky130_fd_sc_hd__dfxtp_4 _49047_ (.CLK(clk_0_176),
    .D(_00934_),
    .Q(\cpuregs[15][14] ));
 sky130_fd_sc_hd__dfxtp_4 _49048_ (.CLK(clk_0_176),
    .D(_00935_),
    .Q(\cpuregs[15][15] ));
 sky130_fd_sc_hd__dfxtp_4 _49049_ (.CLK(clk_0_176),
    .D(_00936_),
    .Q(\cpuregs[15][16] ));
 sky130_fd_sc_hd__dfxtp_4 _49050_ (.CLK(clk_0_176),
    .D(_00937_),
    .Q(\cpuregs[15][17] ));
 sky130_fd_sc_hd__dfxtp_4 _49051_ (.CLK(clk_0_176),
    .D(_00938_),
    .Q(\cpuregs[15][18] ));
 sky130_fd_sc_hd__dfxtp_4 _49052_ (.CLK(clk_0_176),
    .D(_00939_),
    .Q(\cpuregs[15][19] ));
 sky130_fd_sc_hd__dfxtp_4 _49053_ (.CLK(clk_0_176),
    .D(_00941_),
    .Q(\cpuregs[15][20] ));
 sky130_fd_sc_hd__dfxtp_4 _49054_ (.CLK(clk_0_176),
    .D(_00942_),
    .Q(\cpuregs[15][21] ));
 sky130_fd_sc_hd__dfxtp_4 _49055_ (.CLK(clk_0_176),
    .D(_00943_),
    .Q(\cpuregs[15][22] ));
 sky130_fd_sc_hd__dfxtp_4 _49056_ (.CLK(clk_0_176),
    .D(_00944_),
    .Q(\cpuregs[15][23] ));
 sky130_fd_sc_hd__dfxtp_4 _49057_ (.CLK(clk_0_176),
    .D(_00945_),
    .Q(\cpuregs[15][24] ));
 sky130_fd_sc_hd__dfxtp_4 _49058_ (.CLK(clk_0_176),
    .D(_00946_),
    .Q(\cpuregs[15][25] ));
 sky130_fd_sc_hd__dfxtp_4 _49059_ (.CLK(clk_0_176),
    .D(_00947_),
    .Q(\cpuregs[15][26] ));
 sky130_fd_sc_hd__dfxtp_4 _49060_ (.CLK(clk_0_176),
    .D(_00948_),
    .Q(\cpuregs[15][27] ));
 sky130_fd_sc_hd__dfxtp_4 _49061_ (.CLK(clk_0_176),
    .D(_00949_),
    .Q(\cpuregs[15][28] ));
 sky130_fd_sc_hd__dfxtp_4 _49062_ (.CLK(clk_0_192),
    .D(_00950_),
    .Q(\cpuregs[15][29] ));
 sky130_fd_sc_hd__dfxtp_4 _49063_ (.CLK(clk_0_192),
    .D(_00952_),
    .Q(\cpuregs[15][30] ));
 sky130_fd_sc_hd__dfxtp_4 _49064_ (.CLK(clk_0_192),
    .D(_00953_),
    .Q(\cpuregs[15][31] ));
 sky130_fd_sc_hd__dfxtp_4 _49065_ (.CLK(clk_0_192),
    .D(_01057_),
    .Q(\cpuregs[19][0] ));
 sky130_fd_sc_hd__dfxtp_4 _49066_ (.CLK(clk_0_192),
    .D(_01068_),
    .Q(\cpuregs[19][1] ));
 sky130_fd_sc_hd__dfxtp_4 _49067_ (.CLK(clk_0_192),
    .D(_01079_),
    .Q(\cpuregs[19][2] ));
 sky130_fd_sc_hd__dfxtp_4 _49068_ (.CLK(clk_0_192),
    .D(_01082_),
    .Q(\cpuregs[19][3] ));
 sky130_fd_sc_hd__dfxtp_4 _49069_ (.CLK(clk_0_192),
    .D(_01083_),
    .Q(\cpuregs[19][4] ));
 sky130_fd_sc_hd__dfxtp_4 _49070_ (.CLK(clk_0_192),
    .D(_01084_),
    .Q(\cpuregs[19][5] ));
 sky130_fd_sc_hd__dfxtp_4 _49071_ (.CLK(clk_0_192),
    .D(_01085_),
    .Q(\cpuregs[19][6] ));
 sky130_fd_sc_hd__dfxtp_4 _49072_ (.CLK(clk_0_192),
    .D(_01086_),
    .Q(\cpuregs[19][7] ));
 sky130_fd_sc_hd__dfxtp_4 _49073_ (.CLK(clk_0_192),
    .D(_01087_),
    .Q(\cpuregs[19][8] ));
 sky130_fd_sc_hd__dfxtp_4 _49074_ (.CLK(clk_0_192),
    .D(_01088_),
    .Q(\cpuregs[19][9] ));
 sky130_fd_sc_hd__dfxtp_4 _49075_ (.CLK(clk_0_192),
    .D(_01058_),
    .Q(\cpuregs[19][10] ));
 sky130_fd_sc_hd__dfxtp_4 _49076_ (.CLK(clk_0_192),
    .D(_01059_),
    .Q(\cpuregs[19][11] ));
 sky130_fd_sc_hd__dfxtp_4 _49077_ (.CLK(clk_0_192),
    .D(_01060_),
    .Q(\cpuregs[19][12] ));
 sky130_fd_sc_hd__dfxtp_4 _49078_ (.CLK(clk_0_208),
    .D(_01061_),
    .Q(\cpuregs[19][13] ));
 sky130_fd_sc_hd__dfxtp_4 _49079_ (.CLK(clk_0_208),
    .D(_01062_),
    .Q(\cpuregs[19][14] ));
 sky130_fd_sc_hd__dfxtp_4 _49080_ (.CLK(clk_0_208),
    .D(_01063_),
    .Q(\cpuregs[19][15] ));
 sky130_fd_sc_hd__dfxtp_4 _49081_ (.CLK(clk_0_208),
    .D(_01064_),
    .Q(\cpuregs[19][16] ));
 sky130_fd_sc_hd__dfxtp_4 _49082_ (.CLK(clk_0_208),
    .D(_01065_),
    .Q(\cpuregs[19][17] ));
 sky130_fd_sc_hd__dfxtp_4 _49083_ (.CLK(clk_0_208),
    .D(_01066_),
    .Q(\cpuregs[19][18] ));
 sky130_fd_sc_hd__dfxtp_4 _49084_ (.CLK(clk_0_208),
    .D(_01067_),
    .Q(\cpuregs[19][19] ));
 sky130_fd_sc_hd__dfxtp_4 _49085_ (.CLK(clk_0_208),
    .D(_01069_),
    .Q(\cpuregs[19][20] ));
 sky130_fd_sc_hd__dfxtp_4 _49086_ (.CLK(clk_0_208),
    .D(_01070_),
    .Q(\cpuregs[19][21] ));
 sky130_fd_sc_hd__dfxtp_4 _49087_ (.CLK(clk_0_208),
    .D(_01071_),
    .Q(\cpuregs[19][22] ));
 sky130_fd_sc_hd__dfxtp_4 _49088_ (.CLK(clk_0_208),
    .D(_01072_),
    .Q(\cpuregs[19][23] ));
 sky130_fd_sc_hd__dfxtp_4 _49089_ (.CLK(clk_0_208),
    .D(_01073_),
    .Q(\cpuregs[19][24] ));
 sky130_fd_sc_hd__dfxtp_4 _49090_ (.CLK(clk_0_208),
    .D(_01074_),
    .Q(\cpuregs[19][25] ));
 sky130_fd_sc_hd__dfxtp_4 _49091_ (.CLK(clk_0_208),
    .D(_01075_),
    .Q(\cpuregs[19][26] ));
 sky130_fd_sc_hd__dfxtp_4 _49092_ (.CLK(clk_0_208),
    .D(_01076_),
    .Q(\cpuregs[19][27] ));
 sky130_fd_sc_hd__dfxtp_4 _49093_ (.CLK(clk_0_208),
    .D(_01077_),
    .Q(\cpuregs[19][28] ));
 sky130_fd_sc_hd__dfxtp_4 _49094_ (.CLK(clk_0_224),
    .D(_01078_),
    .Q(\cpuregs[19][29] ));
 sky130_fd_sc_hd__dfxtp_4 _49095_ (.CLK(clk_0_224),
    .D(_01080_),
    .Q(\cpuregs[19][30] ));
 sky130_fd_sc_hd__dfxtp_4 _49096_ (.CLK(clk_0_224),
    .D(_01081_),
    .Q(\cpuregs[19][31] ));
 sky130_fd_sc_hd__dfxtp_4 _49097_ (.CLK(clk_0_224),
    .D(_00658_),
    .Q(trap));
 sky130_fd_sc_hd__dfxtp_4 _49098_ (.CLK(clk_0_224),
    .D(_00497_),
    .Q(pcpi_valid));
 sky130_fd_sc_hd__dfxtp_4 _49099_ (.CLK(clk_0_224),
    .D(_00214_),
    .Q(eoi[0]));
 sky130_fd_sc_hd__dfxtp_4 _49100_ (.CLK(clk_0_224),
    .D(_00225_),
    .Q(eoi[1]));
 sky130_fd_sc_hd__dfxtp_4 _49101_ (.CLK(clk_0_224),
    .D(_00236_),
    .Q(eoi[2]));
 sky130_fd_sc_hd__dfxtp_4 _49102_ (.CLK(clk_0_224),
    .D(_00239_),
    .Q(eoi[3]));
 sky130_fd_sc_hd__dfxtp_4 _49103_ (.CLK(clk_0_224),
    .D(_00240_),
    .Q(eoi[4]));
 sky130_fd_sc_hd__dfxtp_4 _49104_ (.CLK(clk_0_224),
    .D(_00241_),
    .Q(eoi[5]));
 sky130_fd_sc_hd__dfxtp_4 _49105_ (.CLK(clk_0_224),
    .D(_00242_),
    .Q(eoi[6]));
 sky130_fd_sc_hd__dfxtp_4 _49106_ (.CLK(clk_0_224),
    .D(_00243_),
    .Q(eoi[7]));
 sky130_fd_sc_hd__dfxtp_4 _49107_ (.CLK(clk_0_224),
    .D(_00244_),
    .Q(eoi[8]));
 sky130_fd_sc_hd__dfxtp_4 _49108_ (.CLK(clk_0_224),
    .D(_00245_),
    .Q(eoi[9]));
 sky130_fd_sc_hd__dfxtp_4 _49109_ (.CLK(clk_0_224),
    .D(_00215_),
    .Q(eoi[10]));
 sky130_fd_sc_hd__dfxtp_4 _49110_ (.CLK(clk_0_240),
    .D(_00216_),
    .Q(eoi[11]));
 sky130_fd_sc_hd__dfxtp_4 _49111_ (.CLK(clk_0_240),
    .D(_00217_),
    .Q(eoi[12]));
 sky130_fd_sc_hd__dfxtp_4 _49112_ (.CLK(clk_0_240),
    .D(_00218_),
    .Q(eoi[13]));
 sky130_fd_sc_hd__dfxtp_4 _49113_ (.CLK(clk_0_240),
    .D(_00219_),
    .Q(eoi[14]));
 sky130_fd_sc_hd__dfxtp_4 _49114_ (.CLK(clk_0_240),
    .D(_00220_),
    .Q(eoi[15]));
 sky130_fd_sc_hd__dfxtp_4 _49115_ (.CLK(clk_0_240),
    .D(_00221_),
    .Q(eoi[16]));
 sky130_fd_sc_hd__dfxtp_4 _49116_ (.CLK(clk_0_240),
    .D(_00222_),
    .Q(eoi[17]));
 sky130_fd_sc_hd__dfxtp_4 _49117_ (.CLK(clk_0_240),
    .D(_00223_),
    .Q(eoi[18]));
 sky130_fd_sc_hd__dfxtp_4 _49118_ (.CLK(clk_0_240),
    .D(_00224_),
    .Q(eoi[19]));
 sky130_fd_sc_hd__dfxtp_4 _49119_ (.CLK(clk_0_240),
    .D(_00226_),
    .Q(eoi[20]));
 sky130_fd_sc_hd__dfxtp_4 _49120_ (.CLK(clk_0_240),
    .D(_00227_),
    .Q(eoi[21]));
 sky130_fd_sc_hd__dfxtp_4 _49121_ (.CLK(clk_0_240),
    .D(_00228_),
    .Q(eoi[22]));
 sky130_fd_sc_hd__dfxtp_4 _49122_ (.CLK(clk_0_240),
    .D(_00229_),
    .Q(eoi[23]));
 sky130_fd_sc_hd__dfxtp_4 _49123_ (.CLK(clk_0_240),
    .D(_00230_),
    .Q(eoi[24]));
 sky130_fd_sc_hd__dfxtp_4 _49124_ (.CLK(clk_0_240),
    .D(_00231_),
    .Q(eoi[25]));
 sky130_fd_sc_hd__dfxtp_4 _49125_ (.CLK(clk_0_240),
    .D(_00232_),
    .Q(eoi[26]));
 sky130_fd_sc_hd__dfxtp_4 _49126_ (.CLK(clk_0_256),
    .D(_00233_),
    .Q(eoi[27]));
 sky130_fd_sc_hd__dfxtp_4 _49127_ (.CLK(clk_0_256),
    .D(_00234_),
    .Q(eoi[28]));
 sky130_fd_sc_hd__dfxtp_4 _49128_ (.CLK(clk_0_256),
    .D(_00235_),
    .Q(eoi[29]));
 sky130_fd_sc_hd__dfxtp_4 _49129_ (.CLK(clk_0_256),
    .D(_00237_),
    .Q(eoi[30]));
 sky130_fd_sc_hd__dfxtp_4 _49130_ (.CLK(clk_0_256),
    .D(_00238_),
    .Q(eoi[31]));
 sky130_fd_sc_hd__dfxtp_4 _49131_ (.CLK(clk_0_256),
    .D(_00004_),
    .Q(\count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49132_ (.CLK(clk_0_256),
    .D(_00015_),
    .Q(\count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49133_ (.CLK(clk_0_256),
    .D(_00026_),
    .Q(\count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49134_ (.CLK(clk_0_256),
    .D(_00037_),
    .Q(\count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49135_ (.CLK(clk_0_256),
    .D(_00048_),
    .Q(\count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49136_ (.CLK(clk_0_256),
    .D(_00059_),
    .Q(\count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49137_ (.CLK(clk_0_256),
    .D(_00064_),
    .Q(\count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49138_ (.CLK(clk_0_256),
    .D(_00065_),
    .Q(\count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49139_ (.CLK(clk_0_256),
    .D(_00066_),
    .Q(\count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49140_ (.CLK(clk_0_256),
    .D(_00067_),
    .Q(\count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49141_ (.CLK(clk_0_256),
    .D(_00005_),
    .Q(\count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49142_ (.CLK(clk_0_272),
    .D(_00006_),
    .Q(\count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49143_ (.CLK(clk_0_272),
    .D(_00007_),
    .Q(\count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49144_ (.CLK(clk_0_272),
    .D(_00008_),
    .Q(\count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49145_ (.CLK(clk_0_272),
    .D(_00009_),
    .Q(\count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49146_ (.CLK(clk_0_272),
    .D(_00010_),
    .Q(\count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49147_ (.CLK(clk_0_272),
    .D(_00011_),
    .Q(\count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49148_ (.CLK(clk_0_272),
    .D(_00012_),
    .Q(\count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49149_ (.CLK(clk_0_272),
    .D(_00013_),
    .Q(\count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49150_ (.CLK(clk_0_272),
    .D(_00014_),
    .Q(\count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49151_ (.CLK(clk_0_272),
    .D(_00016_),
    .Q(\count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49152_ (.CLK(clk_0_272),
    .D(_00017_),
    .Q(\count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49153_ (.CLK(clk_0_272),
    .D(_00018_),
    .Q(\count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49154_ (.CLK(clk_0_272),
    .D(_00019_),
    .Q(\count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49155_ (.CLK(clk_0_272),
    .D(_00020_),
    .Q(\count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49156_ (.CLK(clk_0_272),
    .D(_00021_),
    .Q(\count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49157_ (.CLK(clk_0_272),
    .D(_00022_),
    .Q(\count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49158_ (.CLK(clk_0_288),
    .D(_00023_),
    .Q(\count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49159_ (.CLK(clk_0_288),
    .D(_00024_),
    .Q(\count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49160_ (.CLK(clk_0_288),
    .D(_00025_),
    .Q(\count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49161_ (.CLK(clk_0_288),
    .D(_00027_),
    .Q(\count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49162_ (.CLK(clk_0_288),
    .D(_00028_),
    .Q(\count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49163_ (.CLK(clk_0_288),
    .D(_00029_),
    .Q(\count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_4 _49164_ (.CLK(clk_0_288),
    .D(_00030_),
    .Q(\count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_4 _49165_ (.CLK(clk_0_288),
    .D(_00031_),
    .Q(\count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_4 _49166_ (.CLK(clk_0_288),
    .D(_00032_),
    .Q(\count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_4 _49167_ (.CLK(clk_0_288),
    .D(_00033_),
    .Q(\count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_4 _49168_ (.CLK(clk_0_288),
    .D(_00034_),
    .Q(\count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_4 _49169_ (.CLK(clk_0_288),
    .D(_00035_),
    .Q(\count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_4 _49170_ (.CLK(clk_0_288),
    .D(_00036_),
    .Q(\count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_4 _49171_ (.CLK(clk_0_288),
    .D(_00038_),
    .Q(\count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_4 _49172_ (.CLK(clk_0_288),
    .D(_00039_),
    .Q(\count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_4 _49173_ (.CLK(clk_0_288),
    .D(_00040_),
    .Q(\count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_4 _49174_ (.CLK(clk_0_304),
    .D(_00041_),
    .Q(\count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_4 _49175_ (.CLK(clk_0_304),
    .D(_00042_),
    .Q(\count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_4 _49176_ (.CLK(clk_0_304),
    .D(_00043_),
    .Q(\count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_4 _49177_ (.CLK(clk_0_304),
    .D(_00044_),
    .Q(\count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_4 _49178_ (.CLK(clk_0_304),
    .D(_00045_),
    .Q(\count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_4 _49179_ (.CLK(clk_0_304),
    .D(_00046_),
    .Q(\count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_4 _49180_ (.CLK(clk_0_304),
    .D(_00047_),
    .Q(\count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_4 _49181_ (.CLK(clk_0_304),
    .D(_00049_),
    .Q(\count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_4 _49182_ (.CLK(clk_0_304),
    .D(_00050_),
    .Q(\count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_4 _49183_ (.CLK(clk_0_304),
    .D(_00051_),
    .Q(\count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_4 _49184_ (.CLK(clk_0_304),
    .D(_00052_),
    .Q(\count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_4 _49185_ (.CLK(clk_0_304),
    .D(_00053_),
    .Q(\count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_4 _49186_ (.CLK(clk_0_304),
    .D(_00054_),
    .Q(\count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_4 _49187_ (.CLK(clk_0_304),
    .D(_00055_),
    .Q(\count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_4 _49188_ (.CLK(clk_0_304),
    .D(_00056_),
    .Q(\count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_4 _49189_ (.CLK(clk_0_304),
    .D(_00057_),
    .Q(\count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_4 _49190_ (.CLK(clk_0_320),
    .D(_00058_),
    .Q(\count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_4 _49191_ (.CLK(clk_0_320),
    .D(_00060_),
    .Q(\count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_4 _49192_ (.CLK(clk_0_320),
    .D(_00061_),
    .Q(\count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_4 _49193_ (.CLK(clk_0_320),
    .D(_00062_),
    .Q(\count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_4 _49194_ (.CLK(clk_0_320),
    .D(_00063_),
    .Q(\count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_4 _49195_ (.CLK(clk_0_320),
    .D(_00068_),
    .Q(\count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49196_ (.CLK(clk_0_320),
    .D(_00079_),
    .Q(\count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49197_ (.CLK(clk_0_320),
    .D(_00090_),
    .Q(\count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49198_ (.CLK(clk_0_320),
    .D(_00101_),
    .Q(\count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49199_ (.CLK(clk_0_320),
    .D(_00112_),
    .Q(\count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49200_ (.CLK(clk_0_320),
    .D(_00123_),
    .Q(\count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49201_ (.CLK(clk_0_320),
    .D(_00128_),
    .Q(\count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49202_ (.CLK(clk_0_320),
    .D(_00129_),
    .Q(\count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49203_ (.CLK(clk_0_320),
    .D(_00130_),
    .Q(\count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49204_ (.CLK(clk_0_320),
    .D(_00131_),
    .Q(\count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49205_ (.CLK(clk_0_320),
    .D(_00069_),
    .Q(\count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49206_ (.CLK(clk_0_336),
    .D(_00070_),
    .Q(\count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49207_ (.CLK(clk_0_336),
    .D(_00071_),
    .Q(\count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49208_ (.CLK(clk_0_336),
    .D(_00072_),
    .Q(\count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49209_ (.CLK(clk_0_336),
    .D(_00073_),
    .Q(\count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49210_ (.CLK(clk_0_336),
    .D(_00074_),
    .Q(\count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49211_ (.CLK(clk_0_336),
    .D(_00075_),
    .Q(\count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49212_ (.CLK(clk_0_336),
    .D(_00076_),
    .Q(\count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49213_ (.CLK(clk_0_336),
    .D(_00077_),
    .Q(\count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49214_ (.CLK(clk_0_336),
    .D(_00078_),
    .Q(\count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49215_ (.CLK(clk_0_336),
    .D(_00080_),
    .Q(\count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49216_ (.CLK(clk_0_336),
    .D(_00081_),
    .Q(\count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49217_ (.CLK(clk_0_336),
    .D(_00082_),
    .Q(\count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49218_ (.CLK(clk_0_336),
    .D(_00083_),
    .Q(\count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49219_ (.CLK(clk_0_336),
    .D(_00084_),
    .Q(\count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49220_ (.CLK(clk_0_336),
    .D(_00085_),
    .Q(\count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49221_ (.CLK(clk_0_336),
    .D(_00086_),
    .Q(\count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49222_ (.CLK(clk_0_352),
    .D(_00087_),
    .Q(\count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49223_ (.CLK(clk_0_352),
    .D(_00088_),
    .Q(\count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49224_ (.CLK(clk_0_352),
    .D(_00089_),
    .Q(\count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49225_ (.CLK(clk_0_352),
    .D(_00091_),
    .Q(\count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49226_ (.CLK(clk_0_352),
    .D(_00092_),
    .Q(\count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49227_ (.CLK(clk_0_352),
    .D(_00093_),
    .Q(\count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_4 _49228_ (.CLK(clk_0_352),
    .D(_00094_),
    .Q(\count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_4 _49229_ (.CLK(clk_0_352),
    .D(_00095_),
    .Q(\count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_4 _49230_ (.CLK(clk_0_352),
    .D(_00096_),
    .Q(\count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_4 _49231_ (.CLK(clk_0_352),
    .D(_00097_),
    .Q(\count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_4 _49232_ (.CLK(clk_0_352),
    .D(_00098_),
    .Q(\count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_4 _49233_ (.CLK(clk_0_352),
    .D(_00099_),
    .Q(\count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_4 _49234_ (.CLK(clk_0_352),
    .D(_00100_),
    .Q(\count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_4 _49235_ (.CLK(clk_0_352),
    .D(_00102_),
    .Q(\count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_4 _49236_ (.CLK(clk_0_352),
    .D(_00103_),
    .Q(\count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_4 _49237_ (.CLK(clk_0_352),
    .D(_00104_),
    .Q(\count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_4 _49238_ (.CLK(clk_0_368),
    .D(_00105_),
    .Q(\count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_4 _49239_ (.CLK(clk_0_368),
    .D(_00106_),
    .Q(\count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_4 _49240_ (.CLK(clk_0_368),
    .D(_00107_),
    .Q(\count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_4 _49241_ (.CLK(clk_0_368),
    .D(_00108_),
    .Q(\count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_4 _49242_ (.CLK(clk_0_368),
    .D(_00109_),
    .Q(\count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_4 _49243_ (.CLK(clk_0_368),
    .D(_00110_),
    .Q(\count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_4 _49244_ (.CLK(clk_0_368),
    .D(_00111_),
    .Q(\count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_4 _49245_ (.CLK(clk_0_368),
    .D(_00113_),
    .Q(\count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_4 _49246_ (.CLK(clk_0_368),
    .D(_00114_),
    .Q(\count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_4 _49247_ (.CLK(clk_0_368),
    .D(_00115_),
    .Q(\count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_4 _49248_ (.CLK(clk_0_368),
    .D(_00116_),
    .Q(\count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_4 _49249_ (.CLK(clk_0_368),
    .D(_00117_),
    .Q(\count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_4 _49250_ (.CLK(clk_0_368),
    .D(_00118_),
    .Q(\count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_4 _49251_ (.CLK(clk_0_368),
    .D(_00119_),
    .Q(\count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_4 _49252_ (.CLK(clk_0_368),
    .D(_00120_),
    .Q(\count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_4 _49253_ (.CLK(clk_0_368),
    .D(_00121_),
    .Q(\count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_4 _49254_ (.CLK(clk_0_384),
    .D(_00122_),
    .Q(\count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_4 _49255_ (.CLK(clk_0_384),
    .D(_00124_),
    .Q(\count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_4 _49256_ (.CLK(clk_0_384),
    .D(_00125_),
    .Q(\count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_4 _49257_ (.CLK(clk_0_384),
    .D(_00126_),
    .Q(\count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_4 _49258_ (.CLK(clk_0_384),
    .D(_00127_),
    .Q(\count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_4 _49259_ (.CLK(clk_0_384),
    .D(_00594_),
    .Q(\reg_pc[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49260_ (.CLK(clk_0_384),
    .D(_00605_),
    .Q(\reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49261_ (.CLK(clk_0_384),
    .D(_00616_),
    .Q(\reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49262_ (.CLK(clk_0_384),
    .D(_00619_),
    .Q(\reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49263_ (.CLK(clk_0_384),
    .D(_00620_),
    .Q(\reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49264_ (.CLK(clk_0_384),
    .D(_00621_),
    .Q(\reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49265_ (.CLK(clk_0_384),
    .D(_00622_),
    .Q(\reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49266_ (.CLK(clk_0_384),
    .D(_00623_),
    .Q(\reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49267_ (.CLK(clk_0_384),
    .D(_00624_),
    .Q(\reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49268_ (.CLK(clk_0_384),
    .D(_00625_),
    .Q(\reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49269_ (.CLK(clk_0_384),
    .D(_00595_),
    .Q(\reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49270_ (.CLK(clk_0_400),
    .D(_00596_),
    .Q(\reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49271_ (.CLK(clk_0_400),
    .D(_00597_),
    .Q(\reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49272_ (.CLK(clk_0_400),
    .D(_00598_),
    .Q(\reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49273_ (.CLK(clk_0_400),
    .D(_00599_),
    .Q(\reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49274_ (.CLK(clk_0_400),
    .D(_00600_),
    .Q(\reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49275_ (.CLK(clk_0_400),
    .D(_00601_),
    .Q(\reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49276_ (.CLK(clk_0_400),
    .D(_00602_),
    .Q(\reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49277_ (.CLK(clk_0_400),
    .D(_00603_),
    .Q(\reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49278_ (.CLK(clk_0_400),
    .D(_00604_),
    .Q(\reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49279_ (.CLK(clk_0_400),
    .D(_00606_),
    .Q(\reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49280_ (.CLK(clk_0_400),
    .D(_00607_),
    .Q(\reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49281_ (.CLK(clk_0_400),
    .D(_00608_),
    .Q(\reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49282_ (.CLK(clk_0_400),
    .D(_00609_),
    .Q(\reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49283_ (.CLK(clk_0_400),
    .D(_00610_),
    .Q(\reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49284_ (.CLK(clk_0_400),
    .D(_00611_),
    .Q(\reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49285_ (.CLK(clk_0_400),
    .D(_00612_),
    .Q(\reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49286_ (.CLK(clk_0_416),
    .D(_00613_),
    .Q(\reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49287_ (.CLK(clk_0_416),
    .D(_00614_),
    .Q(\reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49288_ (.CLK(clk_0_416),
    .D(_00615_),
    .Q(\reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49289_ (.CLK(clk_0_416),
    .D(_00617_),
    .Q(\reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49290_ (.CLK(clk_0_416),
    .D(_00618_),
    .Q(\reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49291_ (.CLK(clk_0_416),
    .D(_00498_),
    .Q(\reg_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49292_ (.CLK(clk_0_416),
    .D(_00509_),
    .Q(\reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49293_ (.CLK(clk_0_416),
    .D(_00520_),
    .Q(\reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49294_ (.CLK(clk_0_416),
    .D(_00523_),
    .Q(\reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49295_ (.CLK(clk_0_416),
    .D(_00524_),
    .Q(\reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49296_ (.CLK(clk_0_416),
    .D(_00525_),
    .Q(\reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49297_ (.CLK(clk_0_416),
    .D(_00526_),
    .Q(\reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49298_ (.CLK(clk_0_416),
    .D(_00527_),
    .Q(\reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49299_ (.CLK(clk_0_416),
    .D(_00528_),
    .Q(\reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49300_ (.CLK(clk_0_416),
    .D(_00529_),
    .Q(\reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49301_ (.CLK(clk_0_416),
    .D(_00499_),
    .Q(\reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49302_ (.CLK(clk_0_432),
    .D(_00500_),
    .Q(\reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49303_ (.CLK(clk_0_432),
    .D(_00501_),
    .Q(\reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49304_ (.CLK(clk_0_432),
    .D(_00502_),
    .Q(\reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49305_ (.CLK(clk_0_432),
    .D(_00503_),
    .Q(\reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49306_ (.CLK(clk_0_432),
    .D(_00504_),
    .Q(\reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49307_ (.CLK(clk_0_432),
    .D(_00505_),
    .Q(\reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49308_ (.CLK(clk_0_432),
    .D(_00506_),
    .Q(\reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49309_ (.CLK(clk_0_432),
    .D(_00507_),
    .Q(\reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49310_ (.CLK(clk_0_432),
    .D(_00508_),
    .Q(\reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49311_ (.CLK(clk_0_432),
    .D(_00510_),
    .Q(\reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49312_ (.CLK(clk_0_432),
    .D(_00511_),
    .Q(\reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49313_ (.CLK(clk_0_432),
    .D(_00512_),
    .Q(\reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49314_ (.CLK(clk_0_432),
    .D(_00513_),
    .Q(\reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49315_ (.CLK(clk_0_432),
    .D(_00514_),
    .Q(\reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49316_ (.CLK(clk_0_432),
    .D(_00515_),
    .Q(\reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49317_ (.CLK(clk_0_432),
    .D(_00516_),
    .Q(\reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49318_ (.CLK(clk_0_448),
    .D(_00517_),
    .Q(\reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49319_ (.CLK(clk_0_448),
    .D(_00518_),
    .Q(\reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49320_ (.CLK(clk_0_448),
    .D(_00519_),
    .Q(\reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49321_ (.CLK(clk_0_448),
    .D(_00521_),
    .Q(\reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49322_ (.CLK(clk_0_448),
    .D(_00522_),
    .Q(\reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49323_ (.CLK(clk_0_448),
    .D(_00530_),
    .Q(pcpi_rs1[0]));
 sky130_fd_sc_hd__dfxtp_4 _49324_ (.CLK(clk_0_448),
    .D(_00541_),
    .Q(pcpi_rs1[1]));
 sky130_fd_sc_hd__dfxtp_4 _49325_ (.CLK(clk_0_448),
    .D(_00552_),
    .Q(pcpi_rs1[2]));
 sky130_fd_sc_hd__dfxtp_4 _49326_ (.CLK(clk_0_448),
    .D(_00555_),
    .Q(pcpi_rs1[3]));
 sky130_fd_sc_hd__dfxtp_4 _49327_ (.CLK(clk_0_448),
    .D(_00556_),
    .Q(pcpi_rs1[4]));
 sky130_fd_sc_hd__dfxtp_4 _49328_ (.CLK(clk_0_448),
    .D(_00557_),
    .Q(pcpi_rs1[5]));
 sky130_fd_sc_hd__dfxtp_4 _49329_ (.CLK(clk_0_448),
    .D(_00558_),
    .Q(pcpi_rs1[6]));
 sky130_fd_sc_hd__dfxtp_4 _49330_ (.CLK(clk_0_448),
    .D(_00559_),
    .Q(pcpi_rs1[7]));
 sky130_fd_sc_hd__dfxtp_4 _49331_ (.CLK(clk_0_448),
    .D(_00560_),
    .Q(pcpi_rs1[8]));
 sky130_fd_sc_hd__dfxtp_4 _49332_ (.CLK(clk_0_448),
    .D(_00561_),
    .Q(pcpi_rs1[9]));
 sky130_fd_sc_hd__dfxtp_4 _49333_ (.CLK(clk_0_448),
    .D(_00531_),
    .Q(pcpi_rs1[10]));
 sky130_fd_sc_hd__dfxtp_4 _49334_ (.CLK(clk_0_464),
    .D(_00532_),
    .Q(pcpi_rs1[11]));
 sky130_fd_sc_hd__dfxtp_4 _49335_ (.CLK(clk_0_464),
    .D(_00533_),
    .Q(pcpi_rs1[12]));
 sky130_fd_sc_hd__dfxtp_4 _49336_ (.CLK(clk_0_464),
    .D(_00534_),
    .Q(pcpi_rs1[13]));
 sky130_fd_sc_hd__dfxtp_4 _49337_ (.CLK(clk_0_464),
    .D(_00535_),
    .Q(pcpi_rs1[14]));
 sky130_fd_sc_hd__dfxtp_4 _49338_ (.CLK(clk_0_464),
    .D(_00536_),
    .Q(pcpi_rs1[15]));
 sky130_fd_sc_hd__dfxtp_4 _49339_ (.CLK(clk_0_464),
    .D(_00537_),
    .Q(pcpi_rs1[16]));
 sky130_fd_sc_hd__dfxtp_4 _49340_ (.CLK(clk_0_464),
    .D(_00538_),
    .Q(pcpi_rs1[17]));
 sky130_fd_sc_hd__dfxtp_4 _49341_ (.CLK(clk_0_464),
    .D(_00539_),
    .Q(pcpi_rs1[18]));
 sky130_fd_sc_hd__dfxtp_4 _49342_ (.CLK(clk_0_464),
    .D(_00540_),
    .Q(pcpi_rs1[19]));
 sky130_fd_sc_hd__dfxtp_4 _49343_ (.CLK(clk_0_464),
    .D(_00542_),
    .Q(pcpi_rs1[20]));
 sky130_fd_sc_hd__dfxtp_4 _49344_ (.CLK(clk_0_464),
    .D(_00543_),
    .Q(pcpi_rs1[21]));
 sky130_fd_sc_hd__dfxtp_4 _49345_ (.CLK(clk_0_464),
    .D(_00544_),
    .Q(pcpi_rs1[22]));
 sky130_fd_sc_hd__dfxtp_4 _49346_ (.CLK(clk_0_464),
    .D(_00545_),
    .Q(pcpi_rs1[23]));
 sky130_fd_sc_hd__dfxtp_4 _49347_ (.CLK(clk_0_464),
    .D(_00546_),
    .Q(pcpi_rs1[24]));
 sky130_fd_sc_hd__dfxtp_4 _49348_ (.CLK(clk_0_464),
    .D(_00547_),
    .Q(pcpi_rs1[25]));
 sky130_fd_sc_hd__dfxtp_4 _49349_ (.CLK(clk_0_464),
    .D(_00548_),
    .Q(pcpi_rs1[26]));
 sky130_fd_sc_hd__dfxtp_4 _49350_ (.CLK(clk_0_480),
    .D(_00549_),
    .Q(pcpi_rs1[27]));
 sky130_fd_sc_hd__dfxtp_4 _49351_ (.CLK(clk_0_480),
    .D(_00550_),
    .Q(pcpi_rs1[28]));
 sky130_fd_sc_hd__dfxtp_4 _49352_ (.CLK(clk_0_480),
    .D(_00551_),
    .Q(pcpi_rs1[29]));
 sky130_fd_sc_hd__dfxtp_4 _49353_ (.CLK(clk_0_480),
    .D(_00553_),
    .Q(pcpi_rs1[30]));
 sky130_fd_sc_hd__dfxtp_4 _49354_ (.CLK(clk_0_480),
    .D(_00554_),
    .Q(pcpi_rs1[31]));
 sky130_fd_sc_hd__dfxtp_4 _49355_ (.CLK(clk_0_480),
    .D(_00562_),
    .Q(mem_la_wdata[0]));
 sky130_fd_sc_hd__dfxtp_4 _49356_ (.CLK(clk_0_480),
    .D(_00573_),
    .Q(mem_la_wdata[1]));
 sky130_fd_sc_hd__dfxtp_4 _49357_ (.CLK(clk_0_480),
    .D(_00584_),
    .Q(mem_la_wdata[2]));
 sky130_fd_sc_hd__dfxtp_4 _49358_ (.CLK(clk_0_480),
    .D(_00587_),
    .Q(mem_la_wdata[3]));
 sky130_fd_sc_hd__dfxtp_4 _49359_ (.CLK(clk_0_480),
    .D(_00588_),
    .Q(mem_la_wdata[4]));
 sky130_fd_sc_hd__dfxtp_4 _49360_ (.CLK(clk_0_480),
    .D(_00589_),
    .Q(mem_la_wdata[5]));
 sky130_fd_sc_hd__dfxtp_4 _49361_ (.CLK(clk_0_480),
    .D(_00590_),
    .Q(mem_la_wdata[6]));
 sky130_fd_sc_hd__dfxtp_4 _49362_ (.CLK(clk_0_480),
    .D(_00591_),
    .Q(mem_la_wdata[7]));
 sky130_fd_sc_hd__dfxtp_4 _49363_ (.CLK(clk_0_480),
    .D(_00592_),
    .Q(pcpi_rs2[8]));
 sky130_fd_sc_hd__dfxtp_4 _49364_ (.CLK(clk_0_480),
    .D(_00593_),
    .Q(pcpi_rs2[9]));
 sky130_fd_sc_hd__dfxtp_4 _49365_ (.CLK(clk_0_480),
    .D(_00563_),
    .Q(pcpi_rs2[10]));
 sky130_fd_sc_hd__dfxtp_4 _49366_ (.CLK(clk_0_496),
    .D(_00564_),
    .Q(pcpi_rs2[11]));
 sky130_fd_sc_hd__dfxtp_4 _49367_ (.CLK(clk_0_496),
    .D(_00565_),
    .Q(pcpi_rs2[12]));
 sky130_fd_sc_hd__dfxtp_4 _49368_ (.CLK(clk_0_496),
    .D(_00566_),
    .Q(pcpi_rs2[13]));
 sky130_fd_sc_hd__dfxtp_4 _49369_ (.CLK(clk_0_496),
    .D(_00567_),
    .Q(pcpi_rs2[14]));
 sky130_fd_sc_hd__dfxtp_4 _49370_ (.CLK(clk_0_496),
    .D(_00568_),
    .Q(pcpi_rs2[15]));
 sky130_fd_sc_hd__dfxtp_4 _49371_ (.CLK(clk_0_496),
    .D(_00569_),
    .Q(pcpi_rs2[16]));
 sky130_fd_sc_hd__dfxtp_4 _49372_ (.CLK(clk_0_496),
    .D(_00570_),
    .Q(pcpi_rs2[17]));
 sky130_fd_sc_hd__dfxtp_4 _49373_ (.CLK(clk_0_496),
    .D(_00571_),
    .Q(pcpi_rs2[18]));
 sky130_fd_sc_hd__dfxtp_4 _49374_ (.CLK(clk_0_496),
    .D(_00572_),
    .Q(pcpi_rs2[19]));
 sky130_fd_sc_hd__dfxtp_4 _49375_ (.CLK(clk_0_496),
    .D(_00574_),
    .Q(pcpi_rs2[20]));
 sky130_fd_sc_hd__dfxtp_4 _49376_ (.CLK(clk_0_496),
    .D(_00575_),
    .Q(pcpi_rs2[21]));
 sky130_fd_sc_hd__dfxtp_4 _49377_ (.CLK(clk_0_496),
    .D(_00576_),
    .Q(pcpi_rs2[22]));
 sky130_fd_sc_hd__dfxtp_4 _49378_ (.CLK(clk_0_496),
    .D(_00577_),
    .Q(pcpi_rs2[23]));
 sky130_fd_sc_hd__dfxtp_4 _49379_ (.CLK(clk_0_496),
    .D(_00578_),
    .Q(pcpi_rs2[24]));
 sky130_fd_sc_hd__dfxtp_4 _49380_ (.CLK(clk_0_496),
    .D(_00579_),
    .Q(pcpi_rs2[25]));
 sky130_fd_sc_hd__dfxtp_4 _49381_ (.CLK(clk_0_496),
    .D(_00580_),
    .Q(pcpi_rs2[26]));
 sky130_fd_sc_hd__dfxtp_4 _49382_ (.CLK(clk_0_512),
    .D(_00581_),
    .Q(pcpi_rs2[27]));
 sky130_fd_sc_hd__dfxtp_4 _49383_ (.CLK(clk_0_512),
    .D(_00582_),
    .Q(pcpi_rs2[28]));
 sky130_fd_sc_hd__dfxtp_4 _49384_ (.CLK(clk_0_512),
    .D(_00583_),
    .Q(pcpi_rs2[29]));
 sky130_fd_sc_hd__dfxtp_4 _49385_ (.CLK(clk_0_512),
    .D(_00585_),
    .Q(pcpi_rs2[30]));
 sky130_fd_sc_hd__dfxtp_4 _49386_ (.CLK(clk_0_512),
    .D(_00586_),
    .Q(pcpi_rs2[31]));
 sky130_fd_sc_hd__dfxtp_4 _49387_ (.CLK(clk_0_512),
    .D(_24253_),
    .Q(\reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49388_ (.CLK(clk_0_512),
    .D(_24264_),
    .Q(\reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49389_ (.CLK(clk_0_512),
    .D(_24275_),
    .Q(\reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49390_ (.CLK(clk_0_512),
    .D(_24278_),
    .Q(\reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49391_ (.CLK(clk_0_512),
    .D(_24279_),
    .Q(\reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49392_ (.CLK(clk_0_512),
    .D(_24280_),
    .Q(\reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49393_ (.CLK(clk_0_512),
    .D(_24281_),
    .Q(\reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49394_ (.CLK(clk_0_512),
    .D(_24282_),
    .Q(\reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49395_ (.CLK(clk_0_512),
    .D(_24283_),
    .Q(\reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49396_ (.CLK(clk_0_512),
    .D(_24284_),
    .Q(\reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49397_ (.CLK(clk_0_512),
    .D(_24254_),
    .Q(\reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49398_ (.CLK(clk_0_528),
    .D(_24255_),
    .Q(\reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49399_ (.CLK(clk_0_528),
    .D(_24256_),
    .Q(\reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49400_ (.CLK(clk_0_528),
    .D(_24257_),
    .Q(\reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49401_ (.CLK(clk_0_528),
    .D(_24258_),
    .Q(\reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49402_ (.CLK(clk_0_528),
    .D(_24259_),
    .Q(\reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49403_ (.CLK(clk_0_528),
    .D(_24260_),
    .Q(\reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49404_ (.CLK(clk_0_528),
    .D(_24261_),
    .Q(\reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49405_ (.CLK(clk_0_528),
    .D(_24262_),
    .Q(\reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49406_ (.CLK(clk_0_528),
    .D(_24263_),
    .Q(\reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49407_ (.CLK(clk_0_528),
    .D(_24265_),
    .Q(\reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49408_ (.CLK(clk_0_528),
    .D(_24266_),
    .Q(\reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49409_ (.CLK(clk_0_528),
    .D(_24267_),
    .Q(\reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49410_ (.CLK(clk_0_528),
    .D(_24268_),
    .Q(\reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49411_ (.CLK(clk_0_528),
    .D(_24269_),
    .Q(\reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49412_ (.CLK(clk_0_528),
    .D(_24270_),
    .Q(\reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49413_ (.CLK(clk_0_528),
    .D(_24271_),
    .Q(\reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49414_ (.CLK(clk_0_544),
    .D(_24272_),
    .Q(\reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49415_ (.CLK(clk_0_544),
    .D(_24273_),
    .Q(\reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49416_ (.CLK(clk_0_544),
    .D(_24274_),
    .Q(\reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49417_ (.CLK(clk_0_544),
    .D(_24276_),
    .Q(\reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49418_ (.CLK(clk_0_544),
    .D(_24277_),
    .Q(\reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49419_ (.CLK(clk_0_544),
    .D(_00295_),
    .Q(irq_delay));
 sky130_fd_sc_hd__dfxtp_4 _49420_ (.CLK(clk_0_544),
    .D(_00294_),
    .Q(irq_active));
 sky130_fd_sc_hd__dfxtp_4 _49421_ (.CLK(clk_0_544),
    .D(_00296_),
    .Q(\irq_mask[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49422_ (.CLK(clk_0_544),
    .D(_00307_),
    .Q(\irq_mask[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49423_ (.CLK(clk_0_544),
    .D(_00318_),
    .Q(\irq_mask[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49424_ (.CLK(clk_0_544),
    .D(_00321_),
    .Q(\irq_mask[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49425_ (.CLK(clk_0_544),
    .D(_00322_),
    .Q(\irq_mask[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49426_ (.CLK(clk_0_544),
    .D(_00323_),
    .Q(\irq_mask[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49427_ (.CLK(clk_0_544),
    .D(_00324_),
    .Q(\irq_mask[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49428_ (.CLK(clk_0_544),
    .D(_00325_),
    .Q(\irq_mask[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49429_ (.CLK(clk_0_544),
    .D(_00326_),
    .Q(\irq_mask[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49430_ (.CLK(clk_0_560),
    .D(_00327_),
    .Q(\irq_mask[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49431_ (.CLK(clk_0_560),
    .D(_00297_),
    .Q(\irq_mask[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49432_ (.CLK(clk_0_560),
    .D(_00298_),
    .Q(\irq_mask[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49433_ (.CLK(clk_0_560),
    .D(_00299_),
    .Q(\irq_mask[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49434_ (.CLK(clk_0_560),
    .D(_00300_),
    .Q(\irq_mask[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49435_ (.CLK(clk_0_560),
    .D(_00301_),
    .Q(\irq_mask[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49436_ (.CLK(clk_0_560),
    .D(_00302_),
    .Q(\irq_mask[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49437_ (.CLK(clk_0_560),
    .D(_00303_),
    .Q(\irq_mask[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49438_ (.CLK(clk_0_560),
    .D(_00304_),
    .Q(\irq_mask[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49439_ (.CLK(clk_0_560),
    .D(_00305_),
    .Q(\irq_mask[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49440_ (.CLK(clk_0_560),
    .D(_00306_),
    .Q(\irq_mask[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49441_ (.CLK(clk_0_560),
    .D(_00308_),
    .Q(\irq_mask[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49442_ (.CLK(clk_0_560),
    .D(_00309_),
    .Q(\irq_mask[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49443_ (.CLK(clk_0_560),
    .D(_00310_),
    .Q(\irq_mask[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49444_ (.CLK(clk_0_560),
    .D(_00311_),
    .Q(\irq_mask[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49445_ (.CLK(clk_0_560),
    .D(_00312_),
    .Q(\irq_mask[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49446_ (.CLK(clk_0_576),
    .D(_00313_),
    .Q(\irq_mask[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49447_ (.CLK(clk_0_576),
    .D(_00314_),
    .Q(\irq_mask[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49448_ (.CLK(clk_0_576),
    .D(_00315_),
    .Q(\irq_mask[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49449_ (.CLK(clk_0_576),
    .D(_00316_),
    .Q(\irq_mask[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49450_ (.CLK(clk_0_576),
    .D(_00317_),
    .Q(\irq_mask[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49451_ (.CLK(clk_0_576),
    .D(_00319_),
    .Q(\irq_mask[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49452_ (.CLK(clk_0_576),
    .D(_00320_),
    .Q(\irq_mask[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49453_ (.CLK(clk_0_576),
    .D(_00328_),
    .Q(\irq_pending[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49454_ (.CLK(clk_0_576),
    .D(_00339_),
    .Q(\irq_pending[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49455_ (.CLK(clk_0_576),
    .D(_00350_),
    .Q(\irq_pending[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49456_ (.CLK(clk_0_576),
    .D(_00353_),
    .Q(\irq_pending[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49457_ (.CLK(clk_0_576),
    .D(_00354_),
    .Q(\irq_pending[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49458_ (.CLK(clk_0_576),
    .D(_00355_),
    .Q(\irq_pending[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49459_ (.CLK(clk_0_576),
    .D(_00356_),
    .Q(\irq_pending[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49460_ (.CLK(clk_0_576),
    .D(_00357_),
    .Q(\irq_pending[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49461_ (.CLK(clk_0_576),
    .D(_00358_),
    .Q(\irq_pending[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49462_ (.CLK(clk_0_592),
    .D(_00359_),
    .Q(\irq_pending[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49463_ (.CLK(clk_0_592),
    .D(_00329_),
    .Q(\irq_pending[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49464_ (.CLK(clk_0_592),
    .D(_00330_),
    .Q(\irq_pending[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49465_ (.CLK(clk_0_592),
    .D(_00331_),
    .Q(\irq_pending[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49466_ (.CLK(clk_0_592),
    .D(_00332_),
    .Q(\irq_pending[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49467_ (.CLK(clk_0_592),
    .D(_00333_),
    .Q(\irq_pending[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49468_ (.CLK(clk_0_592),
    .D(_00334_),
    .Q(\irq_pending[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49469_ (.CLK(clk_0_592),
    .D(_00335_),
    .Q(\irq_pending[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49470_ (.CLK(clk_0_592),
    .D(_00336_),
    .Q(\irq_pending[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49471_ (.CLK(clk_0_592),
    .D(_00337_),
    .Q(\irq_pending[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49472_ (.CLK(clk_0_592),
    .D(_00338_),
    .Q(\irq_pending[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49473_ (.CLK(clk_0_592),
    .D(_00340_),
    .Q(\irq_pending[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49474_ (.CLK(clk_0_592),
    .D(_00341_),
    .Q(\irq_pending[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49475_ (.CLK(clk_0_592),
    .D(_00342_),
    .Q(\irq_pending[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49476_ (.CLK(clk_0_592),
    .D(_00343_),
    .Q(\irq_pending[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49477_ (.CLK(clk_0_592),
    .D(_00344_),
    .Q(\irq_pending[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49478_ (.CLK(clk_0_608),
    .D(_00345_),
    .Q(\irq_pending[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49479_ (.CLK(clk_0_608),
    .D(_00346_),
    .Q(\irq_pending[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49480_ (.CLK(clk_0_608),
    .D(_00347_),
    .Q(\irq_pending[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49481_ (.CLK(clk_0_608),
    .D(_00348_),
    .Q(\irq_pending[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49482_ (.CLK(clk_0_608),
    .D(_00349_),
    .Q(\irq_pending[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49483_ (.CLK(clk_0_608),
    .D(_00351_),
    .Q(\irq_pending[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49484_ (.CLK(clk_0_608),
    .D(_00352_),
    .Q(\irq_pending[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49485_ (.CLK(clk_0_608),
    .D(_00626_),
    .Q(\timer[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49486_ (.CLK(clk_0_608),
    .D(_00637_),
    .Q(\timer[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49487_ (.CLK(clk_0_608),
    .D(_00648_),
    .Q(\timer[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49488_ (.CLK(clk_0_608),
    .D(_00651_),
    .Q(\timer[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49489_ (.CLK(clk_0_608),
    .D(_00652_),
    .Q(\timer[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49490_ (.CLK(clk_0_608),
    .D(_00653_),
    .Q(\timer[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49491_ (.CLK(clk_0_608),
    .D(_00654_),
    .Q(\timer[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49492_ (.CLK(clk_0_608),
    .D(_00655_),
    .Q(\timer[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49493_ (.CLK(clk_0_608),
    .D(_00656_),
    .Q(\timer[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49494_ (.CLK(clk_0_624),
    .D(_00657_),
    .Q(\timer[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49495_ (.CLK(clk_0_624),
    .D(_00627_),
    .Q(\timer[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49496_ (.CLK(clk_0_624),
    .D(_00628_),
    .Q(\timer[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49497_ (.CLK(clk_0_624),
    .D(_00629_),
    .Q(\timer[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49498_ (.CLK(clk_0_624),
    .D(_00630_),
    .Q(\timer[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49499_ (.CLK(clk_0_624),
    .D(_00631_),
    .Q(\timer[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49500_ (.CLK(clk_0_624),
    .D(_00632_),
    .Q(\timer[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49501_ (.CLK(clk_0_624),
    .D(_00633_),
    .Q(\timer[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49502_ (.CLK(clk_0_624),
    .D(_00634_),
    .Q(\timer[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49503_ (.CLK(clk_0_624),
    .D(_00635_),
    .Q(\timer[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49504_ (.CLK(clk_0_624),
    .D(_00636_),
    .Q(\timer[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49505_ (.CLK(clk_0_624),
    .D(_00638_),
    .Q(\timer[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49506_ (.CLK(clk_0_624),
    .D(_00639_),
    .Q(\timer[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49507_ (.CLK(clk_0_624),
    .D(_00640_),
    .Q(\timer[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49508_ (.CLK(clk_0_624),
    .D(_00641_),
    .Q(\timer[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49509_ (.CLK(clk_0_624),
    .D(_00642_),
    .Q(\timer[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49510_ (.CLK(clk_0_640),
    .D(_00643_),
    .Q(\timer[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49511_ (.CLK(clk_0_640),
    .D(_00644_),
    .Q(\timer[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49512_ (.CLK(clk_0_640),
    .D(_00645_),
    .Q(\timer[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49513_ (.CLK(clk_0_640),
    .D(_00646_),
    .Q(\timer[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49514_ (.CLK(clk_0_640),
    .D(_00647_),
    .Q(\timer[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49515_ (.CLK(clk_0_640),
    .D(_00649_),
    .Q(\timer[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49516_ (.CLK(clk_0_640),
    .D(_00650_),
    .Q(\timer[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49517_ (.CLK(clk_0_640),
    .D(_00416_),
    .Q(mem_do_prefetch));
 sky130_fd_sc_hd__dfxtp_4 _49518_ (.CLK(clk_0_640),
    .D(_00418_),
    .Q(mem_do_rinst));
 sky130_fd_sc_hd__dfxtp_4 _49519_ (.CLK(clk_0_640),
    .D(_00417_),
    .Q(mem_do_rdata));
 sky130_fd_sc_hd__dfxtp_4 _49520_ (.CLK(clk_0_640),
    .D(_00419_),
    .Q(mem_do_wdata));
 sky130_fd_sc_hd__dfxtp_4 _49521_ (.CLK(clk_0_640),
    .D(_00212_),
    .Q(decoder_trigger));
 sky130_fd_sc_hd__dfxtp_4 _49522_ (.CLK(clk_0_640),
    .D(_00211_),
    .Q(decoder_pseudo_trigger));
 sky130_fd_sc_hd__dfxtp_4 _49523_ (.CLK(clk_0_640),
    .D(_00360_),
    .Q(\irq_state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49524_ (.CLK(clk_0_640),
    .D(_00361_),
    .Q(\irq_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49525_ (.CLK(clk_0_640),
    .D(_00383_),
    .Q(latched_store));
 sky130_fd_sc_hd__dfxtp_4 _49526_ (.CLK(clk_0_656),
    .D(_00382_),
    .Q(latched_stalu));
 sky130_fd_sc_hd__dfxtp_4 _49527_ (.CLK(clk_0_656),
    .D(_00373_),
    .Q(latched_branch));
 sky130_fd_sc_hd__dfxtp_4 _49528_ (.CLK(clk_0_656),
    .D(_00374_),
    .Q(latched_compr));
 sky130_fd_sc_hd__dfxtp_4 _49529_ (.CLK(clk_0_656),
    .D(_00376_),
    .Q(latched_is_lh));
 sky130_fd_sc_hd__dfxtp_4 _49530_ (.CLK(clk_0_656),
    .D(_00375_),
    .Q(latched_is_lb));
 sky130_fd_sc_hd__dfxtp_4 _49531_ (.CLK(clk_0_656),
    .D(_00377_),
    .Q(\latched_rd[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49532_ (.CLK(clk_0_656),
    .D(_00378_),
    .Q(\latched_rd[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49533_ (.CLK(clk_0_656),
    .D(_00379_),
    .Q(\latched_rd[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49534_ (.CLK(clk_0_656),
    .D(_00380_),
    .Q(\latched_rd[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49535_ (.CLK(clk_0_656),
    .D(_00381_),
    .Q(\latched_rd[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49536_ (.CLK(clk_0_656),
    .D(_00493_),
    .Q(\pcpi_timeout_counter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49537_ (.CLK(clk_0_656),
    .D(_00494_),
    .Q(\pcpi_timeout_counter[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49538_ (.CLK(clk_0_656),
    .D(_00495_),
    .Q(\pcpi_timeout_counter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49539_ (.CLK(clk_0_656),
    .D(_00496_),
    .Q(\pcpi_timeout_counter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49540_ (.CLK(clk_0_656),
    .D(_00492_),
    .Q(pcpi_timeout));
 sky130_fd_sc_hd__dfxtp_4 _49541_ (.CLK(clk_0_656),
    .D(_00213_),
    .Q(do_waitirq));
 sky130_fd_sc_hd__dfxtp_4 _49542_ (.CLK(clk_0_672),
    .D(\alu_out[0] ),
    .Q(\alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49543_ (.CLK(clk_0_672),
    .D(\alu_out[1] ),
    .Q(\alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49544_ (.CLK(clk_0_672),
    .D(\alu_out[2] ),
    .Q(\alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49545_ (.CLK(clk_0_672),
    .D(\alu_out[3] ),
    .Q(\alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49546_ (.CLK(clk_0_672),
    .D(\alu_out[4] ),
    .Q(\alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49547_ (.CLK(clk_0_672),
    .D(\alu_out[5] ),
    .Q(\alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49548_ (.CLK(clk_0_672),
    .D(\alu_out[6] ),
    .Q(\alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49549_ (.CLK(clk_0_672),
    .D(\alu_out[7] ),
    .Q(\alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49550_ (.CLK(clk_0_672),
    .D(\alu_out[8] ),
    .Q(\alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49551_ (.CLK(clk_0_672),
    .D(\alu_out[9] ),
    .Q(\alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49552_ (.CLK(clk_0_672),
    .D(\alu_out[10] ),
    .Q(\alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49553_ (.CLK(clk_0_672),
    .D(\alu_out[11] ),
    .Q(\alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49554_ (.CLK(clk_0_672),
    .D(\alu_out[12] ),
    .Q(\alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49555_ (.CLK(clk_0_672),
    .D(\alu_out[13] ),
    .Q(\alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49556_ (.CLK(clk_0_672),
    .D(\alu_out[14] ),
    .Q(\alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49557_ (.CLK(clk_0_672),
    .D(\alu_out[15] ),
    .Q(\alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49558_ (.CLK(clk_0_688),
    .D(\alu_out[16] ),
    .Q(\alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49559_ (.CLK(clk_0_688),
    .D(\alu_out[17] ),
    .Q(\alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49560_ (.CLK(clk_0_688),
    .D(\alu_out[18] ),
    .Q(\alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49561_ (.CLK(clk_0_688),
    .D(\alu_out[19] ),
    .Q(\alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49562_ (.CLK(clk_0_688),
    .D(\alu_out[20] ),
    .Q(\alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49563_ (.CLK(clk_0_688),
    .D(\alu_out[21] ),
    .Q(\alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49564_ (.CLK(clk_0_688),
    .D(\alu_out[22] ),
    .Q(\alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49565_ (.CLK(clk_0_688),
    .D(\alu_out[23] ),
    .Q(\alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49566_ (.CLK(clk_0_688),
    .D(\alu_out[24] ),
    .Q(\alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49567_ (.CLK(clk_0_688),
    .D(\alu_out[25] ),
    .Q(\alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49568_ (.CLK(clk_0_688),
    .D(\alu_out[26] ),
    .Q(\alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49569_ (.CLK(clk_0_688),
    .D(\alu_out[27] ),
    .Q(\alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49570_ (.CLK(clk_0_688),
    .D(\alu_out[28] ),
    .Q(\alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49571_ (.CLK(clk_0_688),
    .D(\alu_out[29] ),
    .Q(\alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49572_ (.CLK(clk_0_688),
    .D(\alu_out[30] ),
    .Q(\alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49573_ (.CLK(clk_0_688),
    .D(\alu_out[31] ),
    .Q(\alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49574_ (.CLK(clk_0_704),
    .D(_00003_),
    .Q(alu_wait));
 sky130_fd_sc_hd__dfxtp_4 _49575_ (.CLK(clk_0_704),
    .D(_00460_),
    .Q(pcpi_insn[0]));
 sky130_fd_sc_hd__dfxtp_4 _49576_ (.CLK(clk_0_704),
    .D(_00471_),
    .Q(pcpi_insn[1]));
 sky130_fd_sc_hd__dfxtp_4 _49577_ (.CLK(clk_0_704),
    .D(_00482_),
    .Q(pcpi_insn[2]));
 sky130_fd_sc_hd__dfxtp_4 _49578_ (.CLK(clk_0_704),
    .D(_00485_),
    .Q(pcpi_insn[3]));
 sky130_fd_sc_hd__dfxtp_4 _49579_ (.CLK(clk_0_704),
    .D(_00486_),
    .Q(pcpi_insn[4]));
 sky130_fd_sc_hd__dfxtp_4 _49580_ (.CLK(clk_0_704),
    .D(_00487_),
    .Q(pcpi_insn[5]));
 sky130_fd_sc_hd__dfxtp_4 _49581_ (.CLK(clk_0_704),
    .D(_00488_),
    .Q(pcpi_insn[6]));
 sky130_fd_sc_hd__dfxtp_4 _49582_ (.CLK(clk_0_704),
    .D(_00489_),
    .Q(pcpi_insn[7]));
 sky130_fd_sc_hd__dfxtp_4 _49583_ (.CLK(clk_0_704),
    .D(_00490_),
    .Q(pcpi_insn[8]));
 sky130_fd_sc_hd__dfxtp_4 _49584_ (.CLK(clk_0_704),
    .D(_00491_),
    .Q(pcpi_insn[9]));
 sky130_fd_sc_hd__dfxtp_4 _49585_ (.CLK(clk_0_704),
    .D(_00461_),
    .Q(pcpi_insn[10]));
 sky130_fd_sc_hd__dfxtp_4 _49586_ (.CLK(clk_0_704),
    .D(_00462_),
    .Q(pcpi_insn[11]));
 sky130_fd_sc_hd__dfxtp_4 _49587_ (.CLK(clk_0_704),
    .D(_00463_),
    .Q(pcpi_insn[12]));
 sky130_fd_sc_hd__dfxtp_4 _49588_ (.CLK(clk_0_704),
    .D(_00464_),
    .Q(pcpi_insn[13]));
 sky130_fd_sc_hd__dfxtp_4 _49589_ (.CLK(clk_0_704),
    .D(_00465_),
    .Q(pcpi_insn[14]));
 sky130_fd_sc_hd__dfxtp_4 _49590_ (.CLK(clk_0_720),
    .D(_00466_),
    .Q(pcpi_insn[15]));
 sky130_fd_sc_hd__dfxtp_4 _49591_ (.CLK(clk_0_720),
    .D(_00467_),
    .Q(pcpi_insn[16]));
 sky130_fd_sc_hd__dfxtp_4 _49592_ (.CLK(clk_0_720),
    .D(_00468_),
    .Q(pcpi_insn[17]));
 sky130_fd_sc_hd__dfxtp_4 _49593_ (.CLK(clk_0_720),
    .D(_00469_),
    .Q(pcpi_insn[18]));
 sky130_fd_sc_hd__dfxtp_4 _49594_ (.CLK(clk_0_720),
    .D(_00470_),
    .Q(pcpi_insn[19]));
 sky130_fd_sc_hd__dfxtp_4 _49595_ (.CLK(clk_0_720),
    .D(_00472_),
    .Q(pcpi_insn[20]));
 sky130_fd_sc_hd__dfxtp_4 _49596_ (.CLK(clk_0_720),
    .D(_00473_),
    .Q(pcpi_insn[21]));
 sky130_fd_sc_hd__dfxtp_4 _49597_ (.CLK(clk_0_720),
    .D(_00474_),
    .Q(pcpi_insn[22]));
 sky130_fd_sc_hd__dfxtp_4 _49598_ (.CLK(clk_0_720),
    .D(_00475_),
    .Q(pcpi_insn[23]));
 sky130_fd_sc_hd__dfxtp_4 _49599_ (.CLK(clk_0_720),
    .D(_00476_),
    .Q(pcpi_insn[24]));
 sky130_fd_sc_hd__dfxtp_4 _49600_ (.CLK(clk_0_720),
    .D(_00477_),
    .Q(pcpi_insn[25]));
 sky130_fd_sc_hd__dfxtp_4 _49601_ (.CLK(clk_0_720),
    .D(_00478_),
    .Q(pcpi_insn[26]));
 sky130_fd_sc_hd__dfxtp_4 _49602_ (.CLK(clk_0_720),
    .D(_00479_),
    .Q(pcpi_insn[27]));
 sky130_fd_sc_hd__dfxtp_4 _49603_ (.CLK(clk_0_720),
    .D(_00480_),
    .Q(pcpi_insn[28]));
 sky130_fd_sc_hd__dfxtp_4 _49604_ (.CLK(clk_0_720),
    .D(_00481_),
    .Q(pcpi_insn[29]));
 sky130_fd_sc_hd__dfxtp_4 _49605_ (.CLK(clk_0_720),
    .D(_00483_),
    .Q(pcpi_insn[30]));
 sky130_fd_sc_hd__dfxtp_4 _49606_ (.CLK(clk_0_736),
    .D(_00484_),
    .Q(pcpi_insn[31]));
 sky130_fd_sc_hd__dfxtp_4 _49607_ (.CLK(clk_0_736),
    .D(_00265_),
    .Q(instr_lui));
 sky130_fd_sc_hd__dfxtp_4 _49608_ (.CLK(clk_0_736),
    .D(_00250_),
    .Q(instr_auipc));
 sky130_fd_sc_hd__dfxtp_4 _49609_ (.CLK(clk_0_736),
    .D(_00259_),
    .Q(instr_jal));
 sky130_fd_sc_hd__dfxtp_4 _49610_ (.CLK(clk_0_736),
    .D(_00260_),
    .Q(instr_jalr));
 sky130_fd_sc_hd__dfxtp_4 _49611_ (.CLK(clk_0_736),
    .D(_00251_),
    .Q(instr_beq));
 sky130_fd_sc_hd__dfxtp_4 _49612_ (.CLK(clk_0_736),
    .D(_00256_),
    .Q(instr_bne));
 sky130_fd_sc_hd__dfxtp_4 _49613_ (.CLK(clk_0_736),
    .D(_00254_),
    .Q(instr_blt));
 sky130_fd_sc_hd__dfxtp_4 _49614_ (.CLK(clk_0_736),
    .D(_00252_),
    .Q(instr_bge));
 sky130_fd_sc_hd__dfxtp_4 _49615_ (.CLK(clk_0_736),
    .D(_00255_),
    .Q(instr_bltu));
 sky130_fd_sc_hd__dfxtp_4 _49616_ (.CLK(clk_0_736),
    .D(_00253_),
    .Q(instr_bgeu));
 sky130_fd_sc_hd__dfxtp_4 _49617_ (.CLK(clk_0_736),
    .D(_00261_),
    .Q(instr_lb));
 sky130_fd_sc_hd__dfxtp_4 _49618_ (.CLK(clk_0_736),
    .D(_00263_),
    .Q(instr_lh));
 sky130_fd_sc_hd__dfxtp_4 _49619_ (.CLK(clk_0_736),
    .D(_00266_),
    .Q(instr_lw));
 sky130_fd_sc_hd__dfxtp_4 _49620_ (.CLK(clk_0_736),
    .D(_00262_),
    .Q(instr_lbu));
 sky130_fd_sc_hd__dfxtp_4 _49621_ (.CLK(clk_0_736),
    .D(_00264_),
    .Q(instr_lhu));
 sky130_fd_sc_hd__dfxtp_4 _49622_ (.CLK(clk_0_752),
    .D(_00275_),
    .Q(instr_sb));
 sky130_fd_sc_hd__dfxtp_4 _49623_ (.CLK(clk_0_752),
    .D(_00277_),
    .Q(instr_sh));
 sky130_fd_sc_hd__dfxtp_4 _49624_ (.CLK(clk_0_752),
    .D(_00289_),
    .Q(instr_sw));
 sky130_fd_sc_hd__dfxtp_4 _49625_ (.CLK(clk_0_752),
    .D(_00247_),
    .Q(instr_addi));
 sky130_fd_sc_hd__dfxtp_4 _49626_ (.CLK(clk_0_752),
    .D(_00281_),
    .Q(instr_slti));
 sky130_fd_sc_hd__dfxtp_4 _49627_ (.CLK(clk_0_752),
    .D(_00282_),
    .Q(instr_sltiu));
 sky130_fd_sc_hd__dfxtp_4 _49628_ (.CLK(clk_0_752),
    .D(_00293_),
    .Q(instr_xori));
 sky130_fd_sc_hd__dfxtp_4 _49629_ (.CLK(clk_0_752),
    .D(_00269_),
    .Q(instr_ori));
 sky130_fd_sc_hd__dfxtp_4 _49630_ (.CLK(clk_0_752),
    .D(_00249_),
    .Q(instr_andi));
 sky130_fd_sc_hd__dfxtp_4 _49631_ (.CLK(clk_0_752),
    .D(_00279_),
    .Q(instr_slli));
 sky130_fd_sc_hd__dfxtp_4 _49632_ (.CLK(clk_0_752),
    .D(_00287_),
    .Q(instr_srli));
 sky130_fd_sc_hd__dfxtp_4 _49633_ (.CLK(clk_0_752),
    .D(_00285_),
    .Q(instr_srai));
 sky130_fd_sc_hd__dfxtp_4 _49634_ (.CLK(clk_0_752),
    .D(_00246_),
    .Q(instr_add));
 sky130_fd_sc_hd__dfxtp_4 _49635_ (.CLK(clk_0_752),
    .D(_00288_),
    .Q(instr_sub));
 sky130_fd_sc_hd__dfxtp_4 _49636_ (.CLK(clk_0_752),
    .D(_00278_),
    .Q(instr_sll));
 sky130_fd_sc_hd__dfxtp_4 _49637_ (.CLK(clk_0_752),
    .D(_00280_),
    .Q(instr_slt));
 sky130_fd_sc_hd__dfxtp_4 _49638_ (.CLK(clk_0_768),
    .D(_00283_),
    .Q(instr_sltu));
 sky130_fd_sc_hd__dfxtp_4 _49639_ (.CLK(clk_0_768),
    .D(_00292_),
    .Q(instr_xor));
 sky130_fd_sc_hd__dfxtp_4 _49640_ (.CLK(clk_0_768),
    .D(_00286_),
    .Q(instr_srl));
 sky130_fd_sc_hd__dfxtp_4 _49641_ (.CLK(clk_0_768),
    .D(_00284_),
    .Q(instr_sra));
 sky130_fd_sc_hd__dfxtp_4 _49642_ (.CLK(clk_0_768),
    .D(_00268_),
    .Q(instr_or));
 sky130_fd_sc_hd__dfxtp_4 _49643_ (.CLK(clk_0_768),
    .D(_00248_),
    .Q(instr_and));
 sky130_fd_sc_hd__dfxtp_4 _49644_ (.CLK(clk_0_768),
    .D(_00270_),
    .Q(instr_rdcycle));
 sky130_fd_sc_hd__dfxtp_4 _49645_ (.CLK(clk_0_768),
    .D(_00271_),
    .Q(instr_rdcycleh));
 sky130_fd_sc_hd__dfxtp_4 _49646_ (.CLK(clk_0_768),
    .D(_00272_),
    .Q(instr_rdinstr));
 sky130_fd_sc_hd__dfxtp_4 _49647_ (.CLK(clk_0_768),
    .D(_00273_),
    .Q(instr_rdinstrh));
 sky130_fd_sc_hd__dfxtp_4 _49648_ (.CLK(clk_0_768),
    .D(_00257_),
    .Q(instr_ecall_ebreak));
 sky130_fd_sc_hd__dfxtp_4 _49649_ (.CLK(clk_0_768),
    .D(_00258_),
    .Q(instr_getq));
 sky130_fd_sc_hd__dfxtp_4 _49650_ (.CLK(clk_0_768),
    .D(_00276_),
    .Q(instr_setq));
 sky130_fd_sc_hd__dfxtp_4 _49651_ (.CLK(clk_0_768),
    .D(_00274_),
    .Q(instr_retirq));
 sky130_fd_sc_hd__dfxtp_4 _49652_ (.CLK(clk_0_768),
    .D(_00267_),
    .Q(instr_maskirq));
 sky130_fd_sc_hd__dfxtp_4 _49653_ (.CLK(clk_0_768),
    .D(_00291_),
    .Q(instr_waitirq));
 sky130_fd_sc_hd__dfxtp_4 _49654_ (.CLK(clk_0_784),
    .D(_00290_),
    .Q(instr_timer));
 sky130_fd_sc_hd__dfxtp_4 _49655_ (.CLK(clk_0_784),
    .D(_00196_),
    .Q(\decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49656_ (.CLK(clk_0_784),
    .D(_00197_),
    .Q(\decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49657_ (.CLK(clk_0_784),
    .D(_00198_),
    .Q(\decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49658_ (.CLK(clk_0_784),
    .D(_00199_),
    .Q(\decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49659_ (.CLK(clk_0_784),
    .D(_00200_),
    .Q(\decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49660_ (.CLK(clk_0_784),
    .D(_00201_),
    .Q(\decoded_rs1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49661_ (.CLK(clk_0_784),
    .D(_00202_),
    .Q(\decoded_rs1[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49662_ (.CLK(clk_0_784),
    .D(_00203_),
    .Q(\decoded_rs1[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49663_ (.CLK(clk_0_784),
    .D(_00204_),
    .Q(\decoded_rs1[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49664_ (.CLK(clk_0_784),
    .D(_00205_),
    .Q(\decoded_rs1[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49665_ (.CLK(clk_0_784),
    .D(_00206_),
    .Q(\decoded_rs2[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49666_ (.CLK(clk_0_784),
    .D(_00207_),
    .Q(\decoded_rs2[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49667_ (.CLK(clk_0_784),
    .D(_00208_),
    .Q(\decoded_rs2[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49668_ (.CLK(clk_0_784),
    .D(_00209_),
    .Q(\decoded_rs2[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49669_ (.CLK(clk_0_784),
    .D(_00210_),
    .Q(\decoded_rs2[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49670_ (.CLK(clk_0_800),
    .D(_00132_),
    .Q(\decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49671_ (.CLK(clk_0_800),
    .D(_00143_),
    .Q(\decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49672_ (.CLK(clk_0_800),
    .D(_00154_),
    .Q(\decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49673_ (.CLK(clk_0_800),
    .D(_00157_),
    .Q(\decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49674_ (.CLK(clk_0_800),
    .D(_00158_),
    .Q(\decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49675_ (.CLK(clk_0_800),
    .D(_00159_),
    .Q(\decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49676_ (.CLK(clk_0_800),
    .D(_00160_),
    .Q(\decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49677_ (.CLK(clk_0_800),
    .D(_00161_),
    .Q(\decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49678_ (.CLK(clk_0_800),
    .D(_00162_),
    .Q(\decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49679_ (.CLK(clk_0_800),
    .D(_00163_),
    .Q(\decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49680_ (.CLK(clk_0_800),
    .D(_00133_),
    .Q(\decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49681_ (.CLK(clk_0_800),
    .D(_00134_),
    .Q(\decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49682_ (.CLK(clk_0_800),
    .D(_00135_),
    .Q(\decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49683_ (.CLK(clk_0_800),
    .D(_00136_),
    .Q(\decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49684_ (.CLK(clk_0_800),
    .D(_00137_),
    .Q(\decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49685_ (.CLK(clk_0_800),
    .D(_00138_),
    .Q(\decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49686_ (.CLK(clk_0_816),
    .D(_00139_),
    .Q(\decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49687_ (.CLK(clk_0_816),
    .D(_00140_),
    .Q(\decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49688_ (.CLK(clk_0_816),
    .D(_00141_),
    .Q(\decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49689_ (.CLK(clk_0_816),
    .D(_00142_),
    .Q(\decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49690_ (.CLK(clk_0_816),
    .D(_00144_),
    .Q(\decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49691_ (.CLK(clk_0_816),
    .D(_00145_),
    .Q(\decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49692_ (.CLK(clk_0_816),
    .D(_00146_),
    .Q(\decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49693_ (.CLK(clk_0_816),
    .D(_00147_),
    .Q(\decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49694_ (.CLK(clk_0_816),
    .D(_00148_),
    .Q(\decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49695_ (.CLK(clk_0_816),
    .D(_00149_),
    .Q(\decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49696_ (.CLK(clk_0_816),
    .D(_00150_),
    .Q(\decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49697_ (.CLK(clk_0_816),
    .D(_00151_),
    .Q(\decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49698_ (.CLK(clk_0_816),
    .D(_00152_),
    .Q(\decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49699_ (.CLK(clk_0_816),
    .D(_00153_),
    .Q(\decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49700_ (.CLK(clk_0_816),
    .D(_00155_),
    .Q(\decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49701_ (.CLK(clk_0_816),
    .D(_00156_),
    .Q(\decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49702_ (.CLK(clk_0_832),
    .D(_00164_),
    .Q(\decoded_imm_uj[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49703_ (.CLK(clk_0_832),
    .D(_00175_),
    .Q(\decoded_imm_uj[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49704_ (.CLK(clk_0_832),
    .D(_00186_),
    .Q(\decoded_imm_uj[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49705_ (.CLK(clk_0_832),
    .D(_00189_),
    .Q(\decoded_imm_uj[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49706_ (.CLK(clk_0_832),
    .D(_00190_),
    .Q(\decoded_imm_uj[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49707_ (.CLK(clk_0_832),
    .D(_00191_),
    .Q(\decoded_imm_uj[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49708_ (.CLK(clk_0_832),
    .D(_00192_),
    .Q(\decoded_imm_uj[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49709_ (.CLK(clk_0_832),
    .D(_00193_),
    .Q(\decoded_imm_uj[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49710_ (.CLK(clk_0_832),
    .D(_00194_),
    .Q(\decoded_imm_uj[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49711_ (.CLK(clk_0_832),
    .D(_00195_),
    .Q(\decoded_imm_uj[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49712_ (.CLK(clk_0_832),
    .D(_00165_),
    .Q(\decoded_imm_uj[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49713_ (.CLK(clk_0_832),
    .D(_00166_),
    .Q(\decoded_imm_uj[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49714_ (.CLK(clk_0_832),
    .D(_00167_),
    .Q(\decoded_imm_uj[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49715_ (.CLK(clk_0_832),
    .D(_00168_),
    .Q(\decoded_imm_uj[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49716_ (.CLK(clk_0_832),
    .D(_00169_),
    .Q(\decoded_imm_uj[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49717_ (.CLK(clk_0_832),
    .D(_00170_),
    .Q(\decoded_imm_uj[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49718_ (.CLK(clk_0_848),
    .D(_00171_),
    .Q(\decoded_imm_uj[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49719_ (.CLK(clk_0_848),
    .D(_00172_),
    .Q(\decoded_imm_uj[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49720_ (.CLK(clk_0_848),
    .D(_00173_),
    .Q(\decoded_imm_uj[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49721_ (.CLK(clk_0_848),
    .D(_00174_),
    .Q(\decoded_imm_uj[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49722_ (.CLK(clk_0_848),
    .D(_00176_),
    .Q(\decoded_imm_uj[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49723_ (.CLK(clk_0_848),
    .D(_00177_),
    .Q(\decoded_imm_uj[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49724_ (.CLK(clk_0_848),
    .D(_00178_),
    .Q(\decoded_imm_uj[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49725_ (.CLK(clk_0_848),
    .D(_00179_),
    .Q(\decoded_imm_uj[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49726_ (.CLK(clk_0_848),
    .D(_00180_),
    .Q(\decoded_imm_uj[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49727_ (.CLK(clk_0_848),
    .D(_00181_),
    .Q(\decoded_imm_uj[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49728_ (.CLK(clk_0_848),
    .D(_00182_),
    .Q(\decoded_imm_uj[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49729_ (.CLK(clk_0_848),
    .D(_00183_),
    .Q(\decoded_imm_uj[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49730_ (.CLK(clk_0_848),
    .D(_00184_),
    .Q(\decoded_imm_uj[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49731_ (.CLK(clk_0_848),
    .D(_00185_),
    .Q(\decoded_imm_uj[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49732_ (.CLK(clk_0_848),
    .D(_00187_),
    .Q(\decoded_imm_uj[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49733_ (.CLK(clk_0_848),
    .D(_00188_),
    .Q(\decoded_imm_uj[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49734_ (.CLK(clk_0_864),
    .D(_00368_),
    .Q(is_lui_auipc_jal));
 sky130_fd_sc_hd__dfxtp_4 _49735_ (.CLK(clk_0_864),
    .D(_00367_),
    .Q(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__dfxtp_4 _49736_ (.CLK(clk_0_864),
    .D(_00370_),
    .Q(is_slli_srli_srai));
 sky130_fd_sc_hd__dfxtp_4 _49737_ (.CLK(clk_0_864),
    .D(_00366_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
 sky130_fd_sc_hd__dfxtp_4 _49738_ (.CLK(clk_0_864),
    .D(_00369_),
    .Q(is_sb_sh_sw));
 sky130_fd_sc_hd__dfxtp_4 _49739_ (.CLK(clk_0_864),
    .D(_01025_),
    .Q(\cpuregs[18][0] ));
 sky130_fd_sc_hd__dfxtp_4 _49740_ (.CLK(clk_0_864),
    .D(_01036_),
    .Q(\cpuregs[18][1] ));
 sky130_fd_sc_hd__dfxtp_4 _49741_ (.CLK(clk_0_864),
    .D(_01047_),
    .Q(\cpuregs[18][2] ));
 sky130_fd_sc_hd__dfxtp_4 _49742_ (.CLK(clk_0_864),
    .D(_01050_),
    .Q(\cpuregs[18][3] ));
 sky130_fd_sc_hd__dfxtp_4 _49743_ (.CLK(clk_0_864),
    .D(_01051_),
    .Q(\cpuregs[18][4] ));
 sky130_fd_sc_hd__dfxtp_4 _49744_ (.CLK(clk_0_864),
    .D(_01052_),
    .Q(\cpuregs[18][5] ));
 sky130_fd_sc_hd__dfxtp_4 _49745_ (.CLK(clk_0_864),
    .D(_01053_),
    .Q(\cpuregs[18][6] ));
 sky130_fd_sc_hd__dfxtp_4 _49746_ (.CLK(clk_0_864),
    .D(_01054_),
    .Q(\cpuregs[18][7] ));
 sky130_fd_sc_hd__dfxtp_4 _49747_ (.CLK(clk_0_864),
    .D(_01055_),
    .Q(\cpuregs[18][8] ));
 sky130_fd_sc_hd__dfxtp_4 _49748_ (.CLK(clk_0_864),
    .D(_01056_),
    .Q(\cpuregs[18][9] ));
 sky130_fd_sc_hd__dfxtp_4 _49749_ (.CLK(clk_0_864),
    .D(_01026_),
    .Q(\cpuregs[18][10] ));
 sky130_fd_sc_hd__dfxtp_4 _49750_ (.CLK(clk_0_880),
    .D(_01027_),
    .Q(\cpuregs[18][11] ));
 sky130_fd_sc_hd__dfxtp_4 _49751_ (.CLK(clk_0_880),
    .D(_01028_),
    .Q(\cpuregs[18][12] ));
 sky130_fd_sc_hd__dfxtp_4 _49752_ (.CLK(clk_0_880),
    .D(_01029_),
    .Q(\cpuregs[18][13] ));
 sky130_fd_sc_hd__dfxtp_4 _49753_ (.CLK(clk_0_880),
    .D(_01030_),
    .Q(\cpuregs[18][14] ));
 sky130_fd_sc_hd__dfxtp_4 _49754_ (.CLK(clk_0_880),
    .D(_01031_),
    .Q(\cpuregs[18][15] ));
 sky130_fd_sc_hd__dfxtp_4 _49755_ (.CLK(clk_0_880),
    .D(_01032_),
    .Q(\cpuregs[18][16] ));
 sky130_fd_sc_hd__dfxtp_4 _49756_ (.CLK(clk_0_880),
    .D(_01033_),
    .Q(\cpuregs[18][17] ));
 sky130_fd_sc_hd__dfxtp_4 _49757_ (.CLK(clk_0_880),
    .D(_01034_),
    .Q(\cpuregs[18][18] ));
 sky130_fd_sc_hd__dfxtp_4 _49758_ (.CLK(clk_0_880),
    .D(_01035_),
    .Q(\cpuregs[18][19] ));
 sky130_fd_sc_hd__dfxtp_4 _49759_ (.CLK(clk_0_880),
    .D(_01037_),
    .Q(\cpuregs[18][20] ));
 sky130_fd_sc_hd__dfxtp_4 _49760_ (.CLK(clk_0_880),
    .D(_01038_),
    .Q(\cpuregs[18][21] ));
 sky130_fd_sc_hd__dfxtp_4 _49761_ (.CLK(clk_0_880),
    .D(_01039_),
    .Q(\cpuregs[18][22] ));
 sky130_fd_sc_hd__dfxtp_4 _49762_ (.CLK(clk_0_880),
    .D(_01040_),
    .Q(\cpuregs[18][23] ));
 sky130_fd_sc_hd__dfxtp_4 _49763_ (.CLK(clk_0_880),
    .D(_01041_),
    .Q(\cpuregs[18][24] ));
 sky130_fd_sc_hd__dfxtp_4 _49764_ (.CLK(clk_0_880),
    .D(_01042_),
    .Q(\cpuregs[18][25] ));
 sky130_fd_sc_hd__dfxtp_4 _49765_ (.CLK(clk_0_880),
    .D(_01043_),
    .Q(\cpuregs[18][26] ));
 sky130_fd_sc_hd__dfxtp_4 _49766_ (.CLK(clk_0_896),
    .D(_01044_),
    .Q(\cpuregs[18][27] ));
 sky130_fd_sc_hd__dfxtp_4 _49767_ (.CLK(clk_0_896),
    .D(_01045_),
    .Q(\cpuregs[18][28] ));
 sky130_fd_sc_hd__dfxtp_4 _49768_ (.CLK(clk_0_896),
    .D(_01046_),
    .Q(\cpuregs[18][29] ));
 sky130_fd_sc_hd__dfxtp_4 _49769_ (.CLK(clk_0_896),
    .D(_01048_),
    .Q(\cpuregs[18][30] ));
 sky130_fd_sc_hd__dfxtp_4 _49770_ (.CLK(clk_0_896),
    .D(_01049_),
    .Q(\cpuregs[18][31] ));
 sky130_fd_sc_hd__dfxtp_4 _49771_ (.CLK(clk_0_896),
    .D(_00371_),
    .Q(is_slti_blt_slt));
 sky130_fd_sc_hd__dfxtp_4 _49772_ (.CLK(clk_0_896),
    .D(_00372_),
    .Q(is_sltiu_bltu_sltu));
 sky130_fd_sc_hd__dfxtp_4 _49773_ (.CLK(clk_0_896),
    .D(_00364_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__dfxtp_4 _49774_ (.CLK(clk_0_896),
    .D(_00362_),
    .Q(is_alu_reg_imm));
 sky130_fd_sc_hd__dfxtp_4 _49775_ (.CLK(clk_0_896),
    .D(_00363_),
    .Q(is_alu_reg_reg));
 sky130_fd_sc_hd__dfxtp_4 _49776_ (.CLK(clk_0_896),
    .D(_00365_),
    .Q(is_compare));
 sky130_fd_sc_hd__dfxtp_4 _49777_ (.CLK(clk_0_896),
    .D(_00423_),
    .Q(mem_valid));
 sky130_fd_sc_hd__dfxtp_4 _49778_ (.CLK(clk_0_896),
    .D(_00420_),
    .Q(mem_instr));
 sky130_fd_sc_hd__dfxtp_4 _49779_ (.CLK(clk_0_896),
    .D(_00384_),
    .Q(mem_addr[0]));
 sky130_fd_sc_hd__dfxtp_4 _49780_ (.CLK(clk_0_896),
    .D(_00395_),
    .Q(mem_addr[1]));
 sky130_fd_sc_hd__dfxtp_4 _49781_ (.CLK(clk_0_896),
    .D(_00406_),
    .Q(mem_addr[2]));
 sky130_fd_sc_hd__dfxtp_4 _49782_ (.CLK(clk_0_912),
    .D(_00409_),
    .Q(mem_addr[3]));
 sky130_fd_sc_hd__dfxtp_4 _49783_ (.CLK(clk_0_912),
    .D(_00410_),
    .Q(mem_addr[4]));
 sky130_fd_sc_hd__dfxtp_4 _49784_ (.CLK(clk_0_912),
    .D(_00411_),
    .Q(mem_addr[5]));
 sky130_fd_sc_hd__dfxtp_4 _49785_ (.CLK(clk_0_912),
    .D(_00412_),
    .Q(mem_addr[6]));
 sky130_fd_sc_hd__dfxtp_4 _49786_ (.CLK(clk_0_912),
    .D(_00413_),
    .Q(mem_addr[7]));
 sky130_fd_sc_hd__dfxtp_4 _49787_ (.CLK(clk_0_912),
    .D(_00414_),
    .Q(mem_addr[8]));
 sky130_fd_sc_hd__dfxtp_4 _49788_ (.CLK(clk_0_912),
    .D(_00415_),
    .Q(mem_addr[9]));
 sky130_fd_sc_hd__dfxtp_4 _49789_ (.CLK(clk_0_912),
    .D(_00385_),
    .Q(mem_addr[10]));
 sky130_fd_sc_hd__dfxtp_4 _49790_ (.CLK(clk_0_912),
    .D(_00386_),
    .Q(mem_addr[11]));
 sky130_fd_sc_hd__dfxtp_4 _49791_ (.CLK(clk_0_912),
    .D(_00387_),
    .Q(mem_addr[12]));
 sky130_fd_sc_hd__dfxtp_4 _49792_ (.CLK(clk_0_912),
    .D(_00388_),
    .Q(mem_addr[13]));
 sky130_fd_sc_hd__dfxtp_4 _49793_ (.CLK(clk_0_912),
    .D(_00389_),
    .Q(mem_addr[14]));
 sky130_fd_sc_hd__dfxtp_4 _49794_ (.CLK(clk_0_912),
    .D(_00390_),
    .Q(mem_addr[15]));
 sky130_fd_sc_hd__dfxtp_4 _49795_ (.CLK(clk_0_912),
    .D(_00391_),
    .Q(mem_addr[16]));
 sky130_fd_sc_hd__dfxtp_4 _49796_ (.CLK(clk_0_912),
    .D(_00392_),
    .Q(mem_addr[17]));
 sky130_fd_sc_hd__dfxtp_4 _49797_ (.CLK(clk_0_912),
    .D(_00393_),
    .Q(mem_addr[18]));
 sky130_fd_sc_hd__dfxtp_4 _49798_ (.CLK(clk_0_928),
    .D(_00394_),
    .Q(mem_addr[19]));
 sky130_fd_sc_hd__dfxtp_4 _49799_ (.CLK(clk_0_928),
    .D(_00396_),
    .Q(mem_addr[20]));
 sky130_fd_sc_hd__dfxtp_4 _49800_ (.CLK(clk_0_928),
    .D(_00397_),
    .Q(mem_addr[21]));
 sky130_fd_sc_hd__dfxtp_4 _49801_ (.CLK(clk_0_928),
    .D(_00398_),
    .Q(mem_addr[22]));
 sky130_fd_sc_hd__dfxtp_4 _49802_ (.CLK(clk_0_928),
    .D(_00399_),
    .Q(mem_addr[23]));
 sky130_fd_sc_hd__dfxtp_4 _49803_ (.CLK(clk_0_928),
    .D(_00400_),
    .Q(mem_addr[24]));
 sky130_fd_sc_hd__dfxtp_4 _49804_ (.CLK(clk_0_928),
    .D(_00401_),
    .Q(mem_addr[25]));
 sky130_fd_sc_hd__dfxtp_4 _49805_ (.CLK(clk_0_928),
    .D(_00402_),
    .Q(mem_addr[26]));
 sky130_fd_sc_hd__dfxtp_4 _49806_ (.CLK(clk_0_928),
    .D(_00403_),
    .Q(mem_addr[27]));
 sky130_fd_sc_hd__dfxtp_4 _49807_ (.CLK(clk_0_928),
    .D(_00404_),
    .Q(mem_addr[28]));
 sky130_fd_sc_hd__dfxtp_4 _49808_ (.CLK(clk_0_928),
    .D(_00405_),
    .Q(mem_addr[29]));
 sky130_fd_sc_hd__dfxtp_4 _49809_ (.CLK(clk_0_928),
    .D(_00407_),
    .Q(mem_addr[30]));
 sky130_fd_sc_hd__dfxtp_4 _49810_ (.CLK(clk_0_928),
    .D(_00408_),
    .Q(mem_addr[31]));
 sky130_fd_sc_hd__dfxtp_4 _49811_ (.CLK(clk_0_928),
    .D(_00424_),
    .Q(mem_wdata[0]));
 sky130_fd_sc_hd__dfxtp_4 _49812_ (.CLK(clk_0_928),
    .D(_00435_),
    .Q(mem_wdata[1]));
 sky130_fd_sc_hd__dfxtp_4 _49813_ (.CLK(clk_0_928),
    .D(_00446_),
    .Q(mem_wdata[2]));
 sky130_fd_sc_hd__dfxtp_4 _49814_ (.CLK(clk_0_944),
    .D(_00449_),
    .Q(mem_wdata[3]));
 sky130_fd_sc_hd__dfxtp_4 _49815_ (.CLK(clk_0_944),
    .D(_00450_),
    .Q(mem_wdata[4]));
 sky130_fd_sc_hd__dfxtp_4 _49816_ (.CLK(clk_0_944),
    .D(_00451_),
    .Q(mem_wdata[5]));
 sky130_fd_sc_hd__dfxtp_4 _49817_ (.CLK(clk_0_944),
    .D(_00452_),
    .Q(mem_wdata[6]));
 sky130_fd_sc_hd__dfxtp_4 _49818_ (.CLK(clk_0_944),
    .D(_00453_),
    .Q(mem_wdata[7]));
 sky130_fd_sc_hd__dfxtp_4 _49819_ (.CLK(clk_0_944),
    .D(_00454_),
    .Q(mem_wdata[8]));
 sky130_fd_sc_hd__dfxtp_4 _49820_ (.CLK(clk_0_944),
    .D(_00455_),
    .Q(mem_wdata[9]));
 sky130_fd_sc_hd__dfxtp_4 _49821_ (.CLK(clk_0_944),
    .D(_00425_),
    .Q(mem_wdata[10]));
 sky130_fd_sc_hd__dfxtp_4 _49822_ (.CLK(clk_0_944),
    .D(_00426_),
    .Q(mem_wdata[11]));
 sky130_fd_sc_hd__dfxtp_4 _49823_ (.CLK(clk_0_944),
    .D(_00427_),
    .Q(mem_wdata[12]));
 sky130_fd_sc_hd__dfxtp_4 _49824_ (.CLK(clk_0_944),
    .D(_00428_),
    .Q(mem_wdata[13]));
 sky130_fd_sc_hd__dfxtp_4 _49825_ (.CLK(clk_0_944),
    .D(_00429_),
    .Q(mem_wdata[14]));
 sky130_fd_sc_hd__dfxtp_4 _49826_ (.CLK(clk_0_944),
    .D(_00430_),
    .Q(mem_wdata[15]));
 sky130_fd_sc_hd__dfxtp_4 _49827_ (.CLK(clk_0_944),
    .D(_00431_),
    .Q(mem_wdata[16]));
 sky130_fd_sc_hd__dfxtp_4 _49828_ (.CLK(clk_0_944),
    .D(_00432_),
    .Q(mem_wdata[17]));
 sky130_fd_sc_hd__dfxtp_4 _49829_ (.CLK(clk_0_944),
    .D(_00433_),
    .Q(mem_wdata[18]));
 sky130_fd_sc_hd__dfxtp_4 _49830_ (.CLK(clk_0_960),
    .D(_00434_),
    .Q(mem_wdata[19]));
 sky130_fd_sc_hd__dfxtp_4 _49831_ (.CLK(clk_0_960),
    .D(_00436_),
    .Q(mem_wdata[20]));
 sky130_fd_sc_hd__dfxtp_4 _49832_ (.CLK(clk_0_960),
    .D(_00437_),
    .Q(mem_wdata[21]));
 sky130_fd_sc_hd__dfxtp_4 _49833_ (.CLK(clk_0_960),
    .D(_00438_),
    .Q(mem_wdata[22]));
 sky130_fd_sc_hd__dfxtp_4 _49834_ (.CLK(clk_0_960),
    .D(_00439_),
    .Q(mem_wdata[23]));
 sky130_fd_sc_hd__dfxtp_4 _49835_ (.CLK(clk_0_960),
    .D(_00440_),
    .Q(mem_wdata[24]));
 sky130_fd_sc_hd__dfxtp_4 _49836_ (.CLK(clk_0_960),
    .D(_00441_),
    .Q(mem_wdata[25]));
 sky130_fd_sc_hd__dfxtp_4 _49837_ (.CLK(clk_0_960),
    .D(_00442_),
    .Q(mem_wdata[26]));
 sky130_fd_sc_hd__dfxtp_4 _49838_ (.CLK(clk_0_960),
    .D(_00443_),
    .Q(mem_wdata[27]));
 sky130_fd_sc_hd__dfxtp_4 _49839_ (.CLK(clk_0_960),
    .D(_00444_),
    .Q(mem_wdata[28]));
 sky130_fd_sc_hd__dfxtp_4 _49840_ (.CLK(clk_0_960),
    .D(_00445_),
    .Q(mem_wdata[29]));
 sky130_fd_sc_hd__dfxtp_4 _49841_ (.CLK(clk_0_960),
    .D(_00447_),
    .Q(mem_wdata[30]));
 sky130_fd_sc_hd__dfxtp_4 _49842_ (.CLK(clk_0_960),
    .D(_00448_),
    .Q(mem_wdata[31]));
 sky130_fd_sc_hd__dfxtp_4 _49843_ (.CLK(clk_0_960),
    .D(_00456_),
    .Q(mem_wstrb[0]));
 sky130_fd_sc_hd__dfxtp_4 _49844_ (.CLK(clk_0_960),
    .D(_00457_),
    .Q(mem_wstrb[1]));
 sky130_fd_sc_hd__dfxtp_4 _49845_ (.CLK(clk_0_960),
    .D(_00458_),
    .Q(mem_wstrb[2]));
 sky130_fd_sc_hd__dfxtp_4 _49846_ (.CLK(clk_0_976),
    .D(_00459_),
    .Q(mem_wstrb[3]));
 sky130_fd_sc_hd__dfxtp_4 _49847_ (.CLK(clk_0_976),
    .D(_00421_),
    .Q(\mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49848_ (.CLK(clk_0_976),
    .D(_00422_),
    .Q(\mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49849_ (.CLK(clk_0_976),
    .D(_01377_),
    .Q(\alu_add_sub[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49850_ (.CLK(clk_0_976),
    .D(_01388_),
    .Q(\alu_add_sub[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49851_ (.CLK(clk_0_976),
    .D(_01399_),
    .Q(\alu_add_sub[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49852_ (.CLK(clk_0_976),
    .D(_01402_),
    .Q(\alu_add_sub[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49853_ (.CLK(clk_0_976),
    .D(_01403_),
    .Q(\alu_add_sub[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49854_ (.CLK(clk_0_976),
    .D(_01404_),
    .Q(\alu_add_sub[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49855_ (.CLK(clk_0_976),
    .D(_01405_),
    .Q(\alu_add_sub[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49856_ (.CLK(clk_0_976),
    .D(_01406_),
    .Q(\alu_add_sub[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49857_ (.CLK(clk_0_976),
    .D(_01407_),
    .Q(\alu_add_sub[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49858_ (.CLK(clk_0_976),
    .D(_01408_),
    .Q(\alu_add_sub[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49859_ (.CLK(clk_0_976),
    .D(_01378_),
    .Q(\alu_add_sub[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49860_ (.CLK(clk_0_976),
    .D(_01379_),
    .Q(\alu_add_sub[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49861_ (.CLK(clk_0_976),
    .D(_01380_),
    .Q(\alu_add_sub[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49862_ (.CLK(clk_0_992),
    .D(_01381_),
    .Q(\alu_add_sub[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49863_ (.CLK(clk_0_992),
    .D(_01382_),
    .Q(\alu_add_sub[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49864_ (.CLK(clk_0_992),
    .D(_01383_),
    .Q(\alu_add_sub[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49865_ (.CLK(clk_0_992),
    .D(_01384_),
    .Q(\alu_add_sub[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49866_ (.CLK(clk_0_992),
    .D(_01385_),
    .Q(\alu_add_sub[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49867_ (.CLK(clk_0_992),
    .D(_01386_),
    .Q(\alu_add_sub[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49868_ (.CLK(clk_0_992),
    .D(_01387_),
    .Q(\alu_add_sub[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49869_ (.CLK(clk_0_992),
    .D(_01389_),
    .Q(\alu_add_sub[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49870_ (.CLK(clk_0_992),
    .D(_01390_),
    .Q(\alu_add_sub[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49871_ (.CLK(clk_0_992),
    .D(_01391_),
    .Q(\alu_add_sub[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49872_ (.CLK(clk_0_992),
    .D(_01392_),
    .Q(\alu_add_sub[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49873_ (.CLK(clk_0_992),
    .D(_01393_),
    .Q(\alu_add_sub[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49874_ (.CLK(clk_0_992),
    .D(_01394_),
    .Q(\alu_add_sub[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49875_ (.CLK(clk_0_992),
    .D(_01395_),
    .Q(\alu_add_sub[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49876_ (.CLK(clk_0_992),
    .D(_01396_),
    .Q(\alu_add_sub[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49877_ (.CLK(clk_0_992),
    .D(_01397_),
    .Q(\alu_add_sub[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49878_ (.CLK(clk_0_1008),
    .D(_01398_),
    .Q(\alu_add_sub[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49879_ (.CLK(clk_0_1008),
    .D(_01400_),
    .Q(\alu_add_sub[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49880_ (.CLK(clk_0_1008),
    .D(_01401_),
    .Q(\alu_add_sub[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49881_ (.CLK(clk_0_1008),
    .D(_24285_),
    .Q(\alu_shl[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49882_ (.CLK(clk_0_1008),
    .D(_24296_),
    .Q(\alu_shl[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49883_ (.CLK(clk_0_1008),
    .D(_24307_),
    .Q(\alu_shl[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49884_ (.CLK(clk_0_1008),
    .D(_24310_),
    .Q(\alu_shl[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49885_ (.CLK(clk_0_1008),
    .D(_24311_),
    .Q(\alu_shl[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49886_ (.CLK(clk_0_1008),
    .D(_24312_),
    .Q(\alu_shl[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49887_ (.CLK(clk_0_1008),
    .D(_24313_),
    .Q(\alu_shl[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49888_ (.CLK(clk_0_1008),
    .D(_24314_),
    .Q(\alu_shl[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49889_ (.CLK(clk_0_1008),
    .D(_24315_),
    .Q(\alu_shl[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49890_ (.CLK(clk_0_1008),
    .D(_24316_),
    .Q(\alu_shl[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49891_ (.CLK(clk_0_1008),
    .D(_24286_),
    .Q(\alu_shl[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49892_ (.CLK(clk_0_1008),
    .D(_24287_),
    .Q(\alu_shl[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49893_ (.CLK(clk_0_1008),
    .D(_24288_),
    .Q(\alu_shl[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49894_ (.CLK(clk_0_1024),
    .D(_24289_),
    .Q(\alu_shl[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49895_ (.CLK(clk_0_1024),
    .D(_24290_),
    .Q(\alu_shl[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49896_ (.CLK(clk_0_1024),
    .D(_24291_),
    .Q(\alu_shl[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49897_ (.CLK(clk_0_1024),
    .D(_24292_),
    .Q(\alu_shl[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49898_ (.CLK(clk_0_1024),
    .D(_24293_),
    .Q(\alu_shl[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49899_ (.CLK(clk_0_1024),
    .D(_24294_),
    .Q(\alu_shl[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49900_ (.CLK(clk_0_1024),
    .D(_24295_),
    .Q(\alu_shl[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49901_ (.CLK(clk_0_1024),
    .D(_24297_),
    .Q(\alu_shl[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49902_ (.CLK(clk_0_1024),
    .D(_24298_),
    .Q(\alu_shl[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49903_ (.CLK(clk_0_1024),
    .D(_24299_),
    .Q(\alu_shl[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49904_ (.CLK(clk_0_1024),
    .D(_24300_),
    .Q(\alu_shl[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49905_ (.CLK(clk_0_1024),
    .D(_24301_),
    .Q(\alu_shl[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49906_ (.CLK(clk_0_1024),
    .D(_24302_),
    .Q(\alu_shl[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49907_ (.CLK(clk_0_1024),
    .D(_24303_),
    .Q(\alu_shl[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49908_ (.CLK(clk_0_1024),
    .D(_24304_),
    .Q(\alu_shl[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49909_ (.CLK(clk_0_1024),
    .D(_24305_),
    .Q(\alu_shl[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49910_ (.CLK(clk_0_1040),
    .D(_24306_),
    .Q(\alu_shl[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49911_ (.CLK(clk_0_1040),
    .D(_24308_),
    .Q(\alu_shl[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49912_ (.CLK(clk_0_1040),
    .D(_24309_),
    .Q(\alu_shl[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49913_ (.CLK(clk_0_1040),
    .D(_24317_),
    .Q(\alu_shr[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49914_ (.CLK(clk_0_1040),
    .D(_24328_),
    .Q(\alu_shr[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49915_ (.CLK(clk_0_1040),
    .D(_24339_),
    .Q(\alu_shr[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49916_ (.CLK(clk_0_1040),
    .D(_24342_),
    .Q(\alu_shr[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49917_ (.CLK(clk_0_1040),
    .D(_24343_),
    .Q(\alu_shr[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49918_ (.CLK(clk_0_1040),
    .D(_24344_),
    .Q(\alu_shr[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49919_ (.CLK(clk_0_1040),
    .D(_24345_),
    .Q(\alu_shr[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49920_ (.CLK(clk_0_1040),
    .D(_24346_),
    .Q(\alu_shr[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49921_ (.CLK(clk_0_1040),
    .D(_24347_),
    .Q(\alu_shr[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49922_ (.CLK(clk_0_1040),
    .D(_24348_),
    .Q(\alu_shr[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49923_ (.CLK(clk_0_1040),
    .D(_24318_),
    .Q(\alu_shr[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49924_ (.CLK(clk_0_1040),
    .D(_24319_),
    .Q(\alu_shr[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49925_ (.CLK(clk_0_1040),
    .D(_24320_),
    .Q(\alu_shr[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49926_ (.CLK(clk_0_1056),
    .D(_24321_),
    .Q(\alu_shr[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49927_ (.CLK(clk_0_1056),
    .D(_24322_),
    .Q(\alu_shr[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49928_ (.CLK(clk_0_1056),
    .D(_24323_),
    .Q(\alu_shr[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49929_ (.CLK(clk_0_1056),
    .D(_24324_),
    .Q(\alu_shr[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49930_ (.CLK(clk_0_1056),
    .D(_24325_),
    .Q(\alu_shr[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49931_ (.CLK(clk_0_1056),
    .D(_24326_),
    .Q(\alu_shr[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49932_ (.CLK(clk_0_1056),
    .D(_24327_),
    .Q(\alu_shr[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49933_ (.CLK(clk_0_1056),
    .D(_24329_),
    .Q(\alu_shr[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49934_ (.CLK(clk_0_1056),
    .D(_24330_),
    .Q(\alu_shr[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49935_ (.CLK(clk_0_1056),
    .D(_24331_),
    .Q(\alu_shr[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49936_ (.CLK(clk_0_1056),
    .D(_24332_),
    .Q(\alu_shr[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49937_ (.CLK(clk_0_1056),
    .D(_24333_),
    .Q(\alu_shr[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49938_ (.CLK(clk_0_1056),
    .D(_24334_),
    .Q(\alu_shr[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49939_ (.CLK(clk_0_1056),
    .D(_24335_),
    .Q(\alu_shr[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49940_ (.CLK(clk_0_1056),
    .D(_24336_),
    .Q(\alu_shr[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49941_ (.CLK(clk_0_1056),
    .D(_24337_),
    .Q(\alu_shr[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49942_ (.CLK(clk_0_1072),
    .D(_24338_),
    .Q(\alu_shr[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49943_ (.CLK(clk_0_1072),
    .D(_24340_),
    .Q(\alu_shr[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49944_ (.CLK(clk_0_1072),
    .D(_24341_),
    .Q(\alu_shr[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49945_ (.CLK(clk_0_1072),
    .D(_00000_),
    .Q(alu_eq));
 sky130_fd_sc_hd__dfxtp_4 _49946_ (.CLK(clk_0_1072),
    .D(_00002_),
    .Q(alu_ltu));
 sky130_fd_sc_hd__dfxtp_4 _49947_ (.CLK(clk_0_1072),
    .D(_00001_),
    .Q(alu_lts));
 sky130_fd_sc_hd__dfxtp_4 _49948_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[0] ),
    .Q(\mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_4 _49949_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[1] ),
    .Q(\mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_4 _49950_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[2] ),
    .Q(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_4 _49951_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[3] ),
    .Q(\mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_4 _49952_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[4] ),
    .Q(\mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_4 _49953_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[5] ),
    .Q(\mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_4 _49954_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[6] ),
    .Q(\mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_4 _49955_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[7] ),
    .Q(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_4 _49956_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[8] ),
    .Q(\mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_4 _49957_ (.CLK(clk_0_1072),
    .D(\mem_rdata_latched[9] ),
    .Q(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_4 _49958_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[10] ),
    .Q(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_4 _49959_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[11] ),
    .Q(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_4 _49960_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[12] ),
    .Q(\mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_4 _49961_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[13] ),
    .Q(\mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_4 _49962_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[14] ),
    .Q(\mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_4 _49963_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[15] ),
    .Q(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_4 _49964_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[16] ),
    .Q(\mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_4 _49965_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[17] ),
    .Q(\mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_4 _49966_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[18] ),
    .Q(\mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_4 _49967_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[19] ),
    .Q(\mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_4 _49968_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[20] ),
    .Q(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_4 _49969_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[21] ),
    .Q(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_4 _49970_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[22] ),
    .Q(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_4 _49971_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[23] ),
    .Q(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_4 _49972_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[24] ),
    .Q(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_4 _49973_ (.CLK(clk_0_1088),
    .D(\mem_rdata_latched[25] ),
    .Q(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_4 _49974_ (.CLK(clk_0_1104),
    .D(\mem_rdata_latched[26] ),
    .Q(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_4 _49975_ (.CLK(clk_0_1104),
    .D(\mem_rdata_latched[27] ),
    .Q(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_4 _49976_ (.CLK(clk_0_1104),
    .D(\mem_rdata_latched[28] ),
    .Q(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_4 _49977_ (.CLK(clk_0_1104),
    .D(\mem_rdata_latched[29] ),
    .Q(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_4 _49978_ (.CLK(clk_0_1104),
    .D(\mem_rdata_latched[30] ),
    .Q(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_4 _49979_ (.CLK(clk_0_1104),
    .D(\mem_rdata_latched[31] ),
    .Q(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_4 _49980_ (.CLK(clk_0_1104),
    .D(_00769_),
    .Q(\cpuregs[10][0] ));
 sky130_fd_sc_hd__dfxtp_4 _49981_ (.CLK(clk_0_1104),
    .D(_00780_),
    .Q(\cpuregs[10][1] ));
 sky130_fd_sc_hd__dfxtp_4 _49982_ (.CLK(clk_0_1104),
    .D(_00791_),
    .Q(\cpuregs[10][2] ));
 sky130_fd_sc_hd__dfxtp_4 _49983_ (.CLK(clk_0_1104),
    .D(_00794_),
    .Q(\cpuregs[10][3] ));
 sky130_fd_sc_hd__dfxtp_4 _49984_ (.CLK(clk_0_1104),
    .D(_00795_),
    .Q(\cpuregs[10][4] ));
 sky130_fd_sc_hd__dfxtp_4 _49985_ (.CLK(clk_0_1104),
    .D(_00796_),
    .Q(\cpuregs[10][5] ));
 sky130_fd_sc_hd__dfxtp_4 _49986_ (.CLK(clk_0_1104),
    .D(_00797_),
    .Q(\cpuregs[10][6] ));
 sky130_fd_sc_hd__dfxtp_4 _49987_ (.CLK(clk_0_1104),
    .D(_00798_),
    .Q(\cpuregs[10][7] ));
 sky130_fd_sc_hd__dfxtp_4 _49988_ (.CLK(clk_0_1104),
    .D(_00799_),
    .Q(\cpuregs[10][8] ));
 sky130_fd_sc_hd__dfxtp_4 _49989_ (.CLK(clk_0_1104),
    .D(_00800_),
    .Q(\cpuregs[10][9] ));
 sky130_fd_sc_hd__dfxtp_4 _49990_ (.CLK(clk_0_1120),
    .D(_00770_),
    .Q(\cpuregs[10][10] ));
 sky130_fd_sc_hd__dfxtp_4 _49991_ (.CLK(clk_0_1120),
    .D(_00771_),
    .Q(\cpuregs[10][11] ));
 sky130_fd_sc_hd__dfxtp_4 _49992_ (.CLK(clk_0_1120),
    .D(_00772_),
    .Q(\cpuregs[10][12] ));
 sky130_fd_sc_hd__dfxtp_4 _49993_ (.CLK(clk_0_1120),
    .D(_00773_),
    .Q(\cpuregs[10][13] ));
 sky130_fd_sc_hd__dfxtp_4 _49994_ (.CLK(clk_0_1120),
    .D(_00774_),
    .Q(\cpuregs[10][14] ));
 sky130_fd_sc_hd__dfxtp_4 _49995_ (.CLK(clk_0_1120),
    .D(_00775_),
    .Q(\cpuregs[10][15] ));
 sky130_fd_sc_hd__dfxtp_4 _49996_ (.CLK(clk_0_1120),
    .D(_00776_),
    .Q(\cpuregs[10][16] ));
 sky130_fd_sc_hd__dfxtp_4 _49997_ (.CLK(clk_0_1120),
    .D(_00777_),
    .Q(\cpuregs[10][17] ));
 sky130_fd_sc_hd__dfxtp_4 _49998_ (.CLK(clk_0_1120),
    .D(_00778_),
    .Q(\cpuregs[10][18] ));
 sky130_fd_sc_hd__dfxtp_4 _49999_ (.CLK(clk_0_1120),
    .D(_00779_),
    .Q(\cpuregs[10][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50000_ (.CLK(clk_0_1120),
    .D(_00781_),
    .Q(\cpuregs[10][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50001_ (.CLK(clk_0_1120),
    .D(_00782_),
    .Q(\cpuregs[10][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50002_ (.CLK(clk_0_1120),
    .D(_00783_),
    .Q(\cpuregs[10][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50003_ (.CLK(clk_0_1120),
    .D(_00784_),
    .Q(\cpuregs[10][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50004_ (.CLK(clk_0_1120),
    .D(_00785_),
    .Q(\cpuregs[10][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50005_ (.CLK(clk_0_1120),
    .D(_00786_),
    .Q(\cpuregs[10][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50006_ (.CLK(clk_0_1136),
    .D(_00787_),
    .Q(\cpuregs[10][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50007_ (.CLK(clk_0_1136),
    .D(_00788_),
    .Q(\cpuregs[10][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50008_ (.CLK(clk_0_1136),
    .D(_00789_),
    .Q(\cpuregs[10][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50009_ (.CLK(clk_0_1136),
    .D(_00790_),
    .Q(\cpuregs[10][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50010_ (.CLK(clk_0_1136),
    .D(_00792_),
    .Q(\cpuregs[10][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50011_ (.CLK(clk_0_1136),
    .D(_00793_),
    .Q(\cpuregs[10][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50012_ (.CLK(clk_0_1136),
    .D(_01409_),
    .Q(\pcpi_mul.rd[0] ));
 sky130_fd_sc_hd__dfxtp_4 _50013_ (.CLK(clk_0_1136),
    .D(_01410_),
    .Q(\pcpi_mul.rd[1] ));
 sky130_fd_sc_hd__dfxtp_4 _50014_ (.CLK(clk_0_1136),
    .D(_01411_),
    .Q(\pcpi_mul.rd[2] ));
 sky130_fd_sc_hd__dfxtp_4 _50015_ (.CLK(clk_0_1136),
    .D(_01412_),
    .Q(\pcpi_mul.rd[3] ));
 sky130_fd_sc_hd__dfxtp_4 _50016_ (.CLK(clk_0_1136),
    .D(_01413_),
    .Q(\pcpi_mul.rd[4] ));
 sky130_fd_sc_hd__dfxtp_4 _50017_ (.CLK(clk_0_1136),
    .D(_01414_),
    .Q(\pcpi_mul.rd[5] ));
 sky130_fd_sc_hd__dfxtp_4 _50018_ (.CLK(clk_0_1136),
    .D(_01469_),
    .Q(\pcpi_mul.rd[6] ));
 sky130_fd_sc_hd__dfxtp_4 _50019_ (.CLK(clk_0_1136),
    .D(_01470_),
    .Q(\pcpi_mul.rd[7] ));
 sky130_fd_sc_hd__dfxtp_4 _50020_ (.CLK(clk_0_1136),
    .D(_01471_),
    .Q(\pcpi_mul.rd[8] ));
 sky130_fd_sc_hd__dfxtp_4 _50021_ (.CLK(clk_0_1136),
    .D(_01472_),
    .Q(\pcpi_mul.rd[9] ));
 sky130_fd_sc_hd__dfxtp_4 _50022_ (.CLK(clk_0_1152),
    .D(_01415_),
    .Q(\pcpi_mul.rd[10] ));
 sky130_fd_sc_hd__dfxtp_4 _50023_ (.CLK(clk_0_1152),
    .D(_01416_),
    .Q(\pcpi_mul.rd[11] ));
 sky130_fd_sc_hd__dfxtp_4 _50024_ (.CLK(clk_0_1152),
    .D(_01417_),
    .Q(\pcpi_mul.rd[12] ));
 sky130_fd_sc_hd__dfxtp_4 _50025_ (.CLK(clk_0_1152),
    .D(_01418_),
    .Q(\pcpi_mul.rd[13] ));
 sky130_fd_sc_hd__dfxtp_4 _50026_ (.CLK(clk_0_1152),
    .D(_01419_),
    .Q(\pcpi_mul.rd[14] ));
 sky130_fd_sc_hd__dfxtp_4 _50027_ (.CLK(clk_0_1152),
    .D(_01420_),
    .Q(\pcpi_mul.rd[15] ));
 sky130_fd_sc_hd__dfxtp_4 _50028_ (.CLK(clk_0_1152),
    .D(_01421_),
    .Q(\pcpi_mul.rd[16] ));
 sky130_fd_sc_hd__dfxtp_4 _50029_ (.CLK(clk_0_1152),
    .D(_01422_),
    .Q(\pcpi_mul.rd[17] ));
 sky130_fd_sc_hd__dfxtp_4 _50030_ (.CLK(clk_0_1152),
    .D(_01423_),
    .Q(\pcpi_mul.rd[18] ));
 sky130_fd_sc_hd__dfxtp_4 _50031_ (.CLK(clk_0_1152),
    .D(_01424_),
    .Q(\pcpi_mul.rd[19] ));
 sky130_fd_sc_hd__dfxtp_4 _50032_ (.CLK(clk_0_1152),
    .D(_01425_),
    .Q(\pcpi_mul.rd[20] ));
 sky130_fd_sc_hd__dfxtp_4 _50033_ (.CLK(clk_0_1152),
    .D(_01426_),
    .Q(\pcpi_mul.rd[21] ));
 sky130_fd_sc_hd__dfxtp_4 _50034_ (.CLK(clk_0_1152),
    .D(_01427_),
    .Q(\pcpi_mul.rd[22] ));
 sky130_fd_sc_hd__dfxtp_4 _50035_ (.CLK(clk_0_1152),
    .D(_01428_),
    .Q(\pcpi_mul.rd[23] ));
 sky130_fd_sc_hd__dfxtp_4 _50036_ (.CLK(clk_0_1152),
    .D(_01429_),
    .Q(\pcpi_mul.rd[24] ));
 sky130_fd_sc_hd__dfxtp_4 _50037_ (.CLK(clk_0_1152),
    .D(_01430_),
    .Q(\pcpi_mul.rd[25] ));
 sky130_fd_sc_hd__dfxtp_4 _50038_ (.CLK(clk_0_1168),
    .D(_01431_),
    .Q(\pcpi_mul.rd[26] ));
 sky130_fd_sc_hd__dfxtp_4 _50039_ (.CLK(clk_0_1168),
    .D(_01432_),
    .Q(\pcpi_mul.rd[27] ));
 sky130_fd_sc_hd__dfxtp_4 _50040_ (.CLK(clk_0_1168),
    .D(_01433_),
    .Q(\pcpi_mul.rd[28] ));
 sky130_fd_sc_hd__dfxtp_4 _50041_ (.CLK(clk_0_1168),
    .D(_01434_),
    .Q(\pcpi_mul.rd[29] ));
 sky130_fd_sc_hd__dfxtp_4 _50042_ (.CLK(clk_0_1168),
    .D(_01435_),
    .Q(\pcpi_mul.rd[30] ));
 sky130_fd_sc_hd__dfxtp_4 _50043_ (.CLK(clk_0_1168),
    .D(_01436_),
    .Q(\pcpi_mul.rd[31] ));
 sky130_fd_sc_hd__dfxtp_4 _50044_ (.CLK(clk_0_1168),
    .D(_01437_),
    .Q(\pcpi_mul.rd[32] ));
 sky130_fd_sc_hd__dfxtp_4 _50045_ (.CLK(clk_0_1168),
    .D(_01438_),
    .Q(\pcpi_mul.rd[33] ));
 sky130_fd_sc_hd__dfxtp_4 _50046_ (.CLK(clk_0_1168),
    .D(_01439_),
    .Q(\pcpi_mul.rd[34] ));
 sky130_fd_sc_hd__dfxtp_4 _50047_ (.CLK(clk_0_1168),
    .D(_01440_),
    .Q(\pcpi_mul.rd[35] ));
 sky130_fd_sc_hd__dfxtp_4 _50048_ (.CLK(clk_0_1168),
    .D(_01441_),
    .Q(\pcpi_mul.rd[36] ));
 sky130_fd_sc_hd__dfxtp_4 _50049_ (.CLK(clk_0_1168),
    .D(_01442_),
    .Q(\pcpi_mul.rd[37] ));
 sky130_fd_sc_hd__dfxtp_4 _50050_ (.CLK(clk_0_1168),
    .D(_01443_),
    .Q(\pcpi_mul.rd[38] ));
 sky130_fd_sc_hd__dfxtp_4 _50051_ (.CLK(clk_0_1168),
    .D(_01444_),
    .Q(\pcpi_mul.rd[39] ));
 sky130_fd_sc_hd__dfxtp_4 _50052_ (.CLK(clk_0_1168),
    .D(_01445_),
    .Q(\pcpi_mul.rd[40] ));
 sky130_fd_sc_hd__dfxtp_4 _50053_ (.CLK(clk_0_1168),
    .D(_01446_),
    .Q(\pcpi_mul.rd[41] ));
 sky130_fd_sc_hd__dfxtp_4 _50054_ (.CLK(clk_0_1184),
    .D(_01447_),
    .Q(\pcpi_mul.rd[42] ));
 sky130_fd_sc_hd__dfxtp_4 _50055_ (.CLK(clk_0_1184),
    .D(_01448_),
    .Q(\pcpi_mul.rd[43] ));
 sky130_fd_sc_hd__dfxtp_4 _50056_ (.CLK(clk_0_1184),
    .D(_01449_),
    .Q(\pcpi_mul.rd[44] ));
 sky130_fd_sc_hd__dfxtp_4 _50057_ (.CLK(clk_0_1184),
    .D(_01450_),
    .Q(\pcpi_mul.rd[45] ));
 sky130_fd_sc_hd__dfxtp_4 _50058_ (.CLK(clk_0_1184),
    .D(_01451_),
    .Q(\pcpi_mul.rd[46] ));
 sky130_fd_sc_hd__dfxtp_4 _50059_ (.CLK(clk_0_1184),
    .D(_01452_),
    .Q(\pcpi_mul.rd[47] ));
 sky130_fd_sc_hd__dfxtp_4 _50060_ (.CLK(clk_0_1184),
    .D(_01453_),
    .Q(\pcpi_mul.rd[48] ));
 sky130_fd_sc_hd__dfxtp_4 _50061_ (.CLK(clk_0_1184),
    .D(_01454_),
    .Q(\pcpi_mul.rd[49] ));
 sky130_fd_sc_hd__dfxtp_4 _50062_ (.CLK(clk_0_1184),
    .D(_01455_),
    .Q(\pcpi_mul.rd[50] ));
 sky130_fd_sc_hd__dfxtp_4 _50063_ (.CLK(clk_0_1184),
    .D(_01456_),
    .Q(\pcpi_mul.rd[51] ));
 sky130_fd_sc_hd__dfxtp_4 _50064_ (.CLK(clk_0_1184),
    .D(_01457_),
    .Q(\pcpi_mul.rd[52] ));
 sky130_fd_sc_hd__dfxtp_4 _50065_ (.CLK(clk_0_1184),
    .D(_01458_),
    .Q(\pcpi_mul.rd[53] ));
 sky130_fd_sc_hd__dfxtp_4 _50066_ (.CLK(clk_0_1184),
    .D(_01459_),
    .Q(\pcpi_mul.rd[54] ));
 sky130_fd_sc_hd__dfxtp_4 _50067_ (.CLK(clk_0_1184),
    .D(_01460_),
    .Q(\pcpi_mul.rd[55] ));
 sky130_fd_sc_hd__dfxtp_4 _50068_ (.CLK(clk_0_1184),
    .D(_01461_),
    .Q(\pcpi_mul.rd[56] ));
 sky130_fd_sc_hd__dfxtp_4 _50069_ (.CLK(clk_0_1184),
    .D(_01462_),
    .Q(\pcpi_mul.rd[57] ));
 sky130_fd_sc_hd__dfxtp_4 _50070_ (.CLK(clk_0_1200),
    .D(_01463_),
    .Q(\pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__dfxtp_4 _50071_ (.CLK(clk_0_1200),
    .D(_01464_),
    .Q(\pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__dfxtp_4 _50072_ (.CLK(clk_0_1200),
    .D(_01465_),
    .Q(\pcpi_mul.rd[60] ));
 sky130_fd_sc_hd__dfxtp_4 _50073_ (.CLK(clk_0_1200),
    .D(_01466_),
    .Q(\pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__dfxtp_4 _50074_ (.CLK(clk_0_1200),
    .D(_01467_),
    .Q(\pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__dfxtp_4 _50075_ (.CLK(clk_0_1200),
    .D(_01468_),
    .Q(\pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__dfxtp_4 _50076_ (.CLK(clk_0_1200),
    .D(_00669_),
    .Q(\pcpi_mul.active[0] ));
 sky130_fd_sc_hd__dfxtp_4 _50077_ (.CLK(clk_0_1200),
    .D(_00670_),
    .Q(\pcpi_mul.active[1] ));
 sky130_fd_sc_hd__dfxtp_4 _50078_ (.CLK(clk_0_1200),
    .D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ));
 sky130_fd_sc_hd__dfxtp_4 _50079_ (.CLK(clk_0_1200),
    .D(_00704_),
    .Q(\pcpi_mul.rs2[0] ));
 sky130_fd_sc_hd__dfxtp_4 _50080_ (.CLK(clk_0_1200),
    .D(_00715_),
    .Q(\pcpi_mul.rs2[1] ));
 sky130_fd_sc_hd__dfxtp_4 _50081_ (.CLK(clk_0_1200),
    .D(_00726_),
    .Q(\pcpi_mul.rs2[2] ));
 sky130_fd_sc_hd__dfxtp_4 _50082_ (.CLK(clk_0_1200),
    .D(_00730_),
    .Q(\pcpi_mul.rs2[3] ));
 sky130_fd_sc_hd__dfxtp_4 _50083_ (.CLK(clk_0_1200),
    .D(_00731_),
    .Q(\pcpi_mul.rs2[4] ));
 sky130_fd_sc_hd__dfxtp_4 _50084_ (.CLK(clk_0_1200),
    .D(_00732_),
    .Q(\pcpi_mul.rs2[5] ));
 sky130_fd_sc_hd__dfxtp_4 _50085_ (.CLK(clk_0_1200),
    .D(_00733_),
    .Q(\pcpi_mul.rs2[6] ));
 sky130_fd_sc_hd__dfxtp_4 _50086_ (.CLK(clk_0_1216),
    .D(_00734_),
    .Q(\pcpi_mul.rs2[7] ));
 sky130_fd_sc_hd__dfxtp_4 _50087_ (.CLK(clk_0_1216),
    .D(_00735_),
    .Q(\pcpi_mul.rs2[8] ));
 sky130_fd_sc_hd__dfxtp_4 _50088_ (.CLK(clk_0_1216),
    .D(_00736_),
    .Q(\pcpi_mul.rs2[9] ));
 sky130_fd_sc_hd__dfxtp_4 _50089_ (.CLK(clk_0_1216),
    .D(_00705_),
    .Q(\pcpi_mul.rs2[10] ));
 sky130_fd_sc_hd__dfxtp_4 _50090_ (.CLK(clk_0_1216),
    .D(_00706_),
    .Q(\pcpi_mul.rs2[11] ));
 sky130_fd_sc_hd__dfxtp_4 _50091_ (.CLK(clk_0_1216),
    .D(_00707_),
    .Q(\pcpi_mul.rs2[12] ));
 sky130_fd_sc_hd__dfxtp_4 _50092_ (.CLK(clk_0_1216),
    .D(_00708_),
    .Q(\pcpi_mul.rs2[13] ));
 sky130_fd_sc_hd__dfxtp_4 _50093_ (.CLK(clk_0_1216),
    .D(_00709_),
    .Q(\pcpi_mul.rs2[14] ));
 sky130_fd_sc_hd__dfxtp_4 _50094_ (.CLK(clk_0_1216),
    .D(_00710_),
    .Q(\pcpi_mul.rs2[15] ));
 sky130_fd_sc_hd__dfxtp_4 _50095_ (.CLK(clk_0_1216),
    .D(_00711_),
    .Q(\pcpi_mul.rs2[16] ));
 sky130_fd_sc_hd__dfxtp_4 _50096_ (.CLK(clk_0_1216),
    .D(_00712_),
    .Q(\pcpi_mul.rs2[17] ));
 sky130_fd_sc_hd__dfxtp_4 _50097_ (.CLK(clk_0_1216),
    .D(_00713_),
    .Q(\pcpi_mul.rs2[18] ));
 sky130_fd_sc_hd__dfxtp_4 _50098_ (.CLK(clk_0_1216),
    .D(_00714_),
    .Q(\pcpi_mul.rs2[19] ));
 sky130_fd_sc_hd__dfxtp_4 _50099_ (.CLK(clk_0_1216),
    .D(_00716_),
    .Q(\pcpi_mul.rs2[20] ));
 sky130_fd_sc_hd__dfxtp_4 _50100_ (.CLK(clk_0_1216),
    .D(_00717_),
    .Q(\pcpi_mul.rs2[21] ));
 sky130_fd_sc_hd__dfxtp_4 _50101_ (.CLK(clk_0_1216),
    .D(_00718_),
    .Q(\pcpi_mul.rs2[22] ));
 sky130_fd_sc_hd__dfxtp_4 _50102_ (.CLK(clk_0_1232),
    .D(_00719_),
    .Q(\pcpi_mul.rs2[23] ));
 sky130_fd_sc_hd__dfxtp_4 _50103_ (.CLK(clk_0_1232),
    .D(_00720_),
    .Q(\pcpi_mul.rs2[24] ));
 sky130_fd_sc_hd__dfxtp_4 _50104_ (.CLK(clk_0_1232),
    .D(_00721_),
    .Q(\pcpi_mul.rs2[25] ));
 sky130_fd_sc_hd__dfxtp_4 _50105_ (.CLK(clk_0_1232),
    .D(_00722_),
    .Q(\pcpi_mul.rs2[26] ));
 sky130_fd_sc_hd__dfxtp_4 _50106_ (.CLK(clk_0_1232),
    .D(_00723_),
    .Q(\pcpi_mul.rs2[27] ));
 sky130_fd_sc_hd__dfxtp_4 _50107_ (.CLK(clk_0_1232),
    .D(_00724_),
    .Q(\pcpi_mul.rs2[28] ));
 sky130_fd_sc_hd__dfxtp_4 _50108_ (.CLK(clk_0_1232),
    .D(_00725_),
    .Q(\pcpi_mul.rs2[29] ));
 sky130_fd_sc_hd__dfxtp_4 _50109_ (.CLK(clk_0_1232),
    .D(_00727_),
    .Q(\pcpi_mul.rs2[30] ));
 sky130_fd_sc_hd__dfxtp_4 _50110_ (.CLK(clk_0_1232),
    .D(_00728_),
    .Q(\pcpi_mul.rs2[31] ));
 sky130_fd_sc_hd__dfxtp_4 _50111_ (.CLK(clk_0_1232),
    .D(_00729_),
    .Q(\pcpi_mul.rs2[32] ));
 sky130_fd_sc_hd__dfxtp_4 _50112_ (.CLK(clk_0_1232),
    .D(_00671_),
    .Q(\pcpi_mul.rs1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _50113_ (.CLK(clk_0_1232),
    .D(_00682_),
    .Q(\pcpi_mul.rs1[1] ));
 sky130_fd_sc_hd__dfxtp_4 _50114_ (.CLK(clk_0_1232),
    .D(_00693_),
    .Q(\pcpi_mul.rs1[2] ));
 sky130_fd_sc_hd__dfxtp_4 _50115_ (.CLK(clk_0_1232),
    .D(_00697_),
    .Q(\pcpi_mul.rs1[3] ));
 sky130_fd_sc_hd__dfxtp_4 _50116_ (.CLK(clk_0_1232),
    .D(_00698_),
    .Q(\pcpi_mul.rs1[4] ));
 sky130_fd_sc_hd__dfxtp_4 _50117_ (.CLK(clk_0_1232),
    .D(_00699_),
    .Q(\pcpi_mul.rs1[5] ));
 sky130_fd_sc_hd__dfxtp_4 _50118_ (.CLK(clk_0_1248),
    .D(_00700_),
    .Q(\pcpi_mul.rs1[6] ));
 sky130_fd_sc_hd__dfxtp_4 _50119_ (.CLK(clk_0_1248),
    .D(_00701_),
    .Q(\pcpi_mul.rs1[7] ));
 sky130_fd_sc_hd__dfxtp_4 _50120_ (.CLK(clk_0_1248),
    .D(_00702_),
    .Q(\pcpi_mul.rs1[8] ));
 sky130_fd_sc_hd__dfxtp_4 _50121_ (.CLK(clk_0_1248),
    .D(_00703_),
    .Q(\pcpi_mul.rs1[9] ));
 sky130_fd_sc_hd__dfxtp_4 _50122_ (.CLK(clk_0_1248),
    .D(_00672_),
    .Q(\pcpi_mul.rs1[10] ));
 sky130_fd_sc_hd__dfxtp_4 _50123_ (.CLK(clk_0_1248),
    .D(_00673_),
    .Q(\pcpi_mul.rs1[11] ));
 sky130_fd_sc_hd__dfxtp_4 _50124_ (.CLK(clk_0_1248),
    .D(_00674_),
    .Q(\pcpi_mul.rs1[12] ));
 sky130_fd_sc_hd__dfxtp_4 _50125_ (.CLK(clk_0_1248),
    .D(_00675_),
    .Q(\pcpi_mul.rs1[13] ));
 sky130_fd_sc_hd__dfxtp_4 _50126_ (.CLK(clk_0_1248),
    .D(_00676_),
    .Q(\pcpi_mul.rs1[14] ));
 sky130_fd_sc_hd__dfxtp_4 _50127_ (.CLK(clk_0_1248),
    .D(_00677_),
    .Q(\pcpi_mul.rs1[15] ));
 sky130_fd_sc_hd__dfxtp_4 _50128_ (.CLK(clk_0_1248),
    .D(_00678_),
    .Q(\pcpi_mul.rs1[16] ));
 sky130_fd_sc_hd__dfxtp_4 _50129_ (.CLK(clk_0_1248),
    .D(_00679_),
    .Q(\pcpi_mul.rs1[17] ));
 sky130_fd_sc_hd__dfxtp_4 _50130_ (.CLK(clk_0_1248),
    .D(_00680_),
    .Q(\pcpi_mul.rs1[18] ));
 sky130_fd_sc_hd__dfxtp_4 _50131_ (.CLK(clk_0_1248),
    .D(_00681_),
    .Q(\pcpi_mul.rs1[19] ));
 sky130_fd_sc_hd__dfxtp_4 _50132_ (.CLK(clk_0_1248),
    .D(_00683_),
    .Q(\pcpi_mul.rs1[20] ));
 sky130_fd_sc_hd__dfxtp_4 _50133_ (.CLK(clk_0_1248),
    .D(_00684_),
    .Q(\pcpi_mul.rs1[21] ));
 sky130_fd_sc_hd__dfxtp_4 _50134_ (.CLK(clk_0_1264),
    .D(_00685_),
    .Q(\pcpi_mul.rs1[22] ));
 sky130_fd_sc_hd__dfxtp_4 _50135_ (.CLK(clk_0_1264),
    .D(_00686_),
    .Q(\pcpi_mul.rs1[23] ));
 sky130_fd_sc_hd__dfxtp_4 _50136_ (.CLK(clk_0_1264),
    .D(_00687_),
    .Q(\pcpi_mul.rs1[24] ));
 sky130_fd_sc_hd__dfxtp_4 _50137_ (.CLK(clk_0_1264),
    .D(_00688_),
    .Q(\pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__dfxtp_4 _50138_ (.CLK(clk_0_1264),
    .D(_00689_),
    .Q(\pcpi_mul.rs1[26] ));
 sky130_fd_sc_hd__dfxtp_4 _50139_ (.CLK(clk_0_1264),
    .D(_00690_),
    .Q(\pcpi_mul.rs1[27] ));
 sky130_fd_sc_hd__dfxtp_4 _50140_ (.CLK(clk_0_1264),
    .D(_00691_),
    .Q(\pcpi_mul.rs1[28] ));
 sky130_fd_sc_hd__dfxtp_4 _50141_ (.CLK(clk_0_1264),
    .D(_00692_),
    .Q(\pcpi_mul.rs1[29] ));
 sky130_fd_sc_hd__dfxtp_4 _50142_ (.CLK(clk_0_1264),
    .D(_00694_),
    .Q(\pcpi_mul.rs1[30] ));
 sky130_fd_sc_hd__dfxtp_4 _50143_ (.CLK(clk_0_1264),
    .D(_00695_),
    .Q(\pcpi_mul.rs1[31] ));
 sky130_fd_sc_hd__dfxtp_4 _50144_ (.CLK(clk_0_1264),
    .D(_00696_),
    .Q(\pcpi_mul.rs1[32] ));
 sky130_fd_sc_hd__dfxtp_4 _50145_ (.CLK(clk_0_1264),
    .D(_00993_),
    .Q(\cpuregs[17][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50146_ (.CLK(clk_0_1264),
    .D(_01004_),
    .Q(\cpuregs[17][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50147_ (.CLK(clk_0_1264),
    .D(_01015_),
    .Q(\cpuregs[17][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50148_ (.CLK(clk_0_1264),
    .D(_01018_),
    .Q(\cpuregs[17][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50149_ (.CLK(clk_0_1264),
    .D(_01019_),
    .Q(\cpuregs[17][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50150_ (.CLK(clk_0_1280),
    .D(_01020_),
    .Q(\cpuregs[17][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50151_ (.CLK(clk_0_1280),
    .D(_01021_),
    .Q(\cpuregs[17][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50152_ (.CLK(clk_0_1280),
    .D(_01022_),
    .Q(\cpuregs[17][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50153_ (.CLK(clk_0_1280),
    .D(_01023_),
    .Q(\cpuregs[17][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50154_ (.CLK(clk_0_1280),
    .D(_01024_),
    .Q(\cpuregs[17][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50155_ (.CLK(clk_0_1280),
    .D(_00994_),
    .Q(\cpuregs[17][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50156_ (.CLK(clk_0_1280),
    .D(_00995_),
    .Q(\cpuregs[17][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50157_ (.CLK(clk_0_1280),
    .D(_00996_),
    .Q(\cpuregs[17][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50158_ (.CLK(clk_0_1280),
    .D(_00997_),
    .Q(\cpuregs[17][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50159_ (.CLK(clk_0_1280),
    .D(_00998_),
    .Q(\cpuregs[17][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50160_ (.CLK(clk_0_1280),
    .D(_00999_),
    .Q(\cpuregs[17][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50161_ (.CLK(clk_0_1280),
    .D(_01000_),
    .Q(\cpuregs[17][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50162_ (.CLK(clk_0_1280),
    .D(_01001_),
    .Q(\cpuregs[17][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50163_ (.CLK(clk_0_1280),
    .D(_01002_),
    .Q(\cpuregs[17][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50164_ (.CLK(clk_0_1280),
    .D(_01003_),
    .Q(\cpuregs[17][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50165_ (.CLK(clk_0_1280),
    .D(_01005_),
    .Q(\cpuregs[17][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50166_ (.CLK(clk_0_1296),
    .D(_01006_),
    .Q(\cpuregs[17][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50167_ (.CLK(clk_0_1296),
    .D(_01007_),
    .Q(\cpuregs[17][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50168_ (.CLK(clk_0_1296),
    .D(_01008_),
    .Q(\cpuregs[17][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50169_ (.CLK(clk_0_1296),
    .D(_01009_),
    .Q(\cpuregs[17][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50170_ (.CLK(clk_0_1296),
    .D(_01010_),
    .Q(\cpuregs[17][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50171_ (.CLK(clk_0_1296),
    .D(_01011_),
    .Q(\cpuregs[17][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50172_ (.CLK(clk_0_1296),
    .D(_01012_),
    .Q(\cpuregs[17][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50173_ (.CLK(clk_0_1296),
    .D(_01013_),
    .Q(\cpuregs[17][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50174_ (.CLK(clk_0_1296),
    .D(_01014_),
    .Q(\cpuregs[17][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50175_ (.CLK(clk_0_1296),
    .D(_01016_),
    .Q(\cpuregs[17][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50176_ (.CLK(clk_0_1296),
    .D(_01017_),
    .Q(\cpuregs[17][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50177_ (.CLK(clk_0_1296),
    .D(_01185_),
    .Q(\cpuregs[4][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50178_ (.CLK(clk_0_1296),
    .D(_01196_),
    .Q(\cpuregs[4][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50179_ (.CLK(clk_0_1296),
    .D(_01207_),
    .Q(\cpuregs[4][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50180_ (.CLK(clk_0_1296),
    .D(_01210_),
    .Q(\cpuregs[4][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50181_ (.CLK(clk_0_1296),
    .D(_01211_),
    .Q(\cpuregs[4][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50182_ (.CLK(clk_0_1312),
    .D(_01212_),
    .Q(\cpuregs[4][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50183_ (.CLK(clk_0_1312),
    .D(_01213_),
    .Q(\cpuregs[4][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50184_ (.CLK(clk_0_1312),
    .D(_01214_),
    .Q(\cpuregs[4][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50185_ (.CLK(clk_0_1312),
    .D(_01215_),
    .Q(\cpuregs[4][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50186_ (.CLK(clk_0_1312),
    .D(_01216_),
    .Q(\cpuregs[4][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50187_ (.CLK(clk_0_1312),
    .D(_01186_),
    .Q(\cpuregs[4][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50188_ (.CLK(clk_0_1312),
    .D(_01187_),
    .Q(\cpuregs[4][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50189_ (.CLK(clk_0_1312),
    .D(_01188_),
    .Q(\cpuregs[4][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50190_ (.CLK(clk_0_1312),
    .D(_01189_),
    .Q(\cpuregs[4][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50191_ (.CLK(clk_0_1312),
    .D(_01190_),
    .Q(\cpuregs[4][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50192_ (.CLK(clk_0_1312),
    .D(_01191_),
    .Q(\cpuregs[4][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50193_ (.CLK(clk_0_1312),
    .D(_01192_),
    .Q(\cpuregs[4][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50194_ (.CLK(clk_0_1312),
    .D(_01193_),
    .Q(\cpuregs[4][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50195_ (.CLK(clk_0_1312),
    .D(_01194_),
    .Q(\cpuregs[4][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50196_ (.CLK(clk_0_1312),
    .D(_01195_),
    .Q(\cpuregs[4][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50197_ (.CLK(clk_0_1312),
    .D(_01197_),
    .Q(\cpuregs[4][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50198_ (.CLK(clk_0_1328),
    .D(_01198_),
    .Q(\cpuregs[4][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50199_ (.CLK(clk_0_1328),
    .D(_01199_),
    .Q(\cpuregs[4][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50200_ (.CLK(clk_0_1328),
    .D(_01200_),
    .Q(\cpuregs[4][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50201_ (.CLK(clk_0_1328),
    .D(_01201_),
    .Q(\cpuregs[4][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50202_ (.CLK(clk_0_1328),
    .D(_01202_),
    .Q(\cpuregs[4][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50203_ (.CLK(clk_0_1328),
    .D(_01203_),
    .Q(\cpuregs[4][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50204_ (.CLK(clk_0_1328),
    .D(_01204_),
    .Q(\cpuregs[4][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50205_ (.CLK(clk_0_1328),
    .D(_01205_),
    .Q(\cpuregs[4][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50206_ (.CLK(clk_0_1328),
    .D(_01206_),
    .Q(\cpuregs[4][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50207_ (.CLK(clk_0_1328),
    .D(_01208_),
    .Q(\cpuregs[4][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50208_ (.CLK(clk_0_1328),
    .D(_01209_),
    .Q(\cpuregs[4][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50209_ (.CLK(clk_0_1328),
    .D(_00737_),
    .Q(\cpuregs[0][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50210_ (.CLK(clk_0_1328),
    .D(_00748_),
    .Q(\cpuregs[0][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50211_ (.CLK(clk_0_1328),
    .D(_00759_),
    .Q(\cpuregs[0][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50212_ (.CLK(clk_0_1328),
    .D(_00762_),
    .Q(\cpuregs[0][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50213_ (.CLK(clk_0_1328),
    .D(_00763_),
    .Q(\cpuregs[0][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50214_ (.CLK(clk_0_1344),
    .D(_00764_),
    .Q(\cpuregs[0][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50215_ (.CLK(clk_0_1344),
    .D(_00765_),
    .Q(\cpuregs[0][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50216_ (.CLK(clk_0_1344),
    .D(_00766_),
    .Q(\cpuregs[0][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50217_ (.CLK(clk_0_1344),
    .D(_00767_),
    .Q(\cpuregs[0][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50218_ (.CLK(clk_0_1344),
    .D(_00768_),
    .Q(\cpuregs[0][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50219_ (.CLK(clk_0_1344),
    .D(_00738_),
    .Q(\cpuregs[0][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50220_ (.CLK(clk_0_1344),
    .D(_00739_),
    .Q(\cpuregs[0][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50221_ (.CLK(clk_0_1344),
    .D(_00740_),
    .Q(\cpuregs[0][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50222_ (.CLK(clk_0_1344),
    .D(_00741_),
    .Q(\cpuregs[0][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50223_ (.CLK(clk_0_1344),
    .D(_00742_),
    .Q(\cpuregs[0][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50224_ (.CLK(clk_0_1344),
    .D(_00743_),
    .Q(\cpuregs[0][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50225_ (.CLK(clk_0_1344),
    .D(_00744_),
    .Q(\cpuregs[0][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50226_ (.CLK(clk_0_1344),
    .D(_00745_),
    .Q(\cpuregs[0][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50227_ (.CLK(clk_0_1344),
    .D(_00746_),
    .Q(\cpuregs[0][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50228_ (.CLK(clk_0_1344),
    .D(_00747_),
    .Q(\cpuregs[0][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50229_ (.CLK(clk_0_1344),
    .D(_00749_),
    .Q(\cpuregs[0][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50230_ (.CLK(clk_0_1360),
    .D(_00750_),
    .Q(\cpuregs[0][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50231_ (.CLK(clk_0_1360),
    .D(_00751_),
    .Q(\cpuregs[0][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50232_ (.CLK(clk_0_1360),
    .D(_00752_),
    .Q(\cpuregs[0][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50233_ (.CLK(clk_0_1360),
    .D(_00753_),
    .Q(\cpuregs[0][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50234_ (.CLK(clk_0_1360),
    .D(_00754_),
    .Q(\cpuregs[0][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50235_ (.CLK(clk_0_1360),
    .D(_00755_),
    .Q(\cpuregs[0][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50236_ (.CLK(clk_0_1360),
    .D(_00756_),
    .Q(\cpuregs[0][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50237_ (.CLK(clk_0_1360),
    .D(_00757_),
    .Q(\cpuregs[0][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50238_ (.CLK(clk_0_1360),
    .D(_00758_),
    .Q(\cpuregs[0][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50239_ (.CLK(clk_0_1360),
    .D(_00760_),
    .Q(\cpuregs[0][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50240_ (.CLK(clk_0_1360),
    .D(_00761_),
    .Q(\cpuregs[0][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50241_ (.CLK(clk_0_1360),
    .D(_01121_),
    .Q(\cpuregs[2][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50242_ (.CLK(clk_0_1360),
    .D(_01132_),
    .Q(\cpuregs[2][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50243_ (.CLK(clk_0_1360),
    .D(_01143_),
    .Q(\cpuregs[2][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50244_ (.CLK(clk_0_1360),
    .D(_01146_),
    .Q(\cpuregs[2][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50245_ (.CLK(clk_0_1360),
    .D(_01147_),
    .Q(\cpuregs[2][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50246_ (.CLK(clk_0_1376),
    .D(_01148_),
    .Q(\cpuregs[2][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50247_ (.CLK(clk_0_1376),
    .D(_01149_),
    .Q(\cpuregs[2][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50248_ (.CLK(clk_0_1376),
    .D(_01150_),
    .Q(\cpuregs[2][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50249_ (.CLK(clk_0_1376),
    .D(_01151_),
    .Q(\cpuregs[2][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50250_ (.CLK(clk_0_1376),
    .D(_01152_),
    .Q(\cpuregs[2][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50251_ (.CLK(clk_0_1376),
    .D(_01122_),
    .Q(\cpuregs[2][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50252_ (.CLK(clk_0_1376),
    .D(_01123_),
    .Q(\cpuregs[2][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50253_ (.CLK(clk_0_1376),
    .D(_01124_),
    .Q(\cpuregs[2][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50254_ (.CLK(clk_0_1376),
    .D(_01125_),
    .Q(\cpuregs[2][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50255_ (.CLK(clk_0_1376),
    .D(_01126_),
    .Q(\cpuregs[2][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50256_ (.CLK(clk_0_1376),
    .D(_01127_),
    .Q(\cpuregs[2][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50257_ (.CLK(clk_0_1376),
    .D(_01128_),
    .Q(\cpuregs[2][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50258_ (.CLK(clk_0_1376),
    .D(_01129_),
    .Q(\cpuregs[2][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50259_ (.CLK(clk_0_1376),
    .D(_01130_),
    .Q(\cpuregs[2][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50260_ (.CLK(clk_0_1376),
    .D(_01131_),
    .Q(\cpuregs[2][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50261_ (.CLK(clk_0_1376),
    .D(_01133_),
    .Q(\cpuregs[2][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50262_ (.CLK(clk_0_1392),
    .D(_01134_),
    .Q(\cpuregs[2][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50263_ (.CLK(clk_0_1392),
    .D(_01135_),
    .Q(\cpuregs[2][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50264_ (.CLK(clk_0_1392),
    .D(_01136_),
    .Q(\cpuregs[2][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50265_ (.CLK(clk_0_1392),
    .D(_01137_),
    .Q(\cpuregs[2][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50266_ (.CLK(clk_0_1392),
    .D(_01138_),
    .Q(\cpuregs[2][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50267_ (.CLK(clk_0_1392),
    .D(_01139_),
    .Q(\cpuregs[2][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50268_ (.CLK(clk_0_1392),
    .D(_01140_),
    .Q(\cpuregs[2][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50269_ (.CLK(clk_0_1392),
    .D(_01141_),
    .Q(\cpuregs[2][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50270_ (.CLK(clk_0_1392),
    .D(_01142_),
    .Q(\cpuregs[2][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50271_ (.CLK(clk_0_1392),
    .D(_01144_),
    .Q(\cpuregs[2][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50272_ (.CLK(clk_0_1392),
    .D(_01145_),
    .Q(\cpuregs[2][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50273_ (.CLK(clk_0_1392),
    .D(_01281_),
    .Q(\cpuregs[7][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50274_ (.CLK(clk_0_1392),
    .D(_01292_),
    .Q(\cpuregs[7][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50275_ (.CLK(clk_0_1392),
    .D(_01303_),
    .Q(\cpuregs[7][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50276_ (.CLK(clk_0_1392),
    .D(_01306_),
    .Q(\cpuregs[7][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50277_ (.CLK(clk_0_1392),
    .D(_01307_),
    .Q(\cpuregs[7][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50278_ (.CLK(clk_0_1408),
    .D(_01308_),
    .Q(\cpuregs[7][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50279_ (.CLK(clk_0_1408),
    .D(_01309_),
    .Q(\cpuregs[7][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50280_ (.CLK(clk_0_1408),
    .D(_01310_),
    .Q(\cpuregs[7][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50281_ (.CLK(clk_0_1408),
    .D(_01311_),
    .Q(\cpuregs[7][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50282_ (.CLK(clk_0_1408),
    .D(_01312_),
    .Q(\cpuregs[7][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50283_ (.CLK(clk_0_1408),
    .D(_01282_),
    .Q(\cpuregs[7][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50284_ (.CLK(clk_0_1408),
    .D(_01283_),
    .Q(\cpuregs[7][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50285_ (.CLK(clk_0_1408),
    .D(_01284_),
    .Q(\cpuregs[7][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50286_ (.CLK(clk_0_1408),
    .D(_01285_),
    .Q(\cpuregs[7][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50287_ (.CLK(clk_0_1408),
    .D(_01286_),
    .Q(\cpuregs[7][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50288_ (.CLK(clk_0_1408),
    .D(_01287_),
    .Q(\cpuregs[7][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50289_ (.CLK(clk_0_1408),
    .D(_01288_),
    .Q(\cpuregs[7][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50290_ (.CLK(clk_0_1408),
    .D(_01289_),
    .Q(\cpuregs[7][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50291_ (.CLK(clk_0_1408),
    .D(_01290_),
    .Q(\cpuregs[7][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50292_ (.CLK(clk_0_1408),
    .D(_01291_),
    .Q(\cpuregs[7][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50293_ (.CLK(clk_0_1408),
    .D(_01293_),
    .Q(\cpuregs[7][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50294_ (.CLK(clk_0_1424),
    .D(_01294_),
    .Q(\cpuregs[7][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50295_ (.CLK(clk_0_1424),
    .D(_01295_),
    .Q(\cpuregs[7][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50296_ (.CLK(clk_0_1424),
    .D(_01296_),
    .Q(\cpuregs[7][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50297_ (.CLK(clk_0_1424),
    .D(_01297_),
    .Q(\cpuregs[7][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50298_ (.CLK(clk_0_1424),
    .D(_01298_),
    .Q(\cpuregs[7][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50299_ (.CLK(clk_0_1424),
    .D(_01299_),
    .Q(\cpuregs[7][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50300_ (.CLK(clk_0_1424),
    .D(_01300_),
    .Q(\cpuregs[7][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50301_ (.CLK(clk_0_1424),
    .D(_01301_),
    .Q(\cpuregs[7][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50302_ (.CLK(clk_0_1424),
    .D(_01302_),
    .Q(\cpuregs[7][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50303_ (.CLK(clk_0_1424),
    .D(_01304_),
    .Q(\cpuregs[7][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50304_ (.CLK(clk_0_1424),
    .D(_01305_),
    .Q(\cpuregs[7][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50305_ (.CLK(clk_0_1424),
    .D(_00659_),
    .Q(\cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _50306_ (.CLK(clk_0_1424),
    .D(_00660_),
    .Q(\cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _50307_ (.CLK(clk_0_1424),
    .D(_00661_),
    .Q(\cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _50308_ (.CLK(clk_0_1424),
    .D(_00662_),
    .Q(\cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_4 _50309_ (.CLK(clk_0_1424),
    .D(_00663_),
    .Q(\cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_4 _50310_ (.CLK(clk_0_1440),
    .D(_00664_),
    .Q(\cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_4 _50311_ (.CLK(clk_0_1440),
    .D(_00665_),
    .Q(\cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_4 _50312_ (.CLK(clk_0_1440),
    .D(_01249_),
    .Q(\cpuregs[6][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50313_ (.CLK(clk_0_1440),
    .D(_01260_),
    .Q(\cpuregs[6][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50314_ (.CLK(clk_0_1440),
    .D(_01271_),
    .Q(\cpuregs[6][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50315_ (.CLK(clk_0_1440),
    .D(_01274_),
    .Q(\cpuregs[6][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50316_ (.CLK(clk_0_1440),
    .D(_01275_),
    .Q(\cpuregs[6][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50317_ (.CLK(clk_0_1440),
    .D(_01276_),
    .Q(\cpuregs[6][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50318_ (.CLK(clk_0_1440),
    .D(_01277_),
    .Q(\cpuregs[6][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50319_ (.CLK(clk_0_1440),
    .D(_01278_),
    .Q(\cpuregs[6][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50320_ (.CLK(clk_0_1440),
    .D(_01279_),
    .Q(\cpuregs[6][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50321_ (.CLK(clk_0_1440),
    .D(_01280_),
    .Q(\cpuregs[6][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50322_ (.CLK(clk_0_1440),
    .D(_01250_),
    .Q(\cpuregs[6][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50323_ (.CLK(clk_0_1440),
    .D(_01251_),
    .Q(\cpuregs[6][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50324_ (.CLK(clk_0_1440),
    .D(_01252_),
    .Q(\cpuregs[6][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50325_ (.CLK(clk_0_1440),
    .D(_01253_),
    .Q(\cpuregs[6][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50326_ (.CLK(clk_0_1456),
    .D(_01254_),
    .Q(\cpuregs[6][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50327_ (.CLK(clk_0_1456),
    .D(_01255_),
    .Q(\cpuregs[6][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50328_ (.CLK(clk_0_1456),
    .D(_01256_),
    .Q(\cpuregs[6][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50329_ (.CLK(clk_0_1456),
    .D(_01257_),
    .Q(\cpuregs[6][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50330_ (.CLK(clk_0_1456),
    .D(_01258_),
    .Q(\cpuregs[6][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50331_ (.CLK(clk_0_1456),
    .D(_01259_),
    .Q(\cpuregs[6][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50332_ (.CLK(clk_0_1456),
    .D(_01261_),
    .Q(\cpuregs[6][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50333_ (.CLK(clk_0_1456),
    .D(_01262_),
    .Q(\cpuregs[6][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50334_ (.CLK(clk_0_1456),
    .D(_01263_),
    .Q(\cpuregs[6][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50335_ (.CLK(clk_0_1456),
    .D(_01264_),
    .Q(\cpuregs[6][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50336_ (.CLK(clk_0_1456),
    .D(_01265_),
    .Q(\cpuregs[6][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50337_ (.CLK(clk_0_1456),
    .D(_01266_),
    .Q(\cpuregs[6][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50338_ (.CLK(clk_0_1456),
    .D(_01267_),
    .Q(\cpuregs[6][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50339_ (.CLK(clk_0_1456),
    .D(_01268_),
    .Q(\cpuregs[6][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50340_ (.CLK(clk_0_1456),
    .D(_01269_),
    .Q(\cpuregs[6][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50341_ (.CLK(clk_0_1456),
    .D(_01270_),
    .Q(\cpuregs[6][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50342_ (.CLK(clk_0_1472),
    .D(_01272_),
    .Q(\cpuregs[6][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50343_ (.CLK(clk_0_1472),
    .D(_01273_),
    .Q(\cpuregs[6][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50344_ (.CLK(clk_0_1472),
    .D(_00801_),
    .Q(\cpuregs[11][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50345_ (.CLK(clk_0_1472),
    .D(_00812_),
    .Q(\cpuregs[11][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50346_ (.CLK(clk_0_1472),
    .D(_00823_),
    .Q(\cpuregs[11][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50347_ (.CLK(clk_0_1472),
    .D(_00826_),
    .Q(\cpuregs[11][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50348_ (.CLK(clk_0_1472),
    .D(_00827_),
    .Q(\cpuregs[11][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50349_ (.CLK(clk_0_1472),
    .D(_00828_),
    .Q(\cpuregs[11][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50350_ (.CLK(clk_0_1472),
    .D(_00829_),
    .Q(\cpuregs[11][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50351_ (.CLK(clk_0_1472),
    .D(_00830_),
    .Q(\cpuregs[11][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50352_ (.CLK(clk_0_1472),
    .D(_00831_),
    .Q(\cpuregs[11][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50353_ (.CLK(clk_0_1472),
    .D(_00832_),
    .Q(\cpuregs[11][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50354_ (.CLK(clk_0_1472),
    .D(_00802_),
    .Q(\cpuregs[11][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50355_ (.CLK(clk_0_1472),
    .D(_00803_),
    .Q(\cpuregs[11][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50356_ (.CLK(clk_0_1472),
    .D(_00804_),
    .Q(\cpuregs[11][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50357_ (.CLK(clk_0_1472),
    .D(_00805_),
    .Q(\cpuregs[11][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50358_ (.CLK(clk_0_1488),
    .D(_00806_),
    .Q(\cpuregs[11][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50359_ (.CLK(clk_0_1488),
    .D(_00807_),
    .Q(\cpuregs[11][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50360_ (.CLK(clk_0_1488),
    .D(_00808_),
    .Q(\cpuregs[11][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50361_ (.CLK(clk_0_1488),
    .D(_00809_),
    .Q(\cpuregs[11][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50362_ (.CLK(clk_0_1488),
    .D(_00810_),
    .Q(\cpuregs[11][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50363_ (.CLK(clk_0_1488),
    .D(_00811_),
    .Q(\cpuregs[11][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50364_ (.CLK(clk_0_1488),
    .D(_00813_),
    .Q(\cpuregs[11][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50365_ (.CLK(clk_0_1488),
    .D(_00814_),
    .Q(\cpuregs[11][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50366_ (.CLK(clk_0_1488),
    .D(_00815_),
    .Q(\cpuregs[11][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50367_ (.CLK(clk_0_1488),
    .D(_00816_),
    .Q(\cpuregs[11][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50368_ (.CLK(clk_0_1488),
    .D(_00817_),
    .Q(\cpuregs[11][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50369_ (.CLK(clk_0_1488),
    .D(_00818_),
    .Q(\cpuregs[11][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50370_ (.CLK(clk_0_1488),
    .D(_00819_),
    .Q(\cpuregs[11][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50371_ (.CLK(clk_0_1488),
    .D(_00820_),
    .Q(\cpuregs[11][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50372_ (.CLK(clk_0_1488),
    .D(_00821_),
    .Q(\cpuregs[11][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50373_ (.CLK(clk_0_1488),
    .D(_00822_),
    .Q(\cpuregs[11][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50374_ (.CLK(clk_0_1504),
    .D(_00824_),
    .Q(\cpuregs[11][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50375_ (.CLK(clk_0_1504),
    .D(_00825_),
    .Q(\cpuregs[11][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50376_ (.CLK(clk_0_1504),
    .D(_01217_),
    .Q(\cpuregs[5][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50377_ (.CLK(clk_0_1504),
    .D(_01228_),
    .Q(\cpuregs[5][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50378_ (.CLK(clk_0_1504),
    .D(_01239_),
    .Q(\cpuregs[5][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50379_ (.CLK(clk_0_1504),
    .D(_01242_),
    .Q(\cpuregs[5][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50380_ (.CLK(clk_0_1504),
    .D(_01243_),
    .Q(\cpuregs[5][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50381_ (.CLK(clk_0_1504),
    .D(_01244_),
    .Q(\cpuregs[5][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50382_ (.CLK(clk_0_1504),
    .D(_01245_),
    .Q(\cpuregs[5][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50383_ (.CLK(clk_0_1504),
    .D(_01246_),
    .Q(\cpuregs[5][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50384_ (.CLK(clk_0_1504),
    .D(_01247_),
    .Q(\cpuregs[5][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50385_ (.CLK(clk_0_1504),
    .D(_01248_),
    .Q(\cpuregs[5][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50386_ (.CLK(clk_0_1504),
    .D(_01218_),
    .Q(\cpuregs[5][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50387_ (.CLK(clk_0_1504),
    .D(_01219_),
    .Q(\cpuregs[5][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50388_ (.CLK(clk_0_1504),
    .D(_01220_),
    .Q(\cpuregs[5][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50389_ (.CLK(clk_0_1504),
    .D(_01221_),
    .Q(\cpuregs[5][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50390_ (.CLK(clk_0_1520),
    .D(_01222_),
    .Q(\cpuregs[5][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50391_ (.CLK(clk_0_1520),
    .D(_01223_),
    .Q(\cpuregs[5][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50392_ (.CLK(clk_0_1520),
    .D(_01224_),
    .Q(\cpuregs[5][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50393_ (.CLK(clk_0_1520),
    .D(_01225_),
    .Q(\cpuregs[5][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50394_ (.CLK(clk_0_1520),
    .D(_01226_),
    .Q(\cpuregs[5][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50395_ (.CLK(clk_0_1520),
    .D(_01227_),
    .Q(\cpuregs[5][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50396_ (.CLK(clk_0_1520),
    .D(_01229_),
    .Q(\cpuregs[5][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50397_ (.CLK(clk_0_1520),
    .D(_01230_),
    .Q(\cpuregs[5][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50398_ (.CLK(clk_0_1520),
    .D(_01231_),
    .Q(\cpuregs[5][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50399_ (.CLK(clk_0_1520),
    .D(_01232_),
    .Q(\cpuregs[5][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50400_ (.CLK(clk_0_1520),
    .D(_01233_),
    .Q(\cpuregs[5][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50401_ (.CLK(clk_0_1520),
    .D(_01234_),
    .Q(\cpuregs[5][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50402_ (.CLK(clk_0_1520),
    .D(_01235_),
    .Q(\cpuregs[5][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50403_ (.CLK(clk_0_1520),
    .D(_01236_),
    .Q(\cpuregs[5][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50404_ (.CLK(clk_0_1520),
    .D(_01237_),
    .Q(\cpuregs[5][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50405_ (.CLK(clk_0_1520),
    .D(_01238_),
    .Q(\cpuregs[5][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50406_ (.CLK(clk_0_1536),
    .D(_01240_),
    .Q(\cpuregs[5][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50407_ (.CLK(clk_0_1536),
    .D(_01241_),
    .Q(\cpuregs[5][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50408_ (.CLK(clk_0_1536),
    .D(_01089_),
    .Q(\cpuregs[1][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50409_ (.CLK(clk_0_1536),
    .D(_01100_),
    .Q(\cpuregs[1][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50410_ (.CLK(clk_0_1536),
    .D(_01111_),
    .Q(\cpuregs[1][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50411_ (.CLK(clk_0_1536),
    .D(_01114_),
    .Q(\cpuregs[1][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50412_ (.CLK(clk_0_1536),
    .D(_01115_),
    .Q(\cpuregs[1][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50413_ (.CLK(clk_0_1536),
    .D(_01116_),
    .Q(\cpuregs[1][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50414_ (.CLK(clk_0_1536),
    .D(_01117_),
    .Q(\cpuregs[1][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50415_ (.CLK(clk_0_1536),
    .D(_01118_),
    .Q(\cpuregs[1][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50416_ (.CLK(clk_0_1536),
    .D(_01119_),
    .Q(\cpuregs[1][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50417_ (.CLK(clk_0_1536),
    .D(_01120_),
    .Q(\cpuregs[1][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50418_ (.CLK(clk_0_1536),
    .D(_01090_),
    .Q(\cpuregs[1][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50419_ (.CLK(clk_0_1536),
    .D(_01091_),
    .Q(\cpuregs[1][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50420_ (.CLK(clk_0_1536),
    .D(_01092_),
    .Q(\cpuregs[1][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50421_ (.CLK(clk_0_1536),
    .D(_01093_),
    .Q(\cpuregs[1][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50422_ (.CLK(clk_0_1552),
    .D(_01094_),
    .Q(\cpuregs[1][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50423_ (.CLK(clk_0_1552),
    .D(_01095_),
    .Q(\cpuregs[1][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50424_ (.CLK(clk_0_1552),
    .D(_01096_),
    .Q(\cpuregs[1][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50425_ (.CLK(clk_0_1552),
    .D(_01097_),
    .Q(\cpuregs[1][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50426_ (.CLK(clk_0_1552),
    .D(_01098_),
    .Q(\cpuregs[1][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50427_ (.CLK(clk_0_1552),
    .D(_01099_),
    .Q(\cpuregs[1][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50428_ (.CLK(clk_0_1552),
    .D(_01101_),
    .Q(\cpuregs[1][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50429_ (.CLK(clk_0_1552),
    .D(_01102_),
    .Q(\cpuregs[1][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50430_ (.CLK(clk_0_1552),
    .D(_01103_),
    .Q(\cpuregs[1][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50431_ (.CLK(clk_0_1552),
    .D(_01104_),
    .Q(\cpuregs[1][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50432_ (.CLK(clk_0_1552),
    .D(_01105_),
    .Q(\cpuregs[1][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50433_ (.CLK(clk_0_1552),
    .D(_01106_),
    .Q(\cpuregs[1][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50434_ (.CLK(clk_0_1552),
    .D(_01107_),
    .Q(\cpuregs[1][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50435_ (.CLK(clk_0_1552),
    .D(_01108_),
    .Q(\cpuregs[1][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50436_ (.CLK(clk_0_1552),
    .D(_01109_),
    .Q(\cpuregs[1][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50437_ (.CLK(clk_0_1552),
    .D(_01110_),
    .Q(\cpuregs[1][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50438_ (.CLK(clk_0_1568),
    .D(_01112_),
    .Q(\cpuregs[1][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50439_ (.CLK(clk_0_1568),
    .D(_01113_),
    .Q(\cpuregs[1][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50440_ (.CLK(clk_0_1568),
    .D(_00961_),
    .Q(\cpuregs[16][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50441_ (.CLK(clk_0_1568),
    .D(_00972_),
    .Q(\cpuregs[16][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50442_ (.CLK(clk_0_1568),
    .D(_00983_),
    .Q(\cpuregs[16][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50443_ (.CLK(clk_0_1568),
    .D(_00986_),
    .Q(\cpuregs[16][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50444_ (.CLK(clk_0_1568),
    .D(_00987_),
    .Q(\cpuregs[16][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50445_ (.CLK(clk_0_1568),
    .D(_00988_),
    .Q(\cpuregs[16][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50446_ (.CLK(clk_0_1568),
    .D(_00989_),
    .Q(\cpuregs[16][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50447_ (.CLK(clk_0_1568),
    .D(_00990_),
    .Q(\cpuregs[16][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50448_ (.CLK(clk_0_1568),
    .D(_00991_),
    .Q(\cpuregs[16][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50449_ (.CLK(clk_0_1568),
    .D(_00992_),
    .Q(\cpuregs[16][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50450_ (.CLK(clk_0_1568),
    .D(_00962_),
    .Q(\cpuregs[16][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50451_ (.CLK(clk_0_1568),
    .D(_00963_),
    .Q(\cpuregs[16][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50452_ (.CLK(clk_0_1568),
    .D(_00964_),
    .Q(\cpuregs[16][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50453_ (.CLK(clk_0_1568),
    .D(_00965_),
    .Q(\cpuregs[16][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50454_ (.CLK(clk_0_1584),
    .D(_00966_),
    .Q(\cpuregs[16][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50455_ (.CLK(clk_0_1584),
    .D(_00967_),
    .Q(\cpuregs[16][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50456_ (.CLK(clk_0_1584),
    .D(_00968_),
    .Q(\cpuregs[16][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50457_ (.CLK(clk_0_1584),
    .D(_00969_),
    .Q(\cpuregs[16][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50458_ (.CLK(clk_0_1584),
    .D(_00970_),
    .Q(\cpuregs[16][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50459_ (.CLK(clk_0_1584),
    .D(_00971_),
    .Q(\cpuregs[16][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50460_ (.CLK(clk_0_1584),
    .D(_00973_),
    .Q(\cpuregs[16][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50461_ (.CLK(clk_0_1584),
    .D(_00974_),
    .Q(\cpuregs[16][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50462_ (.CLK(clk_0_1584),
    .D(_00975_),
    .Q(\cpuregs[16][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50463_ (.CLK(clk_0_1584),
    .D(_00976_),
    .Q(\cpuregs[16][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50464_ (.CLK(clk_0_1584),
    .D(_00977_),
    .Q(\cpuregs[16][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50465_ (.CLK(clk_0_1584),
    .D(_00978_),
    .Q(\cpuregs[16][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50466_ (.CLK(clk_0_1584),
    .D(_00979_),
    .Q(\cpuregs[16][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50467_ (.CLK(clk_0_1584),
    .D(_00980_),
    .Q(\cpuregs[16][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50468_ (.CLK(clk_0_1584),
    .D(_00981_),
    .Q(\cpuregs[16][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50469_ (.CLK(clk_0_1584),
    .D(_00982_),
    .Q(\cpuregs[16][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50470_ (.CLK(clk_0_1600),
    .D(_00984_),
    .Q(\cpuregs[16][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50471_ (.CLK(clk_0_1600),
    .D(_00985_),
    .Q(\cpuregs[16][31] ));
 sky130_fd_sc_hd__dfxtp_4 _50472_ (.CLK(clk_0_1600),
    .D(_01313_),
    .Q(\cpuregs[8][0] ));
 sky130_fd_sc_hd__dfxtp_4 _50473_ (.CLK(clk_0_1600),
    .D(_01324_),
    .Q(\cpuregs[8][1] ));
 sky130_fd_sc_hd__dfxtp_4 _50474_ (.CLK(clk_0_1600),
    .D(_01335_),
    .Q(\cpuregs[8][2] ));
 sky130_fd_sc_hd__dfxtp_4 _50475_ (.CLK(clk_0_1600),
    .D(_01338_),
    .Q(\cpuregs[8][3] ));
 sky130_fd_sc_hd__dfxtp_4 _50476_ (.CLK(clk_0_1600),
    .D(_01339_),
    .Q(\cpuregs[8][4] ));
 sky130_fd_sc_hd__dfxtp_4 _50477_ (.CLK(clk_0_1600),
    .D(_01340_),
    .Q(\cpuregs[8][5] ));
 sky130_fd_sc_hd__dfxtp_4 _50478_ (.CLK(clk_0_1600),
    .D(_01341_),
    .Q(\cpuregs[8][6] ));
 sky130_fd_sc_hd__dfxtp_4 _50479_ (.CLK(clk_0_1600),
    .D(_01342_),
    .Q(\cpuregs[8][7] ));
 sky130_fd_sc_hd__dfxtp_4 _50480_ (.CLK(clk_0_1600),
    .D(_01343_),
    .Q(\cpuregs[8][8] ));
 sky130_fd_sc_hd__dfxtp_4 _50481_ (.CLK(clk_0_1600),
    .D(_01344_),
    .Q(\cpuregs[8][9] ));
 sky130_fd_sc_hd__dfxtp_4 _50482_ (.CLK(clk_0_1600),
    .D(_01314_),
    .Q(\cpuregs[8][10] ));
 sky130_fd_sc_hd__dfxtp_4 _50483_ (.CLK(clk_0_1600),
    .D(_01315_),
    .Q(\cpuregs[8][11] ));
 sky130_fd_sc_hd__dfxtp_4 _50484_ (.CLK(clk_0_1600),
    .D(_01316_),
    .Q(\cpuregs[8][12] ));
 sky130_fd_sc_hd__dfxtp_4 _50485_ (.CLK(clk_0_1600),
    .D(_01317_),
    .Q(\cpuregs[8][13] ));
 sky130_fd_sc_hd__dfxtp_4 _50486_ (.CLK(clk_0_1616),
    .D(_01318_),
    .Q(\cpuregs[8][14] ));
 sky130_fd_sc_hd__dfxtp_4 _50487_ (.CLK(clk_0_1616),
    .D(_01319_),
    .Q(\cpuregs[8][15] ));
 sky130_fd_sc_hd__dfxtp_4 _50488_ (.CLK(clk_0_1616),
    .D(_01320_),
    .Q(\cpuregs[8][16] ));
 sky130_fd_sc_hd__dfxtp_4 _50489_ (.CLK(clk_0_1616),
    .D(_01321_),
    .Q(\cpuregs[8][17] ));
 sky130_fd_sc_hd__dfxtp_4 _50490_ (.CLK(clk_0_1616),
    .D(_01322_),
    .Q(\cpuregs[8][18] ));
 sky130_fd_sc_hd__dfxtp_4 _50491_ (.CLK(clk_0_1616),
    .D(_01323_),
    .Q(\cpuregs[8][19] ));
 sky130_fd_sc_hd__dfxtp_4 _50492_ (.CLK(clk_0_1616),
    .D(_01325_),
    .Q(\cpuregs[8][20] ));
 sky130_fd_sc_hd__dfxtp_4 _50493_ (.CLK(clk_0_1616),
    .D(_01326_),
    .Q(\cpuregs[8][21] ));
 sky130_fd_sc_hd__dfxtp_4 _50494_ (.CLK(clk_0_1616),
    .D(_01327_),
    .Q(\cpuregs[8][22] ));
 sky130_fd_sc_hd__dfxtp_4 _50495_ (.CLK(clk_0_1616),
    .D(_01328_),
    .Q(\cpuregs[8][23] ));
 sky130_fd_sc_hd__dfxtp_4 _50496_ (.CLK(clk_0_1616),
    .D(_01329_),
    .Q(\cpuregs[8][24] ));
 sky130_fd_sc_hd__dfxtp_4 _50497_ (.CLK(clk_0_1616),
    .D(_01330_),
    .Q(\cpuregs[8][25] ));
 sky130_fd_sc_hd__dfxtp_4 _50498_ (.CLK(clk_0_1616),
    .D(_01331_),
    .Q(\cpuregs[8][26] ));
 sky130_fd_sc_hd__dfxtp_4 _50499_ (.CLK(clk_0_1616),
    .D(_01332_),
    .Q(\cpuregs[8][27] ));
 sky130_fd_sc_hd__dfxtp_4 _50500_ (.CLK(clk_0_1616),
    .D(_01333_),
    .Q(\cpuregs[8][28] ));
 sky130_fd_sc_hd__dfxtp_4 _50501_ (.CLK(clk_0_1616),
    .D(_01334_),
    .Q(\cpuregs[8][29] ));
 sky130_fd_sc_hd__dfxtp_4 _50502_ (.CLK(clk_0_1632),
    .D(_01336_),
    .Q(\cpuregs[8][30] ));
 sky130_fd_sc_hd__dfxtp_4 _50503_ (.CLK(clk_0_1632),
    .D(_01337_),
    .Q(\cpuregs[8][31] ));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_0 (.A(clk_1_0),
    .X(clk_0_0));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1008 (.A(clk_1_768),
    .X(clk_0_1008));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1024 (.A(clk_1_1024),
    .X(clk_0_1024));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1040 (.A(clk_1_1024),
    .X(clk_0_1040));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1056 (.A(clk_1_1024),
    .X(clk_0_1056));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1072 (.A(clk_1_1024),
    .X(clk_0_1072));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1088 (.A(clk_1_1024),
    .X(clk_0_1088));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1104 (.A(clk_1_1024),
    .X(clk_0_1104));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_112 (.A(clk_1_0),
    .X(clk_0_112));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1120 (.A(clk_1_1024),
    .X(clk_0_1120));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1136 (.A(clk_1_1024),
    .X(clk_0_1136));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1152 (.A(clk_1_1024),
    .X(clk_0_1152));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1168 (.A(clk_1_1024),
    .X(clk_0_1168));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1184 (.A(clk_1_1024),
    .X(clk_0_1184));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1200 (.A(clk_1_1024),
    .X(clk_0_1200));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1216 (.A(clk_1_1024),
    .X(clk_0_1216));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1232 (.A(clk_1_1024),
    .X(clk_0_1232));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1248 (.A(clk_1_1024),
    .X(clk_0_1248));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1264 (.A(clk_1_1024),
    .X(clk_0_1264));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_128 (.A(clk_1_0),
    .X(clk_0_128));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1280 (.A(clk_1_1280),
    .X(clk_0_1280));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1296 (.A(clk_1_1280),
    .X(clk_0_1296));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1312 (.A(clk_1_1280),
    .X(clk_0_1312));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1328 (.A(clk_1_1280),
    .X(clk_0_1328));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1344 (.A(clk_1_1280),
    .X(clk_0_1344));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1360 (.A(clk_1_1280),
    .X(clk_0_1360));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1376 (.A(clk_1_1280),
    .X(clk_0_1376));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1392 (.A(clk_1_1280),
    .X(clk_0_1392));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1408 (.A(clk_1_1280),
    .X(clk_0_1408));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1424 (.A(clk_1_1280),
    .X(clk_0_1424));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_144 (.A(clk_1_0),
    .X(clk_0_144));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1440 (.A(clk_1_1280),
    .X(clk_0_1440));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1456 (.A(clk_1_1280),
    .X(clk_0_1456));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1472 (.A(clk_1_1280),
    .X(clk_0_1472));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1488 (.A(clk_1_1280),
    .X(clk_0_1488));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1504 (.A(clk_1_1280),
    .X(clk_0_1504));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1520 (.A(clk_1_1280),
    .X(clk_0_1520));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1536 (.A(clk_1_1536),
    .X(clk_0_1536));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1552 (.A(clk_1_1536),
    .X(clk_0_1552));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1568 (.A(clk_1_1536),
    .X(clk_0_1568));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1584 (.A(clk_1_1536),
    .X(clk_0_1584));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_16 (.A(clk_1_0),
    .X(clk_0_16));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_160 (.A(clk_1_0),
    .X(clk_0_160));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1600 (.A(clk_1_1536),
    .X(clk_0_1600));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1616 (.A(clk_1_1536),
    .X(clk_0_1616));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_1632 (.A(clk_1_1536),
    .X(clk_0_1632));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_176 (.A(clk_1_0),
    .X(clk_0_176));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_192 (.A(clk_1_0),
    .X(clk_0_192));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_208 (.A(clk_1_0),
    .X(clk_0_208));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_224 (.A(clk_1_0),
    .X(clk_0_224));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_240 (.A(clk_1_0),
    .X(clk_0_240));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_256 (.A(clk_1_256),
    .X(clk_0_256));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_272 (.A(clk_1_256),
    .X(clk_0_272));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_288 (.A(clk_1_256),
    .X(clk_0_288));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_304 (.A(clk_1_256),
    .X(clk_0_304));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_32 (.A(clk_1_0),
    .X(clk_0_32));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_320 (.A(clk_1_256),
    .X(clk_0_320));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_336 (.A(clk_1_256),
    .X(clk_0_336));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_352 (.A(clk_1_256),
    .X(clk_0_352));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_368 (.A(clk_1_256),
    .X(clk_0_368));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_384 (.A(clk_1_256),
    .X(clk_0_384));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_400 (.A(clk_1_256),
    .X(clk_0_400));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_416 (.A(clk_1_256),
    .X(clk_0_416));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_432 (.A(clk_1_256),
    .X(clk_0_432));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_448 (.A(clk_1_256),
    .X(clk_0_448));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_464 (.A(clk_1_256),
    .X(clk_0_464));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_48 (.A(clk_1_0),
    .X(clk_0_48));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_480 (.A(clk_1_256),
    .X(clk_0_480));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_496 (.A(clk_1_256),
    .X(clk_0_496));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_512 (.A(clk_1_512),
    .X(clk_0_512));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_528 (.A(clk_1_512),
    .X(clk_0_528));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_544 (.A(clk_1_512),
    .X(clk_0_544));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_560 (.A(clk_1_512),
    .X(clk_0_560));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_576 (.A(clk_1_512),
    .X(clk_0_576));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_592 (.A(clk_1_512),
    .X(clk_0_592));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_608 (.A(clk_1_512),
    .X(clk_0_608));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_624 (.A(clk_1_512),
    .X(clk_0_624));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_64 (.A(clk_1_0),
    .X(clk_0_64));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_640 (.A(clk_1_512),
    .X(clk_0_640));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_656 (.A(clk_1_512),
    .X(clk_0_656));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_672 (.A(clk_1_512),
    .X(clk_0_672));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_688 (.A(clk_1_512),
    .X(clk_0_688));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_704 (.A(clk_1_512),
    .X(clk_0_704));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_720 (.A(clk_1_512),
    .X(clk_0_720));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_736 (.A(clk_1_512),
    .X(clk_0_736));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_752 (.A(clk_1_512),
    .X(clk_0_752));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_768 (.A(clk_1_768),
    .X(clk_0_768));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_784 (.A(clk_1_768),
    .X(clk_0_784));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_80 (.A(clk_1_0),
    .X(clk_0_80));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_800 (.A(clk_1_768),
    .X(clk_0_800));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_816 (.A(clk_1_768),
    .X(clk_0_816));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_832 (.A(clk_1_768),
    .X(clk_0_832));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_848 (.A(clk_1_768),
    .X(clk_0_848));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_864 (.A(clk_1_768),
    .X(clk_0_864));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_880 (.A(clk_1_768),
    .X(clk_0_880));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_896 (.A(clk_1_768),
    .X(clk_0_896));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_912 (.A(clk_1_768),
    .X(clk_0_912));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_928 (.A(clk_1_768),
    .X(clk_0_928));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_944 (.A(clk_1_768),
    .X(clk_0_944));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_96 (.A(clk_1_0),
    .X(clk_0_96));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_960 (.A(clk_1_768),
    .X(clk_0_960));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_976 (.A(clk_1_768),
    .X(clk_0_976));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_992 (.A(clk_1_768),
    .X(clk_0_992));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_2_0 (.A(clk_2_0),
    .X(clk_1_0));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_2_1024 (.A(clk_2_0),
    .X(clk_1_1024));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_2_1280 (.A(clk_2_0),
    .X(clk_1_1280));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_2_1536 (.A(clk_2_0),
    .X(clk_1_1536));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_2_256 (.A(clk_2_0),
    .X(clk_1_256));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_2_512 (.A(clk_2_0),
    .X(clk_1_512));
 sky130_fd_sc_hd__clkbuf_4 _CTS_buf_2_768 (.A(clk_2_0),
    .X(clk_1_768));
 sky130_fd_sc_hd__clkbuf_16 _CTS_root (.A(clk),
    .X(clk_2_0));
endmodule
