magic
tech sky130A
timestamp 1614977522
<< nwell >>
rect -121 24 289 116
<< nmos >>
rect -67 -170 -44 -126
rect 5 -170 25 -126
rect 70 -170 95 -126
rect 117 -170 139 -126
rect 211 -170 231 -126
<< pmos >>
rect -60 56 -40 87
rect 5 56 25 87
rect 70 56 95 87
rect 142 56 165 87
rect 211 56 231 87
<< ndiff >>
rect -95 -133 -67 -126
rect -95 -154 -90 -133
rect -73 -154 -67 -133
rect -95 -170 -67 -154
rect -44 -170 5 -126
rect 25 -170 70 -126
rect 95 -170 117 -126
rect 139 -139 211 -126
rect 139 -160 165 -139
rect 183 -160 211 -139
rect 139 -170 211 -160
rect 231 -141 270 -126
rect 231 -162 245 -141
rect 263 -162 270 -141
rect 231 -170 270 -162
<< pdiff >>
rect 240 87 268 89
rect -97 81 -60 87
rect -97 61 -91 81
rect -74 61 -60 81
rect -97 56 -60 61
rect -40 82 5 87
rect -40 62 -25 82
rect -8 62 5 82
rect -40 56 5 62
rect 25 81 70 87
rect 25 61 39 81
rect 56 61 70 81
rect 25 56 70 61
rect 95 80 142 87
rect 95 60 110 80
rect 127 60 142 80
rect 95 56 142 60
rect 165 80 211 87
rect 165 60 179 80
rect 196 60 211 80
rect 165 56 211 60
rect 231 81 268 87
rect 231 59 245 81
rect 262 59 268 81
rect 231 56 268 59
rect -97 55 -68 56
rect 240 53 268 56
<< ndiffc >>
rect -90 -154 -73 -133
rect 165 -160 183 -139
rect 245 -162 263 -141
<< pdiffc >>
rect -91 61 -74 81
rect -25 62 -8 82
rect 39 61 56 81
rect 110 60 127 80
rect 179 60 196 80
rect 245 59 262 81
<< poly >>
rect -60 87 -40 114
rect 5 87 25 113
rect 70 87 95 115
rect 142 87 165 116
rect 211 87 231 100
rect -60 30 -40 56
rect -90 6 -40 30
rect -90 -20 -70 6
rect 5 -19 25 56
rect 70 -19 95 56
rect 142 -7 165 56
rect 118 -13 165 -7
rect -95 -25 -65 -20
rect -95 -50 -90 -25
rect -70 -50 -65 -25
rect -95 -55 -65 -50
rect 3 -27 35 -19
rect 3 -52 9 -27
rect 29 -52 35 -27
rect -90 -95 -70 -55
rect 3 -60 35 -52
rect 67 -28 97 -19
rect 67 -53 72 -28
rect 92 -53 97 -28
rect 67 -60 97 -53
rect 118 -20 170 -13
rect 118 -45 145 -20
rect 165 -45 170 -20
rect 118 -53 170 -45
rect -90 -115 -44 -95
rect -67 -126 -44 -115
rect 5 -126 25 -60
rect 70 -126 95 -60
rect 118 -81 139 -53
rect 211 -69 231 56
rect 117 -126 139 -81
rect 194 -77 231 -69
rect 194 -98 202 -77
rect 219 -98 231 -77
rect 194 -106 231 -98
rect 211 -126 231 -106
rect -67 -189 -44 -170
rect 5 -189 25 -170
rect 70 -192 95 -170
rect 117 -191 139 -170
rect 211 -203 231 -170
<< polycont >>
rect -90 -50 -70 -25
rect 9 -52 29 -27
rect 72 -53 92 -28
rect 145 -45 165 -20
rect 202 -98 219 -77
<< locali >>
rect -94 121 275 158
rect -93 87 -70 121
rect -99 81 -66 87
rect -99 61 -91 81
rect -74 61 -66 81
rect -99 56 -66 61
rect -33 82 0 91
rect 35 87 60 121
rect -33 62 -25 82
rect -8 62 0 82
rect -33 56 0 62
rect 31 81 64 87
rect 31 61 39 81
rect 56 61 64 81
rect -99 53 -68 56
rect -30 39 -5 56
rect 31 53 64 61
rect 105 80 131 88
rect 175 85 200 121
rect 105 60 110 80
rect 127 60 131 80
rect -40 35 -5 39
rect 105 35 131 60
rect 171 80 204 85
rect 171 60 179 80
rect 196 60 204 80
rect 171 52 204 60
rect 240 81 266 89
rect 240 59 245 81
rect 262 59 266 81
rect -40 15 131 35
rect -40 5 130 15
rect -98 -25 -62 -17
rect -98 -50 -90 -25
rect -70 -50 -62 -25
rect -98 -58 -62 -50
rect -40 -81 -15 5
rect 2 -27 38 -19
rect 2 -52 9 -27
rect 29 -52 38 -27
rect 2 -60 38 -52
rect 63 -28 100 -19
rect 63 -53 72 -28
rect 92 -53 100 -28
rect 63 -60 100 -53
rect 135 -20 173 -12
rect 135 -45 145 -20
rect 165 -45 173 -20
rect 240 -40 266 59
rect 135 -54 173 -45
rect 194 -77 228 -69
rect 194 -81 202 -77
rect -40 -98 202 -81
rect 219 -98 228 -77
rect -40 -106 228 -98
rect -40 -107 218 -106
rect -40 -125 -15 -107
rect 245 -123 266 -40
rect -98 -133 -15 -125
rect -98 -154 -90 -133
rect -73 -154 -15 -133
rect -98 -159 -15 -154
rect 159 -139 191 -125
rect -98 -162 -69 -159
rect 159 -160 165 -139
rect 183 -160 191 -139
rect 159 -213 191 -160
rect 240 -126 266 -123
rect 240 -141 270 -126
rect 240 -162 245 -141
rect 263 -162 270 -141
rect 240 -170 270 -162
rect -92 -270 271 -213
<< metal1 >>
rect -100 118 278 161
rect -100 -278 280 -207
<< end >>
