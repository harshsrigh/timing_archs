.subckt vsdcell_nand3_2x A B C VGND VPWR Y
X0 Y A NET1 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X1 Y A NET1  VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X2 NET1 B NET2 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X3 NET1 B NET2 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X4 NET2 C VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X5 NET2 C VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X6 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X7 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u

X8 Y B VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X9 Y B VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u

X10 Y C VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X11 Y C VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
.ends