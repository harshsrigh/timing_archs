magic
tech sky130A
timestamp 1616056921
<< nwell >>
rect -2 169 436 301
rect 1 168 424 169
<< nmos >>
rect 46 40 61 82
rect 90 40 105 82
rect 137 40 152 82
rect 183 40 198 82
rect 230 40 245 82
rect 277 40 292 82
rect 326 40 341 82
rect 373 40 388 82
<< pmos >>
rect 46 205 61 255
rect 90 205 105 255
rect 137 205 152 255
rect 183 205 198 255
rect 230 205 245 255
rect 277 205 292 255
rect 326 205 341 255
rect 373 205 388 255
<< ndiff >>
rect 18 65 46 82
rect 18 48 22 65
rect 39 48 46 65
rect 18 40 46 48
rect 61 66 90 82
rect 61 49 67 66
rect 84 49 90 66
rect 61 40 90 49
rect 105 62 137 82
rect 105 45 114 62
rect 131 45 137 62
rect 105 40 137 45
rect 152 67 183 82
rect 152 50 159 67
rect 176 50 183 67
rect 152 40 183 50
rect 198 62 230 82
rect 198 45 206 62
rect 223 45 230 62
rect 198 40 230 45
rect 245 67 277 82
rect 245 50 254 67
rect 271 50 277 67
rect 245 40 277 50
rect 292 62 326 82
rect 292 45 300 62
rect 317 45 326 62
rect 292 40 326 45
rect 341 67 373 82
rect 341 50 349 67
rect 366 50 373 67
rect 341 40 373 50
rect 388 63 417 82
rect 388 46 396 63
rect 413 46 417 63
rect 388 40 417 46
<< pdiff >>
rect 16 244 46 255
rect 16 227 20 244
rect 37 227 46 244
rect 16 205 46 227
rect 61 241 90 255
rect 61 224 67 241
rect 84 224 90 241
rect 61 205 90 224
rect 105 244 137 255
rect 105 227 112 244
rect 129 227 137 244
rect 105 205 137 227
rect 152 241 183 255
rect 152 224 159 241
rect 176 224 183 241
rect 152 205 183 224
rect 198 244 230 255
rect 198 227 205 244
rect 222 227 230 244
rect 198 205 230 227
rect 245 240 277 255
rect 245 223 253 240
rect 270 223 277 240
rect 245 205 277 223
rect 292 244 326 255
rect 292 227 300 244
rect 317 227 326 244
rect 292 205 326 227
rect 341 240 373 255
rect 341 223 349 240
rect 366 223 373 240
rect 341 205 373 223
rect 388 244 418 255
rect 388 227 397 244
rect 414 227 418 244
rect 388 205 418 227
<< ndiffc >>
rect 22 48 39 65
rect 67 49 84 66
rect 114 45 131 62
rect 159 50 176 67
rect 206 45 223 62
rect 254 50 271 67
rect 300 45 317 62
rect 349 50 366 67
rect 396 46 413 63
<< pdiffc >>
rect 20 227 37 244
rect 67 224 84 241
rect 112 227 129 244
rect 159 224 176 241
rect 205 227 222 244
rect 253 223 270 240
rect 300 227 317 244
rect 349 223 366 240
rect 397 227 414 244
<< poly >>
rect 46 255 61 268
rect 90 255 105 268
rect 137 255 152 268
rect 183 255 198 268
rect 230 255 245 268
rect 277 255 292 268
rect 326 255 341 269
rect 373 255 388 269
rect 46 147 61 205
rect 90 147 105 205
rect 137 147 152 205
rect 183 147 198 205
rect 230 147 245 205
rect 277 147 292 205
rect 326 147 341 205
rect 373 147 388 205
rect 38 142 388 147
rect 38 125 46 142
rect 63 125 80 142
rect 97 125 114 142
rect 131 125 148 142
rect 165 125 182 142
rect 199 125 217 142
rect 234 125 251 142
rect 268 125 285 142
rect 302 125 319 142
rect 336 125 353 142
rect 370 125 388 142
rect 38 120 388 125
rect 46 82 61 120
rect 90 82 105 120
rect 137 82 152 120
rect 183 82 198 120
rect 230 82 245 120
rect 277 82 292 120
rect 326 82 341 120
rect 373 82 388 120
rect 46 23 61 40
rect 90 23 105 40
rect 137 23 152 40
rect 183 23 198 40
rect 230 23 245 40
rect 277 23 292 40
rect 326 24 341 40
rect 373 24 388 40
<< polycont >>
rect 46 125 63 142
rect 80 125 97 142
rect 114 125 131 142
rect 148 125 165 142
rect 182 125 199 142
rect 217 125 234 142
rect 251 125 268 142
rect 285 125 302 142
rect 319 125 336 142
rect 353 125 370 142
<< locali >>
rect 2 289 422 291
rect 2 272 4 289
rect 21 272 46 289
rect 63 272 84 289
rect 101 272 129 289
rect 146 272 171 289
rect 188 272 216 289
rect 233 272 255 289
rect 272 288 397 289
rect 272 272 301 288
rect 2 271 301 272
rect 318 271 348 288
rect 365 272 397 288
rect 414 272 422 289
rect 365 271 422 272
rect 2 270 422 271
rect 20 244 37 270
rect 20 219 37 227
rect 67 241 84 250
rect 67 188 84 224
rect 112 244 129 270
rect 112 219 129 227
rect 159 241 176 250
rect 159 188 176 224
rect 205 244 222 270
rect 205 218 222 227
rect 253 240 270 250
rect 253 188 270 223
rect 300 244 317 270
rect 300 218 317 227
rect 349 240 366 250
rect 349 188 366 223
rect 397 244 414 270
rect 397 218 414 227
rect 1 168 426 188
rect 1 108 18 168
rect 374 143 391 146
rect 38 142 391 143
rect 38 125 46 142
rect 63 125 80 142
rect 97 125 114 142
rect 131 125 148 142
rect 165 125 182 142
rect 199 125 217 142
rect 234 125 251 142
rect 268 125 285 142
rect 302 125 319 142
rect 336 125 353 142
rect 370 125 391 142
rect 409 108 426 168
rect 1 91 426 108
rect 14 65 43 73
rect 14 48 22 65
rect 39 48 43 65
rect 14 40 43 48
rect 67 66 84 91
rect 67 40 84 49
rect 114 62 131 70
rect 20 11 37 40
rect 3 10 37 11
rect 114 10 131 45
rect 159 67 176 91
rect 159 40 176 50
rect 206 62 223 70
rect 206 10 223 45
rect 254 67 271 91
rect 254 40 271 50
rect 300 62 317 70
rect 300 10 317 45
rect 349 67 366 91
rect 349 40 366 50
rect 396 63 413 71
rect 396 10 413 46
rect 3 9 421 10
rect 20 -8 45 9
rect 62 -8 87 9
rect 104 -8 129 9
rect 146 -8 172 9
rect 189 -8 216 9
rect 233 -8 258 9
rect 275 -8 301 9
rect 318 -8 347 9
rect 364 -8 396 9
rect 413 -8 421 9
rect 3 -10 421 -8
<< viali >>
rect 4 272 21 289
rect 46 272 63 289
rect 84 272 101 289
rect 129 272 146 289
rect 171 272 188 289
rect 216 272 233 289
rect 255 272 272 289
rect 301 271 318 288
rect 348 271 365 288
rect 397 272 414 289
rect 3 -8 20 9
rect 45 -8 62 9
rect 87 -8 104 9
rect 129 -8 146 9
rect 172 -8 189 9
rect 216 -8 233 9
rect 258 -8 275 9
rect 301 -8 318 9
rect 347 -8 364 9
rect 396 -8 413 9
<< metal1 >>
rect 0 289 431 299
rect 0 272 4 289
rect 21 272 46 289
rect 63 272 84 289
rect 101 272 129 289
rect 146 272 171 289
rect 188 272 216 289
rect 233 272 255 289
rect 272 288 397 289
rect 272 272 301 288
rect 0 271 301 272
rect 318 271 348 288
rect 365 272 397 288
rect 414 272 431 289
rect 365 271 431 272
rect 0 261 431 271
rect 20 219 37 261
rect 0 9 430 19
rect 0 -8 3 9
rect 20 -8 45 9
rect 62 -8 87 9
rect 104 -8 129 9
rect 146 -8 172 9
rect 189 -8 216 9
rect 233 -8 258 9
rect 275 -8 301 9
rect 318 -8 347 9
rect 364 -8 396 9
rect 413 -8 430 9
rect 0 -20 430 -8
<< labels >>
flabel locali 370 125 391 143 0 FreeSans 120 0 0 0 A
port 0 nsew signal input
flabel locali 409 91 426 188 0 FreeSans 120 0 0 0 Y
port 1 nsew signal output
flabel metal1 188 270 216 291 0 FreeSans 120 0 0 0 VPWR
port 3 nsew power bidirectional
flabel metal1 189 -10 216 10 0 FreeSans 120 0 0 0 VGND
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 428 278
<< end >>
