VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vsdcell_nand2_1x
  CLASS CORE ;
  FOREIGN vsdcell_nand2_1x ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.320 BY 2.720 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.305900 ;
    PORT
      LAYER li1 ;
        RECT 0.320 0.910 0.670 1.250 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.305900 ;
    PORT
      LAYER li1 ;
        RECT 1.690 0.960 2.030 1.240 ;
    END
  END B
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.200 1.220 2.420 3.050 ;
      LAYER li1 ;
        RECT -0.200 2.580 2.420 2.900 ;
        RECT 0.180 2.330 0.350 2.580 ;
        RECT 1.930 2.340 2.100 2.580 ;
        RECT 0.100 1.970 0.440 2.330 ;
        RECT 1.850 1.970 2.190 2.340 ;
      LAYER mcon ;
        RECT 0.530 2.640 0.700 2.810 ;
        RECT 1.330 2.650 1.500 2.820 ;
      LAYER met1 ;
        RECT -0.200 2.480 2.420 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.410 0.450 0.690 ;
        RECT 0.150 0.210 0.380 0.410 ;
        RECT -0.210 -0.150 2.420 0.210 ;
      LAYER mcon ;
        RECT 0.510 -0.090 0.680 0.080 ;
        RECT 1.300 -0.080 1.470 0.090 ;
      LAYER met1 ;
        RECT -0.210 -0.180 2.420 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.942900 ;
    PORT
      LAYER li1 ;
        RECT 0.940 1.960 1.280 2.330 ;
        RECT 1.060 1.790 1.230 1.960 ;
        RECT 0.950 1.280 1.400 1.790 ;
        RECT 1.060 0.760 1.230 1.280 ;
        RECT 1.060 0.410 2.180 0.760 ;
    END
  END Y
END vsdcell_nand2_1x
END LIBRARY

