* SPICE3 file created from nand_4.ext - technology: sky130A

.option scale=10000u

.subckt nand_4 A VPWR VGND B C D Y
X0 a_67_30# A VGND SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X1 a_176_30# C a_127_30# SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X2 VPWR B Y w_n10_170# sky130_fd_pr__pfet_01v8 w=50 l=15
X3 Y A VPWR w_n10_170# sky130_fd_pr__pfet_01v8 w=50 l=15
X4 VPWR D Y w_n10_170# sky130_fd_pr__pfet_01v8 w=50 l=16
X5 a_127_30# B a_67_30# SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X6 Y C VPWR w_n10_170# sky130_fd_pr__pfet_01v8 w=50 l=15
X7 Y D a_176_30# SUB sky130_fd_pr__nfet_01v8 w=42 l=16
.ends
