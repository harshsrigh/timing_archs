* SPICE3 file created from sky130_vsd_buf2.ext - technology: sky130A

.option scale=10000u

.subckt sky130_vsd_buf2 X A VPWR VGND
X0 VPWR a_42_7# X w_n8_158# sky130_fd_pr__pfet_01v8 w=60 l=15
X1 a_42_7# A VGND SUB sky130_fd_pr__nfet_01v8 w=42 l=17
X2 a_42_7# A VPWR w_n8_158# sky130_fd_pr__pfet_01v8 w=60 l=17
X3 VGND a_42_7# X SUB sky130_fd_pr__nfet_01v8 w=42 l=15
.ends
