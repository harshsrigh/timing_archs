
.subckt vsdcell_and4_2x A B C D VGND VPWR Y

X6 net4 A net3 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X0 net4 A VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X1 net4 A VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X2 net4 B VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X3 net4 B VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X5 net4 A net3 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X7 net3 B net2 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X8 net3 B net2 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X10 net4 C VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X11 net4 C VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X12 net2 C net8 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X13 net2 C net8 VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X4 Y net4 VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X9 Y net4 VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X14 net4 D VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X15 net4 D VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u 
X16 net8 D VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 
X17 net8 D VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u 

.ends
