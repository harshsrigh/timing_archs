magic
tech sky130A
timestamp 1616064524
<< nwell >>
rect -10 170 185 300
<< nmos >>
rect 52 30 67 72
rect 112 30 127 72
<< pmos >>
rect 52 190 67 240
rect 112 190 127 240
<< ndiff >>
rect 10 60 52 72
rect 10 40 20 60
rect 40 40 52 60
rect 10 30 52 40
rect 67 30 112 72
rect 127 63 164 72
rect 127 43 135 63
rect 155 43 164 63
rect 127 30 164 43
<< pdiff >>
rect 10 230 52 240
rect 10 210 20 230
rect 40 210 52 230
rect 10 190 52 210
rect 67 229 112 240
rect 67 209 84 229
rect 104 209 112 229
rect 67 190 112 209
rect 127 230 165 240
rect 127 210 135 230
rect 155 210 165 230
rect 127 190 165 210
<< ndiffc >>
rect 20 40 40 60
rect 135 43 155 63
<< pdiffc >>
rect 20 210 40 230
rect 84 209 104 229
rect 135 210 155 230
<< poly >>
rect 52 240 67 253
rect 112 240 127 253
rect 52 141 67 190
rect 31 131 67 141
rect 31 110 36 131
rect 56 110 67 131
rect 31 102 67 110
rect 52 72 67 102
rect 112 165 127 190
rect 112 157 150 165
rect 112 136 125 157
rect 145 136 150 157
rect 112 126 150 136
rect 112 72 127 126
rect 52 17 67 30
rect 112 17 127 30
<< polycont >>
rect 36 110 56 131
rect 125 136 145 157
<< locali >>
rect 0 287 173 291
rect 0 270 31 287
rect 48 270 132 287
rect 149 270 173 287
rect 0 264 173 270
rect 20 230 40 264
rect 12 210 20 230
rect 40 210 48 230
rect 12 202 48 210
rect 84 229 104 240
rect 31 131 59 141
rect 31 110 36 131
rect 56 110 59 131
rect 31 102 59 110
rect 84 109 104 209
rect 135 230 155 264
rect 135 200 155 210
rect 122 157 150 165
rect 122 136 125 157
rect 145 136 150 157
rect 122 126 150 136
rect 84 83 155 109
rect 12 60 48 69
rect 12 40 20 60
rect 40 40 48 60
rect 12 39 48 40
rect 135 63 155 83
rect 20 10 40 39
rect 135 35 155 43
rect 10 9 175 10
rect 10 -8 36 9
rect 53 -8 133 9
rect 150 -8 175 9
rect 10 -10 175 -8
<< viali >>
rect 31 270 48 287
rect 132 270 149 287
rect 36 -8 53 9
rect 133 -8 150 9
<< metal1 >>
rect 0 287 178 300
rect 0 270 31 287
rect 48 270 132 287
rect 149 270 178 287
rect 0 255 178 270
rect 0 9 180 20
rect 0 -8 36 9
rect 53 -8 133 9
rect 150 -8 180 9
rect 0 -20 180 -8
<< labels >>
flabel polycont 36 110 56 131 0 FreeSans 120 0 0 0 A
port 0 nsew signal input
flabel polycont 125 136 145 157 0 FreeSans 120 0 0 0 B
port 1 nsew signal input
flabel locali 84 83 104 209 0 FreeSans 120 0 0 0 Y
port 2 nsew signal output
flabel locali 0 264 173 291 0 FreeSans 120 0 0 0 VPWR
port 3 nsew power bidirectional
flabel locali 10 -10 175 10 0 FreeSans 120 0 0 0 VGND
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 175 278
<< end >>
