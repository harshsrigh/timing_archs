* SPICE3 file created from sky130_vsdclkbuf_1x.ext - technology: sky130A

.option scale=0.01u

.subckt sky130_vsdclkbuf_1x A Y VGND VPWR VPB
X0 a_34_100# A VPWR VPB sky130_fd_pr__pfet_01v8 w=70 l=15
X1 VGND a_34_100# Y VGND sky130_fd_pr__nfet_01v8 w=43 l=15
X2 a_34_100# A VGND VGND sky130_fd_pr__nfet_01v8 w=43 l=15
X3 VPWR a_34_100# Y VPB sky130_fd_pr__pfet_01v8 w=70 l=15
C0 VPWR a_34_100# 0.19fF
C1 VPWR A 0.03fF
C2 Y VPB 0.00fF
C3 Y a_34_100# 0.12fF
C4 Y A 0.01fF
C5 VPB a_34_100# 0.00fF
C6 Y VPWR 0.12fF
C7 A a_34_100# 0.13fF
C8 VPWR VPB 0.02fF
C9 VPWR VGND 0.33fF
C10 Y VGND 0.21fF
C11 VPB VGND 0.25fF
C12 a_34_100# VGND 0.53fF
.ends
