VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_vsdclkbuf_1x
  CLASS CORE ;
  FOREIGN sky130_vsdclkbuf_1x ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.690 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.169500 ;
    PORT
      LAYER li1 ;
        RECT 0.880 1.190 1.210 1.470 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.421300 ;
    PORT
      LAYER li1 ;
        RECT 0.000 1.660 0.300 2.360 ;
        RECT 0.000 0.830 0.170 1.660 ;
        RECT 0.000 0.400 0.360 0.830 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.590 0.180 0.940 0.830 ;
        RECT 0.000 -0.120 1.680 0.180 ;
      LAYER mcon ;
        RECT 0.210 -0.080 0.380 0.100 ;
        RECT 0.570 -0.080 0.740 0.100 ;
        RECT 0.930 -0.080 1.100 0.100 ;
        RECT 1.290 -0.080 1.460 0.100 ;
      LAYER met1 ;
        RECT 0.000 -0.170 1.680 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.570 1.690 2.870 ;
        RECT 0.650 1.670 0.940 2.570 ;
      LAYER mcon ;
        RECT 0.220 2.630 0.390 2.810 ;
        RECT 0.580 2.630 0.750 2.810 ;
        RECT 0.940 2.630 1.110 2.810 ;
        RECT 1.300 2.630 1.470 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.490 1.690 2.910 ;
    END
  END VPWR
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.130 1.460 1.800 2.880 ;
    END
  END VPB
  OBS
      LAYER li1 ;
        RECT 1.280 1.660 1.640 2.360 ;
        RECT 0.340 1.000 0.670 1.280 ;
        RECT 1.460 0.830 1.640 1.660 ;
        RECT 1.310 0.400 1.640 0.830 ;
      LAYER mcon ;
        RECT 0.420 1.050 0.590 1.230 ;
        RECT 1.460 1.010 1.640 1.180 ;
      LAYER met1 ;
        RECT 0.340 1.170 0.670 1.280 ;
        RECT 1.410 1.170 1.680 1.240 ;
        RECT 0.340 1.000 1.680 1.170 ;
        RECT 1.410 0.950 1.680 1.000 ;
  END
END sky130_vsdclkbuf_1x
END LIBRARY

