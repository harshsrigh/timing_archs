* SPICE3 file created from sky130_vsd_conb.ext - technology: sky130A

.option scale=10000u

.subckt sky130_vsd_conb HI LO VGND VPWR
X0 VPWR LO HI w_n13_156# sky130_fd_pr__pfet_01v8 w=60 l=15
X1 VGND LO LO SUB sky130_fd_pr__nfet_01v8 w=42 l=15
X2 HI HI VPWR w_n13_156# sky130_fd_pr__pfet_01v8 w=60 l=15
X3 LO HI VGND SUB sky130_fd_pr__nfet_01v8 w=42 l=15
.ends
