magic
tech sky130A
timestamp 1615276334
<< nwell >>
rect -20 122 242 305
<< nmos >>
rect 49 41 72 83
rect 159 41 182 83
<< pmos >>
rect 49 143 72 234
rect 159 143 182 234
<< ndiff >>
rect 10 62 49 83
rect 10 45 19 62
rect 36 45 49 62
rect 10 41 49 45
rect 72 41 159 83
rect 182 62 218 83
rect 182 45 192 62
rect 209 45 218 62
rect 182 41 218 45
<< pdiff >>
rect 7 228 49 234
rect 7 203 18 228
rect 36 203 49 228
rect 7 143 49 203
rect 72 227 159 234
rect 72 202 102 227
rect 120 202 159 227
rect 72 143 159 202
rect 182 228 219 234
rect 182 203 193 228
rect 211 203 219 228
rect 182 196 219 203
rect 182 143 218 196
<< ndiffc >>
rect 19 45 36 62
rect 192 45 209 62
<< pdiffc >>
rect 18 203 36 228
rect 102 202 120 227
rect 193 203 211 228
<< psubdiff >>
rect -21 13 129 14
rect -21 -7 76 13
rect 12 -8 76 -7
rect 93 -8 110 13
rect 127 -8 242 13
rect 112 -9 129 -8
<< nsubdiff >>
rect 12 285 130 286
rect 12 261 75 285
rect 93 261 110 285
rect 128 261 203 285
<< psubdiffcont >>
rect 76 -8 93 13
rect 110 -8 127 13
<< nsubdiffcont >>
rect 75 261 93 285
rect 110 261 128 285
<< poly >>
rect 49 234 72 250
rect 159 234 182 250
rect 49 125 72 143
rect 32 119 72 125
rect 32 102 42 119
rect 59 102 72 119
rect 32 91 72 102
rect 49 83 72 91
rect 159 124 182 143
rect 159 119 203 124
rect 159 102 178 119
rect 195 102 203 119
rect 159 96 203 102
rect 159 83 182 96
rect 49 27 72 41
rect 159 26 182 41
<< polycont >>
rect 42 102 59 119
rect 178 102 195 119
<< locali >>
rect -20 285 242 290
rect -20 281 75 285
rect -20 264 53 281
rect 70 264 75 281
rect -20 261 75 264
rect 93 261 110 285
rect 128 282 242 285
rect 128 265 133 282
rect 150 265 242 282
rect 128 261 242 265
rect -20 258 242 261
rect 18 233 35 258
rect 193 234 210 258
rect 10 228 44 233
rect 10 203 18 228
rect 36 203 44 228
rect 10 197 44 203
rect 94 227 128 233
rect 94 202 102 227
rect 120 202 128 227
rect 94 196 128 202
rect 185 228 219 234
rect 185 203 193 228
rect 211 203 219 228
rect 185 197 219 203
rect 106 179 123 196
rect 95 128 140 179
rect 32 119 67 125
rect 32 102 42 119
rect 59 102 67 119
rect 32 91 67 102
rect 106 76 123 128
rect 169 119 203 124
rect 169 102 178 119
rect 195 102 203 119
rect 169 96 203 102
rect 10 62 45 69
rect 10 45 19 62
rect 36 45 45 62
rect 10 41 45 45
rect 106 62 218 76
rect 106 45 192 62
rect 209 45 218 62
rect 106 41 218 45
rect 15 21 38 41
rect -21 13 242 21
rect -21 8 76 13
rect -21 -9 51 8
rect 68 -8 76 8
rect 93 -8 110 13
rect 127 9 242 13
rect 127 -8 130 9
rect 147 -8 242 9
rect 68 -9 242 -8
rect -21 -15 242 -9
<< viali >>
rect 53 264 70 281
rect 133 265 150 282
rect 51 -9 68 8
rect 130 -8 147 9
<< metal1 >>
rect -20 282 242 296
rect -20 281 133 282
rect -20 264 53 281
rect 70 265 133 281
rect 150 265 242 282
rect 70 264 242 265
rect -20 248 242 264
rect -21 9 242 24
rect -21 8 130 9
rect -21 -9 51 8
rect 68 -8 130 8
rect 147 -8 242 9
rect 68 -9 242 -8
rect -21 -18 242 -9
<< labels >>
flabel locali 104 139 135 173 0 FreeSans 184 0 0 0 Y
port 5 nsew signal output
flabel locali 36 93 65 123 0 FreeSans 184 0 0 0 A
port 1 nsew signal input
flabel locali 173 97 200 124 0 FreeSans 184 0 0 0 B
port 2 nsew signal input
flabel metal1 72 255 132 292 0 FreeSans 184 0 0 0 VPWR
port 3 nsew power bidirectional
flabel metal1 73 -14 129 19 0 FreeSans 120 0 0 0 VGND
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 232 272
string LEFsource USER
string LEForigin 0 0
<< end >>
