VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_vsddfxtp_1
  CLASS CORE ;
  FOREIGN sky130_vsddfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.297000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.100 0.380 1.490 ;
        RECT 1.210 1.150 1.500 1.490 ;
      LAYER mcon ;
        RECT 0.150 1.230 0.320 1.410 ;
        RECT 1.270 1.230 1.440 1.410 ;
      LAYER met1 ;
        RECT 0.090 1.410 0.380 1.490 ;
        RECT 1.210 1.410 1.500 1.490 ;
        RECT 0.090 1.230 1.500 1.410 ;
        RECT 0.090 1.100 0.380 1.230 ;
        RECT 1.210 1.150 1.500 1.230 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.508500 ;
    ANTENNADIFFAREA 0.259300 ;
    PORT
      LAYER li1 ;
        RECT 0.580 0.400 0.820 2.360 ;
        RECT 2.130 1.000 3.100 1.300 ;
        RECT 3.680 1.000 4.020 1.280 ;
      LAYER mcon ;
        RECT 2.210 1.050 2.380 1.230 ;
        RECT 2.850 1.060 3.020 1.240 ;
        RECT 3.770 1.050 3.940 1.230 ;
        RECT 0.610 0.800 0.780 0.980 ;
      LAYER met1 ;
        RECT 2.770 1.260 3.100 1.270 ;
        RECT 2.130 1.250 2.460 1.260 ;
        RECT 2.770 1.250 3.120 1.260 ;
        RECT 3.680 1.250 4.020 1.270 ;
        RECT 2.130 1.230 4.020 1.250 ;
        RECT 1.690 1.160 4.020 1.230 ;
        RECT 1.680 1.070 4.020 1.160 ;
        RECT 0.580 1.000 0.820 1.040 ;
        RECT 1.680 1.000 1.920 1.070 ;
        RECT 2.130 1.010 3.100 1.070 ;
        RECT 2.130 1.000 2.800 1.010 ;
        RECT 3.680 1.000 4.020 1.070 ;
        RECT 0.580 0.840 1.920 1.000 ;
        RECT 0.580 0.690 0.820 0.840 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.169500 ;
    ANTENNADIFFAREA 0.403100 ;
    PORT
      LAYER li1 ;
        RECT 5.360 1.000 5.700 1.280 ;
        RECT 6.590 0.760 6.830 2.360 ;
        RECT 7.120 0.760 7.340 0.830 ;
        RECT 6.590 0.570 7.340 0.760 ;
        RECT 7.120 0.480 7.340 0.570 ;
      LAYER mcon ;
        RECT 6.630 1.750 6.800 1.930 ;
        RECT 5.450 1.050 5.620 1.230 ;
      LAYER met1 ;
        RECT 5.360 1.080 5.840 1.270 ;
        RECT 6.590 1.080 6.830 2.050 ;
        RECT 5.360 1.000 6.830 1.080 ;
        RECT 5.700 0.940 6.830 1.000 ;
    END
  END Q
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.060 0.200 0.300 0.830 ;
        RECT 1.100 0.200 1.330 0.830 ;
        RECT 2.700 0.200 2.920 0.830 ;
        RECT 4.380 0.200 4.600 0.830 ;
        RECT 6.020 0.200 6.240 0.830 ;
        RECT 0.020 -0.110 7.400 0.200 ;
        RECT 4.330 -0.120 4.770 -0.110 ;
        RECT 5.970 -0.120 6.410 -0.110 ;
      LAYER mcon ;
        RECT 0.140 -0.100 0.310 0.080 ;
        RECT 0.500 -0.100 0.670 0.080 ;
        RECT 0.860 -0.100 1.030 0.080 ;
        RECT 1.220 -0.100 1.390 0.080 ;
        RECT 1.580 -0.100 1.750 0.080 ;
        RECT 1.940 -0.100 2.110 0.080 ;
        RECT 2.300 -0.100 2.470 0.080 ;
        RECT 2.660 -0.100 2.830 0.080 ;
        RECT 3.020 -0.100 3.190 0.080 ;
        RECT 3.380 -0.100 3.550 0.080 ;
        RECT 3.740 -0.100 3.910 0.080 ;
        RECT 4.100 -0.100 4.270 0.080 ;
        RECT 4.460 -0.100 4.630 0.080 ;
        RECT 4.820 -0.100 4.990 0.080 ;
        RECT 5.180 -0.100 5.350 0.080 ;
        RECT 5.540 -0.100 5.710 0.080 ;
        RECT 5.900 -0.100 6.070 0.080 ;
        RECT 6.260 -0.100 6.430 0.080 ;
        RECT 6.620 -0.100 6.790 0.080 ;
        RECT 6.980 -0.100 7.150 0.080 ;
      LAYER met1 ;
        RECT 0.000 -0.210 7.420 0.250 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.060 0.200 0.300 0.830 ;
        RECT 1.100 0.200 1.330 0.830 ;
        RECT 2.700 0.200 2.920 0.830 ;
        RECT 4.380 0.200 4.600 0.830 ;
        RECT 6.020 0.200 6.240 0.830 ;
        RECT 0.020 -0.110 7.400 0.200 ;
        RECT 4.330 -0.120 4.770 -0.110 ;
        RECT 5.970 -0.120 6.410 -0.110 ;
      LAYER mcon ;
        RECT 0.140 -0.100 0.310 0.080 ;
        RECT 0.500 -0.100 0.670 0.080 ;
        RECT 0.860 -0.100 1.030 0.080 ;
        RECT 1.220 -0.100 1.390 0.080 ;
        RECT 1.580 -0.100 1.750 0.080 ;
        RECT 1.940 -0.100 2.110 0.080 ;
        RECT 2.300 -0.100 2.470 0.080 ;
        RECT 2.660 -0.100 2.830 0.080 ;
        RECT 3.020 -0.100 3.190 0.080 ;
        RECT 3.380 -0.100 3.550 0.080 ;
        RECT 3.740 -0.100 3.910 0.080 ;
        RECT 4.100 -0.100 4.270 0.080 ;
        RECT 4.460 -0.100 4.630 0.080 ;
        RECT 4.820 -0.100 4.990 0.080 ;
        RECT 5.180 -0.100 5.350 0.080 ;
        RECT 5.540 -0.100 5.710 0.080 ;
        RECT 5.900 -0.100 6.070 0.080 ;
        RECT 6.260 -0.100 6.430 0.080 ;
        RECT 6.620 -0.100 6.790 0.080 ;
        RECT 6.980 -0.100 7.150 0.080 ;
      LAYER met1 ;
        RECT 0.000 -0.210 7.420 0.250 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.020 2.570 7.420 2.870 ;
        RECT 0.060 1.970 0.300 2.570 ;
        RECT 1.140 1.660 1.380 2.570 ;
        RECT 2.220 1.660 2.450 2.570 ;
        RECT 2.730 1.660 2.970 2.570 ;
        RECT 3.810 1.660 4.040 2.570 ;
        RECT 4.410 1.660 4.650 2.570 ;
        RECT 5.490 1.660 5.720 2.570 ;
        RECT 6.050 1.660 6.290 2.570 ;
        RECT 7.130 1.660 7.360 2.570 ;
      LAYER mcon ;
        RECT 0.170 2.630 0.340 2.810 ;
        RECT 0.530 2.630 0.700 2.810 ;
        RECT 0.890 2.630 1.060 2.810 ;
        RECT 1.250 2.630 1.420 2.810 ;
        RECT 1.610 2.630 1.780 2.810 ;
        RECT 1.970 2.630 2.140 2.810 ;
        RECT 2.330 2.630 2.500 2.810 ;
        RECT 2.690 2.630 2.860 2.810 ;
        RECT 3.050 2.630 3.220 2.810 ;
        RECT 3.410 2.630 3.580 2.810 ;
        RECT 3.770 2.630 3.940 2.810 ;
        RECT 4.130 2.630 4.300 2.810 ;
        RECT 4.490 2.630 4.660 2.810 ;
        RECT 4.850 2.630 5.020 2.810 ;
        RECT 5.210 2.630 5.380 2.810 ;
        RECT 5.570 2.630 5.740 2.810 ;
        RECT 5.930 2.630 6.100 2.810 ;
        RECT 6.290 2.630 6.460 2.810 ;
        RECT 6.650 2.630 6.820 2.810 ;
        RECT 7.010 2.630 7.180 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.500 7.420 2.900 ;
    END
  END VPWR
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.130 1.420 7.550 2.890 ;
    END
  END VPB
  OBS
      LAYER li1 ;
        RECT 1.680 0.760 1.920 2.360 ;
        RECT 2.210 0.760 2.430 0.830 ;
        RECT 1.680 0.570 2.430 0.760 ;
        RECT 3.270 0.760 3.510 2.360 ;
        RECT 4.440 1.000 4.780 1.280 ;
        RECT 3.770 0.760 4.020 0.830 ;
        RECT 3.270 0.570 4.020 0.760 ;
        RECT 4.950 0.760 5.190 2.360 ;
        RECT 6.130 1.150 6.420 1.490 ;
        RECT 7.000 1.040 7.340 1.320 ;
        RECT 5.460 0.760 5.700 0.830 ;
        RECT 4.950 0.570 5.700 0.760 ;
        RECT 2.210 0.480 2.430 0.570 ;
        RECT 3.770 0.480 4.020 0.570 ;
        RECT 5.480 0.480 5.700 0.570 ;
      LAYER mcon ;
        RECT 1.720 1.810 1.890 1.990 ;
        RECT 1.710 1.440 1.880 1.620 ;
        RECT 4.530 1.050 4.700 1.230 ;
        RECT 3.810 0.570 3.980 0.750 ;
        RECT 6.170 1.310 6.340 1.490 ;
        RECT 7.090 1.090 7.260 1.270 ;
        RECT 5.490 0.560 5.660 0.740 ;
      LAYER met1 ;
        RECT 1.680 1.550 1.920 2.050 ;
        RECT 1.680 1.490 6.370 1.550 ;
        RECT 1.680 1.410 6.420 1.490 ;
        RECT 1.680 1.380 1.920 1.410 ;
        RECT 4.440 1.140 4.780 1.270 ;
        RECT 6.130 1.220 6.420 1.410 ;
        RECT 4.160 1.000 4.780 1.140 ;
        RECT 7.000 1.040 7.350 1.310 ;
        RECT 3.770 0.750 4.020 0.830 ;
        RECT 4.160 0.750 4.320 1.000 ;
        RECT 3.770 0.580 4.320 0.750 ;
        RECT 5.460 0.760 5.700 0.800 ;
        RECT 7.120 0.760 7.350 1.040 ;
        RECT 3.770 0.480 4.020 0.580 ;
        RECT 5.460 0.570 7.350 0.760 ;
        RECT 5.460 0.560 7.340 0.570 ;
        RECT 5.460 0.480 5.700 0.560 ;
  END
END sky130_vsddfxtp_1
END LIBRARY

